magic
tech sky130A
magscale 1 2
timestamp 1685205180
<< viali >>
rect 11989 20553 12023 20587
rect 12725 20553 12759 20587
rect 15301 20553 15335 20587
rect 17785 20553 17819 20587
rect 18705 20553 18739 20587
rect 19717 20553 19751 20587
rect 20085 20553 20119 20587
rect 22017 20553 22051 20587
rect 31677 20553 31711 20587
rect 27445 20485 27479 20519
rect 30205 20485 30239 20519
rect 12173 20417 12207 20451
rect 12909 20417 12943 20451
rect 14657 20417 14691 20451
rect 15485 20417 15519 20451
rect 16313 20417 16347 20451
rect 17049 20417 17083 20451
rect 17969 20417 18003 20451
rect 18889 20417 18923 20451
rect 21097 20417 21131 20451
rect 22201 20417 22235 20451
rect 23397 20417 23431 20451
rect 24777 20417 24811 20451
rect 25421 20417 25455 20451
rect 26065 20417 26099 20451
rect 17233 20349 17267 20383
rect 20177 20349 20211 20383
rect 20269 20349 20303 20383
rect 23213 20349 23247 20383
rect 27169 20349 27203 20383
rect 29929 20349 29963 20383
rect 14473 20281 14507 20315
rect 20913 20281 20947 20315
rect 24593 20281 24627 20315
rect 25881 20281 25915 20315
rect 16129 20213 16163 20247
rect 16865 20213 16899 20247
rect 23581 20213 23615 20247
rect 25237 20213 25271 20247
rect 28917 20213 28951 20247
rect 2237 20009 2271 20043
rect 3065 20009 3099 20043
rect 4353 20009 4387 20043
rect 5089 20009 5123 20043
rect 5825 20009 5859 20043
rect 6561 20009 6595 20043
rect 10517 20009 10551 20043
rect 11253 20009 11287 20043
rect 13553 20009 13587 20043
rect 14381 20009 14415 20043
rect 15301 20009 15335 20043
rect 18889 20009 18923 20043
rect 24593 20009 24627 20043
rect 22569 19941 22603 19975
rect 23673 19941 23707 19975
rect 12173 19873 12207 19907
rect 14749 19873 14783 19907
rect 15945 19873 15979 19907
rect 16589 19873 16623 19907
rect 16773 19873 16807 19907
rect 18613 19873 18647 19907
rect 19993 19873 20027 19907
rect 21189 19873 21223 19907
rect 23397 19873 23431 19907
rect 26157 19873 26191 19907
rect 29193 19873 29227 19907
rect 2421 19805 2455 19839
rect 2881 19805 2915 19839
rect 4169 19805 4203 19839
rect 4905 19805 4939 19839
rect 5641 19805 5675 19839
rect 6377 19805 6411 19839
rect 10701 19805 10735 19839
rect 13737 19805 13771 19839
rect 14565 19805 14599 19839
rect 15669 19805 15703 19839
rect 17877 19805 17911 19839
rect 18521 19805 18555 19839
rect 19809 19805 19843 19839
rect 21005 19805 21039 19839
rect 23305 19805 23339 19839
rect 25421 19805 25455 19839
rect 31493 19805 31527 19839
rect 11529 19737 11563 19771
rect 12449 19737 12483 19771
rect 16865 19737 16899 19771
rect 22201 19737 22235 19771
rect 24777 19737 24811 19771
rect 24961 19737 24995 19771
rect 26433 19737 26467 19771
rect 15761 19669 15795 19703
rect 17233 19669 17267 19703
rect 17693 19669 17727 19703
rect 19441 19669 19475 19703
rect 19901 19669 19935 19703
rect 20637 19669 20671 19703
rect 21097 19669 21131 19703
rect 22661 19669 22695 19703
rect 25605 19669 25639 19703
rect 27905 19669 27939 19703
rect 28549 19669 28583 19703
rect 30205 19669 30239 19703
rect 2421 19465 2455 19499
rect 3893 19465 3927 19499
rect 10977 19465 11011 19499
rect 12449 19465 12483 19499
rect 13185 19465 13219 19499
rect 14841 19465 14875 19499
rect 16129 19465 16163 19499
rect 20453 19465 20487 19499
rect 20821 19465 20855 19499
rect 22017 19465 22051 19499
rect 23121 19465 23155 19499
rect 24133 19465 24167 19499
rect 28917 19465 28951 19499
rect 14013 19397 14047 19431
rect 15209 19397 15243 19431
rect 17325 19397 17359 19431
rect 19625 19397 19659 19431
rect 27445 19397 27479 19431
rect 31769 19397 31803 19431
rect 2605 19329 2639 19363
rect 4077 19329 4111 19363
rect 11161 19329 11195 19363
rect 12633 19329 12667 19363
rect 13369 19329 13403 19363
rect 14197 19329 14231 19363
rect 14381 19329 14415 19363
rect 16313 19329 16347 19363
rect 18245 19329 18279 19363
rect 20913 19329 20947 19363
rect 22201 19329 22235 19363
rect 24133 19329 24167 19363
rect 24317 19329 24351 19363
rect 13553 19261 13587 19295
rect 15301 19261 15335 19295
rect 15485 19261 15519 19295
rect 19717 19261 19751 19295
rect 19901 19261 19935 19295
rect 21005 19261 21039 19295
rect 23305 19261 23339 19295
rect 23397 19261 23431 19295
rect 23489 19261 23523 19295
rect 23581 19261 23615 19295
rect 24869 19261 24903 19295
rect 26341 19261 26375 19295
rect 26617 19261 26651 19295
rect 27169 19261 27203 19295
rect 29745 19261 29779 19295
rect 30021 19261 30055 19295
rect 17049 19193 17083 19227
rect 18061 19193 18095 19227
rect 19257 19193 19291 19227
rect 11529 18921 11563 18955
rect 13369 18921 13403 18955
rect 15025 18921 15059 18955
rect 15853 18921 15887 18955
rect 17141 18921 17175 18955
rect 19717 18921 19751 18955
rect 20729 18921 20763 18955
rect 23029 18921 23063 18955
rect 20269 18853 20303 18887
rect 24041 18853 24075 18887
rect 25237 18853 25271 18887
rect 22753 18785 22787 18819
rect 23581 18785 23615 18819
rect 29193 18785 29227 18819
rect 11713 18717 11747 18751
rect 13553 18717 13587 18751
rect 13737 18717 13771 18751
rect 15209 18717 15243 18751
rect 15393 18717 15427 18751
rect 16037 18717 16071 18751
rect 16221 18717 16255 18751
rect 17325 18717 17359 18751
rect 20085 18717 20119 18751
rect 20913 18717 20947 18751
rect 22661 18717 22695 18751
rect 23673 18717 23707 18751
rect 24593 18717 24627 18751
rect 24777 18717 24811 18751
rect 25421 18717 25455 18751
rect 26341 18717 26375 18751
rect 30021 18717 30055 18751
rect 19993 18649 20027 18683
rect 24685 18649 24719 18683
rect 26617 18649 26651 18683
rect 30297 18649 30331 18683
rect 19901 18581 19935 18615
rect 28089 18581 28123 18615
rect 31769 18581 31803 18615
rect 15669 18377 15703 18411
rect 19809 18377 19843 18411
rect 22845 18377 22879 18411
rect 23765 18377 23799 18411
rect 25145 18377 25179 18411
rect 27629 18377 27663 18411
rect 31309 18377 31343 18411
rect 19625 18309 19659 18343
rect 20177 18309 20211 18343
rect 22997 18309 23031 18343
rect 23213 18309 23247 18343
rect 23949 18309 23983 18343
rect 15853 18241 15887 18275
rect 16037 18241 16071 18275
rect 19901 18241 19935 18275
rect 19993 18241 20027 18275
rect 23673 18241 23707 18275
rect 24409 18241 24443 18275
rect 25053 18241 25087 18275
rect 29377 18241 29411 18275
rect 30021 18241 30055 18275
rect 23949 18105 23983 18139
rect 24593 18105 24627 18139
rect 23029 18037 23063 18071
rect 29113 18037 29147 18071
rect 26341 17833 26375 17867
rect 30849 17833 30883 17867
rect 31493 17833 31527 17867
rect 27813 17629 27847 17663
rect 31033 17629 31067 17663
rect 31677 17629 31711 17663
<< metal1 >>
rect 23658 21020 23664 21072
rect 23716 21060 23722 21072
rect 26050 21060 26056 21072
rect 23716 21032 26056 21060
rect 23716 21020 23722 21032
rect 26050 21020 26056 21032
rect 26108 21020 26114 21072
rect 20070 20952 20076 21004
rect 20128 20992 20134 21004
rect 25222 20992 25228 21004
rect 20128 20964 25228 20992
rect 20128 20952 20134 20964
rect 25222 20952 25228 20964
rect 25280 20952 25286 21004
rect 18506 20884 18512 20936
rect 18564 20924 18570 20936
rect 24854 20924 24860 20936
rect 18564 20896 24860 20924
rect 18564 20884 18570 20896
rect 24854 20884 24860 20896
rect 24912 20884 24918 20936
rect 18874 20816 18880 20868
rect 18932 20856 18938 20868
rect 30190 20856 30196 20868
rect 18932 20828 30196 20856
rect 18932 20816 18938 20828
rect 30190 20816 30196 20828
rect 30248 20816 30254 20868
rect 21082 20748 21088 20800
rect 21140 20788 21146 20800
rect 30834 20788 30840 20800
rect 21140 20760 30840 20788
rect 21140 20748 21146 20760
rect 30834 20748 30840 20760
rect 30892 20748 30898 20800
rect 1104 20698 32632 20720
rect 1104 20646 8792 20698
rect 8844 20646 8856 20698
rect 8908 20646 8920 20698
rect 8972 20646 8984 20698
rect 9036 20646 9048 20698
rect 9100 20646 16634 20698
rect 16686 20646 16698 20698
rect 16750 20646 16762 20698
rect 16814 20646 16826 20698
rect 16878 20646 16890 20698
rect 16942 20646 24476 20698
rect 24528 20646 24540 20698
rect 24592 20646 24604 20698
rect 24656 20646 24668 20698
rect 24720 20646 24732 20698
rect 24784 20646 32318 20698
rect 32370 20646 32382 20698
rect 32434 20646 32446 20698
rect 32498 20646 32510 20698
rect 32562 20646 32574 20698
rect 32626 20646 32632 20698
rect 1104 20624 32632 20646
rect 11974 20544 11980 20596
rect 12032 20544 12038 20596
rect 12710 20544 12716 20596
rect 12768 20544 12774 20596
rect 14826 20544 14832 20596
rect 14884 20584 14890 20596
rect 15289 20587 15347 20593
rect 15289 20584 15301 20587
rect 14884 20556 15301 20584
rect 14884 20544 14890 20556
rect 15289 20553 15301 20556
rect 15335 20553 15347 20587
rect 15289 20547 15347 20553
rect 15562 20544 15568 20596
rect 15620 20584 15626 20596
rect 15620 20556 17724 20584
rect 15620 20544 15626 20556
rect 15838 20516 15844 20528
rect 12176 20488 15844 20516
rect 12176 20457 12204 20488
rect 15838 20476 15844 20488
rect 15896 20476 15902 20528
rect 12161 20451 12219 20457
rect 12161 20417 12173 20451
rect 12207 20417 12219 20451
rect 12161 20411 12219 20417
rect 12897 20451 12955 20457
rect 12897 20417 12909 20451
rect 12943 20448 12955 20451
rect 14366 20448 14372 20460
rect 12943 20420 14372 20448
rect 12943 20417 12955 20420
rect 12897 20411 12955 20417
rect 14366 20408 14372 20420
rect 14424 20408 14430 20460
rect 14642 20408 14648 20460
rect 14700 20408 14706 20460
rect 15286 20408 15292 20460
rect 15344 20448 15350 20460
rect 15473 20451 15531 20457
rect 15473 20448 15485 20451
rect 15344 20420 15485 20448
rect 15344 20408 15350 20420
rect 15473 20417 15485 20420
rect 15519 20417 15531 20451
rect 15473 20411 15531 20417
rect 16301 20451 16359 20457
rect 16301 20417 16313 20451
rect 16347 20417 16359 20451
rect 16301 20411 16359 20417
rect 14458 20272 14464 20324
rect 14516 20272 14522 20324
rect 16316 20312 16344 20411
rect 16942 20408 16948 20460
rect 17000 20446 17006 20460
rect 17037 20451 17095 20457
rect 17037 20446 17049 20451
rect 17000 20418 17049 20446
rect 17000 20408 17006 20418
rect 17037 20417 17049 20418
rect 17083 20417 17095 20451
rect 17037 20411 17095 20417
rect 16390 20340 16396 20392
rect 16448 20380 16454 20392
rect 17221 20383 17279 20389
rect 17221 20380 17233 20383
rect 16448 20352 17233 20380
rect 16448 20340 16454 20352
rect 17221 20349 17233 20352
rect 17267 20349 17279 20383
rect 17696 20380 17724 20556
rect 17770 20544 17776 20596
rect 17828 20544 17834 20596
rect 18690 20544 18696 20596
rect 18748 20544 18754 20596
rect 19705 20587 19763 20593
rect 19705 20553 19717 20587
rect 19751 20553 19763 20587
rect 19705 20547 19763 20553
rect 17957 20451 18015 20457
rect 17957 20417 17969 20451
rect 18003 20448 18015 20451
rect 18782 20448 18788 20460
rect 18003 20420 18788 20448
rect 18003 20417 18015 20420
rect 17957 20411 18015 20417
rect 18782 20408 18788 20420
rect 18840 20408 18846 20460
rect 18877 20451 18935 20457
rect 18877 20417 18889 20451
rect 18923 20448 18935 20451
rect 19720 20448 19748 20547
rect 20070 20544 20076 20596
rect 20128 20544 20134 20596
rect 20162 20544 20168 20596
rect 20220 20584 20226 20596
rect 22005 20587 22063 20593
rect 22005 20584 22017 20587
rect 20220 20556 22017 20584
rect 20220 20544 20226 20556
rect 22005 20553 22017 20556
rect 22051 20553 22063 20587
rect 22005 20547 22063 20553
rect 22186 20544 22192 20596
rect 22244 20584 22250 20596
rect 22244 20556 24808 20584
rect 22244 20544 22250 20556
rect 19978 20476 19984 20528
rect 20036 20516 20042 20528
rect 20036 20488 22232 20516
rect 20036 20476 20042 20488
rect 18923 20420 19748 20448
rect 18923 20417 18935 20420
rect 18877 20411 18935 20417
rect 19794 20408 19800 20460
rect 19852 20448 19858 20460
rect 21082 20448 21088 20460
rect 19852 20420 21088 20448
rect 19852 20408 19858 20420
rect 21082 20408 21088 20420
rect 21140 20408 21146 20460
rect 22204 20457 22232 20488
rect 22189 20451 22247 20457
rect 22189 20417 22201 20451
rect 22235 20417 22247 20451
rect 22189 20411 22247 20417
rect 22922 20408 22928 20460
rect 22980 20448 22986 20460
rect 23385 20451 23443 20457
rect 22980 20420 23336 20448
rect 22980 20408 22986 20420
rect 19518 20380 19524 20392
rect 17696 20352 19524 20380
rect 17221 20343 17279 20349
rect 19518 20340 19524 20352
rect 19576 20380 19582 20392
rect 20165 20383 20223 20389
rect 20165 20380 20177 20383
rect 19576 20352 20177 20380
rect 19576 20340 19582 20352
rect 20165 20349 20177 20352
rect 20211 20349 20223 20383
rect 20165 20343 20223 20349
rect 20257 20383 20315 20389
rect 20257 20349 20269 20383
rect 20303 20349 20315 20383
rect 20257 20343 20315 20349
rect 23201 20383 23259 20389
rect 23201 20349 23213 20383
rect 23247 20349 23259 20383
rect 23308 20380 23336 20420
rect 23385 20417 23397 20451
rect 23431 20448 23443 20451
rect 24578 20448 24584 20460
rect 23431 20420 24584 20448
rect 23431 20417 23443 20420
rect 23385 20411 23443 20417
rect 24578 20408 24584 20420
rect 24636 20408 24642 20460
rect 24780 20457 24808 20556
rect 24854 20544 24860 20596
rect 24912 20584 24918 20596
rect 31665 20587 31723 20593
rect 31665 20584 31677 20587
rect 24912 20556 31677 20584
rect 24912 20544 24918 20556
rect 31665 20553 31677 20556
rect 31711 20553 31723 20587
rect 31665 20547 31723 20553
rect 27433 20519 27491 20525
rect 27433 20516 27445 20519
rect 26206 20488 27445 20516
rect 24765 20451 24823 20457
rect 24765 20417 24777 20451
rect 24811 20417 24823 20451
rect 24765 20411 24823 20417
rect 25409 20451 25467 20457
rect 25409 20417 25421 20451
rect 25455 20417 25467 20451
rect 25409 20411 25467 20417
rect 25424 20380 25452 20411
rect 26050 20408 26056 20460
rect 26108 20408 26114 20460
rect 23308 20352 25452 20380
rect 23201 20343 23259 20349
rect 19794 20312 19800 20324
rect 16316 20284 19800 20312
rect 19794 20272 19800 20284
rect 19852 20272 19858 20324
rect 19886 20272 19892 20324
rect 19944 20312 19950 20324
rect 20272 20312 20300 20343
rect 20901 20315 20959 20321
rect 20901 20312 20913 20315
rect 19944 20284 20913 20312
rect 19944 20272 19950 20284
rect 20901 20281 20913 20284
rect 20947 20281 20959 20315
rect 20901 20275 20959 20281
rect 21082 20272 21088 20324
rect 21140 20312 21146 20324
rect 23216 20312 23244 20343
rect 25590 20340 25596 20392
rect 25648 20380 25654 20392
rect 26206 20380 26234 20488
rect 27433 20485 27445 20488
rect 27479 20485 27491 20519
rect 28718 20516 28724 20528
rect 28658 20488 28724 20516
rect 27433 20479 27491 20485
rect 28718 20476 28724 20488
rect 28776 20476 28782 20528
rect 30190 20476 30196 20528
rect 30248 20476 30254 20528
rect 30742 20476 30748 20528
rect 30800 20476 30806 20528
rect 25648 20352 26234 20380
rect 25648 20340 25654 20352
rect 26510 20340 26516 20392
rect 26568 20380 26574 20392
rect 27157 20383 27215 20389
rect 27157 20380 27169 20383
rect 26568 20352 27169 20380
rect 26568 20340 26574 20352
rect 27157 20349 27169 20352
rect 27203 20349 27215 20383
rect 27157 20343 27215 20349
rect 29914 20340 29920 20392
rect 29972 20340 29978 20392
rect 23382 20312 23388 20324
rect 21140 20284 22094 20312
rect 23216 20284 23388 20312
rect 21140 20272 21146 20284
rect 14642 20204 14648 20256
rect 14700 20244 14706 20256
rect 16117 20247 16175 20253
rect 16117 20244 16129 20247
rect 14700 20216 16129 20244
rect 14700 20204 14706 20216
rect 16117 20213 16129 20216
rect 16163 20213 16175 20247
rect 16117 20207 16175 20213
rect 16206 20204 16212 20256
rect 16264 20244 16270 20256
rect 16853 20247 16911 20253
rect 16853 20244 16865 20247
rect 16264 20216 16865 20244
rect 16264 20204 16270 20216
rect 16853 20213 16865 20216
rect 16899 20213 16911 20247
rect 16853 20207 16911 20213
rect 17034 20204 17040 20256
rect 17092 20244 17098 20256
rect 20162 20244 20168 20256
rect 17092 20216 20168 20244
rect 17092 20204 17098 20216
rect 20162 20204 20168 20216
rect 20220 20204 20226 20256
rect 22066 20244 22094 20284
rect 23382 20272 23388 20284
rect 23440 20272 23446 20324
rect 24581 20315 24639 20321
rect 24581 20312 24593 20315
rect 23492 20284 24593 20312
rect 23492 20244 23520 20284
rect 24581 20281 24593 20284
rect 24627 20281 24639 20315
rect 25869 20315 25927 20321
rect 25869 20312 25881 20315
rect 24581 20275 24639 20281
rect 24688 20284 25881 20312
rect 22066 20216 23520 20244
rect 23569 20247 23627 20253
rect 23569 20213 23581 20247
rect 23615 20244 23627 20247
rect 24394 20244 24400 20256
rect 23615 20216 24400 20244
rect 23615 20213 23627 20216
rect 23569 20207 23627 20213
rect 24394 20204 24400 20216
rect 24452 20204 24458 20256
rect 24486 20204 24492 20256
rect 24544 20244 24550 20256
rect 24688 20244 24716 20284
rect 25869 20281 25881 20284
rect 25915 20281 25927 20315
rect 25869 20275 25927 20281
rect 24544 20216 24716 20244
rect 24544 20204 24550 20216
rect 24854 20204 24860 20256
rect 24912 20244 24918 20256
rect 25225 20247 25283 20253
rect 25225 20244 25237 20247
rect 24912 20216 25237 20244
rect 24912 20204 24918 20216
rect 25225 20213 25237 20216
rect 25271 20213 25283 20247
rect 25225 20207 25283 20213
rect 25314 20204 25320 20256
rect 25372 20244 25378 20256
rect 28905 20247 28963 20253
rect 28905 20244 28917 20247
rect 25372 20216 28917 20244
rect 25372 20204 25378 20216
rect 28905 20213 28917 20216
rect 28951 20213 28963 20247
rect 28905 20207 28963 20213
rect 1104 20154 32476 20176
rect 1104 20102 4871 20154
rect 4923 20102 4935 20154
rect 4987 20102 4999 20154
rect 5051 20102 5063 20154
rect 5115 20102 5127 20154
rect 5179 20102 12713 20154
rect 12765 20102 12777 20154
rect 12829 20102 12841 20154
rect 12893 20102 12905 20154
rect 12957 20102 12969 20154
rect 13021 20102 20555 20154
rect 20607 20102 20619 20154
rect 20671 20102 20683 20154
rect 20735 20102 20747 20154
rect 20799 20102 20811 20154
rect 20863 20102 28397 20154
rect 28449 20102 28461 20154
rect 28513 20102 28525 20154
rect 28577 20102 28589 20154
rect 28641 20102 28653 20154
rect 28705 20102 32476 20154
rect 1104 20080 32476 20102
rect 2222 20000 2228 20052
rect 2280 20000 2286 20052
rect 3050 20000 3056 20052
rect 3108 20000 3114 20052
rect 4338 20000 4344 20052
rect 4396 20000 4402 20052
rect 5077 20043 5135 20049
rect 5077 20009 5089 20043
rect 5123 20040 5135 20043
rect 5258 20040 5264 20052
rect 5123 20012 5264 20040
rect 5123 20009 5135 20012
rect 5077 20003 5135 20009
rect 5258 20000 5264 20012
rect 5316 20000 5322 20052
rect 5810 20000 5816 20052
rect 5868 20000 5874 20052
rect 6546 20000 6552 20052
rect 6604 20000 6610 20052
rect 9122 20000 9128 20052
rect 9180 20040 9186 20052
rect 10505 20043 10563 20049
rect 10505 20040 10517 20043
rect 9180 20012 10517 20040
rect 9180 20000 9186 20012
rect 10505 20009 10517 20012
rect 10551 20009 10563 20043
rect 10505 20003 10563 20009
rect 11054 20000 11060 20052
rect 11112 20040 11118 20052
rect 11241 20043 11299 20049
rect 11241 20040 11253 20043
rect 11112 20012 11253 20040
rect 11112 20000 11118 20012
rect 11241 20009 11253 20012
rect 11287 20009 11299 20043
rect 11241 20003 11299 20009
rect 13541 20043 13599 20049
rect 13541 20009 13553 20043
rect 13587 20040 13599 20043
rect 13722 20040 13728 20052
rect 13587 20012 13728 20040
rect 13587 20009 13599 20012
rect 13541 20003 13599 20009
rect 13722 20000 13728 20012
rect 13780 20000 13786 20052
rect 14366 20000 14372 20052
rect 14424 20000 14430 20052
rect 15286 20000 15292 20052
rect 15344 20000 15350 20052
rect 16022 20000 16028 20052
rect 16080 20040 16086 20052
rect 16080 20012 18828 20040
rect 16080 20000 16086 20012
rect 14642 19972 14648 19984
rect 6886 19944 14648 19972
rect 6886 19904 6914 19944
rect 14642 19932 14648 19944
rect 14700 19972 14706 19984
rect 18800 19972 18828 20012
rect 18874 20000 18880 20052
rect 18932 20000 18938 20052
rect 24486 20040 24492 20052
rect 19812 20012 24492 20040
rect 19610 19972 19616 19984
rect 14700 19944 16620 19972
rect 18800 19944 19616 19972
rect 14700 19932 14706 19944
rect 6380 19876 6914 19904
rect 2409 19839 2467 19845
rect 2409 19805 2421 19839
rect 2455 19836 2467 19839
rect 2869 19839 2927 19845
rect 2869 19836 2881 19839
rect 2455 19808 2881 19836
rect 2455 19805 2467 19808
rect 2409 19799 2467 19805
rect 2869 19805 2881 19808
rect 2915 19836 2927 19839
rect 4062 19836 4068 19848
rect 2915 19808 4068 19836
rect 2915 19805 2927 19808
rect 2869 19799 2927 19805
rect 4062 19796 4068 19808
rect 4120 19836 4126 19848
rect 6380 19845 6408 19876
rect 11054 19864 11060 19916
rect 11112 19904 11118 19916
rect 12161 19907 12219 19913
rect 12161 19904 12173 19907
rect 11112 19876 12173 19904
rect 11112 19864 11118 19876
rect 12161 19873 12173 19876
rect 12207 19873 12219 19907
rect 12161 19867 12219 19873
rect 14458 19864 14464 19916
rect 14516 19904 14522 19916
rect 14737 19907 14795 19913
rect 14737 19904 14749 19907
rect 14516 19876 14749 19904
rect 14516 19864 14522 19876
rect 14737 19873 14749 19876
rect 14783 19904 14795 19907
rect 15470 19904 15476 19916
rect 14783 19876 15476 19904
rect 14783 19873 14795 19876
rect 14737 19867 14795 19873
rect 15470 19864 15476 19876
rect 15528 19904 15534 19916
rect 15933 19907 15991 19913
rect 15933 19904 15945 19907
rect 15528 19876 15945 19904
rect 15528 19864 15534 19876
rect 15933 19873 15945 19876
rect 15979 19904 15991 19907
rect 16390 19904 16396 19916
rect 15979 19876 16396 19904
rect 15979 19873 15991 19876
rect 15933 19867 15991 19873
rect 16390 19864 16396 19876
rect 16448 19864 16454 19916
rect 16592 19913 16620 19944
rect 19610 19932 19616 19944
rect 19668 19932 19674 19984
rect 16577 19907 16635 19913
rect 16577 19873 16589 19907
rect 16623 19873 16635 19907
rect 16577 19867 16635 19873
rect 16761 19907 16819 19913
rect 16761 19873 16773 19907
rect 16807 19904 16819 19907
rect 16942 19904 16948 19916
rect 16807 19876 16948 19904
rect 16807 19873 16819 19876
rect 16761 19867 16819 19873
rect 16942 19864 16948 19876
rect 17000 19904 17006 19916
rect 18601 19907 18659 19913
rect 17000 19876 18552 19904
rect 17000 19864 17006 19876
rect 18524 19848 18552 19876
rect 18601 19873 18613 19907
rect 18647 19873 18659 19907
rect 18601 19867 18659 19873
rect 4157 19839 4215 19845
rect 4157 19836 4169 19839
rect 4120 19808 4169 19836
rect 4120 19796 4126 19808
rect 4157 19805 4169 19808
rect 4203 19836 4215 19839
rect 4893 19839 4951 19845
rect 4893 19836 4905 19839
rect 4203 19808 4905 19836
rect 4203 19805 4215 19808
rect 4157 19799 4215 19805
rect 4893 19805 4905 19808
rect 4939 19836 4951 19839
rect 5629 19839 5687 19845
rect 5629 19836 5641 19839
rect 4939 19808 5641 19836
rect 4939 19805 4951 19808
rect 4893 19799 4951 19805
rect 5629 19805 5641 19808
rect 5675 19836 5687 19839
rect 6365 19839 6423 19845
rect 6365 19836 6377 19839
rect 5675 19808 6377 19836
rect 5675 19805 5687 19808
rect 5629 19799 5687 19805
rect 6365 19805 6377 19808
rect 6411 19805 6423 19839
rect 6365 19799 6423 19805
rect 10689 19839 10747 19845
rect 10689 19805 10701 19839
rect 10735 19836 10747 19839
rect 13170 19836 13176 19848
rect 10735 19808 13176 19836
rect 10735 19805 10747 19808
rect 10689 19799 10747 19805
rect 13170 19796 13176 19808
rect 13228 19796 13234 19848
rect 13722 19796 13728 19848
rect 13780 19796 13786 19848
rect 14553 19839 14611 19845
rect 14553 19805 14565 19839
rect 14599 19836 14611 19839
rect 15562 19836 15568 19848
rect 14599 19808 15568 19836
rect 14599 19805 14611 19808
rect 14553 19799 14611 19805
rect 15562 19796 15568 19808
rect 15620 19796 15626 19848
rect 15657 19839 15715 19845
rect 15657 19805 15669 19839
rect 15703 19836 15715 19839
rect 15703 19808 17816 19836
rect 15703 19805 15715 19808
rect 15657 19799 15715 19805
rect 11517 19771 11575 19777
rect 11517 19737 11529 19771
rect 11563 19768 11575 19771
rect 12437 19771 12495 19777
rect 11563 19740 12388 19768
rect 11563 19737 11575 19740
rect 11517 19731 11575 19737
rect 12360 19700 12388 19740
rect 12437 19737 12449 19771
rect 12483 19768 12495 19771
rect 16206 19768 16212 19780
rect 12483 19740 16212 19768
rect 12483 19737 12495 19740
rect 12437 19731 12495 19737
rect 16206 19728 16212 19740
rect 16264 19728 16270 19780
rect 16853 19771 16911 19777
rect 16853 19737 16865 19771
rect 16899 19768 16911 19771
rect 17788 19768 17816 19808
rect 17862 19796 17868 19848
rect 17920 19796 17926 19848
rect 18506 19796 18512 19848
rect 18564 19796 18570 19848
rect 18616 19836 18644 19867
rect 19702 19836 19708 19848
rect 18616 19808 19708 19836
rect 19702 19796 19708 19808
rect 19760 19796 19766 19848
rect 19812 19845 19840 20012
rect 24486 20000 24492 20012
rect 24544 20000 24550 20052
rect 24578 20000 24584 20052
rect 24636 20000 24642 20052
rect 27430 20040 27436 20052
rect 26206 20012 27436 20040
rect 22557 19975 22615 19981
rect 22557 19941 22569 19975
rect 22603 19972 22615 19975
rect 23106 19972 23112 19984
rect 22603 19944 23112 19972
rect 22603 19941 22615 19944
rect 22557 19935 22615 19941
rect 23106 19932 23112 19944
rect 23164 19932 23170 19984
rect 23661 19975 23719 19981
rect 23661 19941 23673 19975
rect 23707 19972 23719 19975
rect 26206 19972 26234 20012
rect 27430 20000 27436 20012
rect 27488 20000 27494 20052
rect 23707 19944 26234 19972
rect 23707 19941 23719 19944
rect 23661 19935 23719 19941
rect 19886 19864 19892 19916
rect 19944 19904 19950 19916
rect 19981 19907 20039 19913
rect 19981 19904 19993 19907
rect 19944 19876 19993 19904
rect 19944 19864 19950 19876
rect 19981 19873 19993 19876
rect 20027 19904 20039 19907
rect 21177 19907 21235 19913
rect 21177 19904 21189 19907
rect 20027 19876 21189 19904
rect 20027 19873 20039 19876
rect 19981 19867 20039 19873
rect 21177 19873 21189 19876
rect 21223 19873 21235 19907
rect 21177 19867 21235 19873
rect 23382 19864 23388 19916
rect 23440 19864 23446 19916
rect 25958 19904 25964 19916
rect 23492 19876 25964 19904
rect 19797 19839 19855 19845
rect 19797 19805 19809 19839
rect 19843 19805 19855 19839
rect 19797 19799 19855 19805
rect 20993 19839 21051 19845
rect 20993 19805 21005 19839
rect 21039 19836 21051 19839
rect 21082 19836 21088 19848
rect 21039 19808 21088 19836
rect 21039 19805 21051 19808
rect 20993 19799 21051 19805
rect 21082 19796 21088 19808
rect 21140 19796 21146 19848
rect 23290 19796 23296 19848
rect 23348 19836 23354 19848
rect 23492 19836 23520 19876
rect 25958 19864 25964 19876
rect 26016 19864 26022 19916
rect 26145 19907 26203 19913
rect 26145 19873 26157 19907
rect 26191 19904 26203 19907
rect 26510 19904 26516 19916
rect 26191 19876 26516 19904
rect 26191 19873 26203 19876
rect 26145 19867 26203 19873
rect 26510 19864 26516 19876
rect 26568 19864 26574 19916
rect 26786 19864 26792 19916
rect 26844 19904 26850 19916
rect 29181 19907 29239 19913
rect 26844 19876 27660 19904
rect 26844 19864 26850 19876
rect 25409 19839 25467 19845
rect 25409 19836 25421 19839
rect 23348 19808 23520 19836
rect 24044 19808 25421 19836
rect 23348 19796 23354 19808
rect 16899 19740 17724 19768
rect 17788 19740 21036 19768
rect 16899 19737 16911 19740
rect 16853 19731 16911 19737
rect 13354 19700 13360 19712
rect 12360 19672 13360 19700
rect 13354 19660 13360 19672
rect 13412 19660 13418 19712
rect 15194 19660 15200 19712
rect 15252 19700 15258 19712
rect 15749 19703 15807 19709
rect 15749 19700 15761 19703
rect 15252 19672 15761 19700
rect 15252 19660 15258 19672
rect 15749 19669 15761 19672
rect 15795 19669 15807 19703
rect 15749 19663 15807 19669
rect 17221 19703 17279 19709
rect 17221 19669 17233 19703
rect 17267 19700 17279 19703
rect 17310 19700 17316 19712
rect 17267 19672 17316 19700
rect 17267 19669 17279 19672
rect 17221 19663 17279 19669
rect 17310 19660 17316 19672
rect 17368 19660 17374 19712
rect 17696 19709 17724 19740
rect 21008 19712 21036 19740
rect 22186 19728 22192 19780
rect 22244 19728 22250 19780
rect 17681 19703 17739 19709
rect 17681 19669 17693 19703
rect 17727 19669 17739 19703
rect 17681 19663 17739 19669
rect 18230 19660 18236 19712
rect 18288 19700 18294 19712
rect 19429 19703 19487 19709
rect 19429 19700 19441 19703
rect 18288 19672 19441 19700
rect 18288 19660 18294 19672
rect 19429 19669 19441 19672
rect 19475 19669 19487 19703
rect 19429 19663 19487 19669
rect 19610 19660 19616 19712
rect 19668 19700 19674 19712
rect 19794 19700 19800 19712
rect 19668 19672 19800 19700
rect 19668 19660 19674 19672
rect 19794 19660 19800 19672
rect 19852 19700 19858 19712
rect 19889 19703 19947 19709
rect 19889 19700 19901 19703
rect 19852 19672 19901 19700
rect 19852 19660 19858 19672
rect 19889 19669 19901 19672
rect 19935 19669 19947 19703
rect 19889 19663 19947 19669
rect 20622 19660 20628 19712
rect 20680 19660 20686 19712
rect 20990 19660 20996 19712
rect 21048 19660 21054 19712
rect 21085 19703 21143 19709
rect 21085 19669 21097 19703
rect 21131 19700 21143 19703
rect 21174 19700 21180 19712
rect 21131 19672 21180 19700
rect 21131 19669 21143 19672
rect 21085 19663 21143 19669
rect 21174 19660 21180 19672
rect 21232 19660 21238 19712
rect 22649 19703 22707 19709
rect 22649 19669 22661 19703
rect 22695 19700 22707 19703
rect 24044 19700 24072 19808
rect 25409 19805 25421 19808
rect 25455 19805 25467 19839
rect 25409 19799 25467 19805
rect 24118 19728 24124 19780
rect 24176 19768 24182 19780
rect 24765 19771 24823 19777
rect 24765 19768 24777 19771
rect 24176 19740 24777 19768
rect 24176 19728 24182 19740
rect 24765 19737 24777 19740
rect 24811 19737 24823 19771
rect 24765 19731 24823 19737
rect 24949 19771 25007 19777
rect 24949 19737 24961 19771
rect 24995 19737 25007 19771
rect 24949 19731 25007 19737
rect 22695 19672 24072 19700
rect 22695 19669 22707 19672
rect 22649 19663 22707 19669
rect 24302 19660 24308 19712
rect 24360 19700 24366 19712
rect 24964 19700 24992 19731
rect 25038 19728 25044 19780
rect 25096 19768 25102 19780
rect 26421 19771 26479 19777
rect 26421 19768 26433 19771
rect 25096 19740 26433 19768
rect 25096 19728 25102 19740
rect 26421 19737 26433 19740
rect 26467 19737 26479 19771
rect 27632 19768 27660 19876
rect 29181 19873 29193 19907
rect 29227 19904 29239 19907
rect 31662 19904 31668 19916
rect 29227 19876 31668 19904
rect 29227 19873 29239 19876
rect 29181 19867 29239 19873
rect 31662 19864 31668 19876
rect 31720 19864 31726 19916
rect 31481 19839 31539 19845
rect 31481 19805 31493 19839
rect 31527 19836 31539 19839
rect 31754 19836 31760 19848
rect 31527 19808 31760 19836
rect 31527 19805 31539 19808
rect 31481 19799 31539 19805
rect 31754 19796 31760 19808
rect 31812 19796 31818 19848
rect 27632 19754 28580 19768
rect 27646 19740 28580 19754
rect 26421 19731 26479 19737
rect 25314 19700 25320 19712
rect 24360 19672 25320 19700
rect 24360 19660 24366 19672
rect 25314 19660 25320 19672
rect 25372 19660 25378 19712
rect 25593 19703 25651 19709
rect 25593 19669 25605 19703
rect 25639 19700 25651 19703
rect 26234 19700 26240 19712
rect 25639 19672 26240 19700
rect 25639 19669 25651 19672
rect 25593 19663 25651 19669
rect 26234 19660 26240 19672
rect 26292 19660 26298 19712
rect 26326 19660 26332 19712
rect 26384 19700 26390 19712
rect 26786 19700 26792 19712
rect 26384 19672 26792 19700
rect 26384 19660 26390 19672
rect 26786 19660 26792 19672
rect 26844 19660 26850 19712
rect 27062 19660 27068 19712
rect 27120 19700 27126 19712
rect 28552 19709 28580 19740
rect 27893 19703 27951 19709
rect 27893 19700 27905 19703
rect 27120 19672 27905 19700
rect 27120 19660 27126 19672
rect 27893 19669 27905 19672
rect 27939 19669 27951 19703
rect 27893 19663 27951 19669
rect 28537 19703 28595 19709
rect 28537 19669 28549 19703
rect 28583 19700 28595 19703
rect 28718 19700 28724 19712
rect 28583 19672 28724 19700
rect 28583 19669 28595 19672
rect 28537 19663 28595 19669
rect 28718 19660 28724 19672
rect 28776 19660 28782 19712
rect 30190 19660 30196 19712
rect 30248 19660 30254 19712
rect 1104 19610 32632 19632
rect 1104 19558 8792 19610
rect 8844 19558 8856 19610
rect 8908 19558 8920 19610
rect 8972 19558 8984 19610
rect 9036 19558 9048 19610
rect 9100 19558 16634 19610
rect 16686 19558 16698 19610
rect 16750 19558 16762 19610
rect 16814 19558 16826 19610
rect 16878 19558 16890 19610
rect 16942 19558 24476 19610
rect 24528 19558 24540 19610
rect 24592 19558 24604 19610
rect 24656 19558 24668 19610
rect 24720 19558 24732 19610
rect 24784 19558 32318 19610
rect 32370 19558 32382 19610
rect 32434 19558 32446 19610
rect 32498 19558 32510 19610
rect 32562 19558 32574 19610
rect 32626 19558 32632 19610
rect 1104 19536 32632 19558
rect 2406 19456 2412 19508
rect 2464 19456 2470 19508
rect 3878 19456 3884 19508
rect 3936 19456 3942 19508
rect 10962 19456 10968 19508
rect 11020 19456 11026 19508
rect 11882 19456 11888 19508
rect 11940 19496 11946 19508
rect 12437 19499 12495 19505
rect 12437 19496 12449 19499
rect 11940 19468 12449 19496
rect 11940 19456 11946 19468
rect 12437 19465 12449 19468
rect 12483 19465 12495 19499
rect 12437 19459 12495 19465
rect 13170 19456 13176 19508
rect 13228 19456 13234 19508
rect 13280 19468 13584 19496
rect 13280 19428 13308 19468
rect 13446 19428 13452 19440
rect 12636 19400 13308 19428
rect 13372 19400 13452 19428
rect 2593 19363 2651 19369
rect 2593 19329 2605 19363
rect 2639 19360 2651 19363
rect 4062 19360 4068 19372
rect 2639 19332 4068 19360
rect 2639 19329 2651 19332
rect 2593 19323 2651 19329
rect 4062 19320 4068 19332
rect 4120 19320 4126 19372
rect 11146 19320 11152 19372
rect 11204 19320 11210 19372
rect 12636 19369 12664 19400
rect 13372 19369 13400 19400
rect 13446 19388 13452 19400
rect 13504 19388 13510 19440
rect 13556 19428 13584 19468
rect 13722 19456 13728 19508
rect 13780 19496 13786 19508
rect 14829 19499 14887 19505
rect 14829 19496 14841 19499
rect 13780 19468 14841 19496
rect 13780 19456 13786 19468
rect 14829 19465 14841 19468
rect 14875 19465 14887 19499
rect 16022 19496 16028 19508
rect 14829 19459 14887 19465
rect 15120 19468 16028 19496
rect 14001 19431 14059 19437
rect 14001 19428 14013 19431
rect 13556 19400 14013 19428
rect 14001 19397 14013 19400
rect 14047 19397 14059 19431
rect 15120 19428 15148 19468
rect 16022 19456 16028 19468
rect 16080 19456 16086 19508
rect 16114 19456 16120 19508
rect 16172 19456 16178 19508
rect 17954 19456 17960 19508
rect 18012 19496 18018 19508
rect 20441 19499 20499 19505
rect 20441 19496 20453 19499
rect 18012 19468 20453 19496
rect 18012 19456 18018 19468
rect 20441 19465 20453 19468
rect 20487 19465 20499 19499
rect 20441 19459 20499 19465
rect 20809 19499 20867 19505
rect 20809 19465 20821 19499
rect 20855 19496 20867 19499
rect 22005 19499 22063 19505
rect 22005 19496 22017 19499
rect 20855 19468 22017 19496
rect 20855 19465 20867 19468
rect 20809 19459 20867 19465
rect 22005 19465 22017 19468
rect 22051 19465 22063 19499
rect 22005 19459 22063 19465
rect 23106 19456 23112 19508
rect 23164 19456 23170 19508
rect 23382 19456 23388 19508
rect 23440 19496 23446 19508
rect 24121 19499 24179 19505
rect 24121 19496 24133 19499
rect 23440 19468 24133 19496
rect 23440 19456 23446 19468
rect 24121 19465 24133 19468
rect 24167 19465 24179 19499
rect 24121 19459 24179 19465
rect 24946 19456 24952 19508
rect 25004 19496 25010 19508
rect 27062 19496 27068 19508
rect 25004 19468 27068 19496
rect 25004 19456 25010 19468
rect 27062 19456 27068 19468
rect 27120 19456 27126 19508
rect 28905 19499 28963 19505
rect 28905 19496 28917 19499
rect 27356 19468 28917 19496
rect 14001 19391 14059 19397
rect 14200 19400 15148 19428
rect 15197 19431 15255 19437
rect 14200 19369 14228 19400
rect 15197 19397 15209 19431
rect 15243 19428 15255 19431
rect 17034 19428 17040 19440
rect 15243 19400 17040 19428
rect 15243 19397 15255 19400
rect 15197 19391 15255 19397
rect 17034 19388 17040 19400
rect 17092 19388 17098 19440
rect 17310 19388 17316 19440
rect 17368 19388 17374 19440
rect 19613 19431 19671 19437
rect 17696 19400 19380 19428
rect 12621 19363 12679 19369
rect 12621 19329 12633 19363
rect 12667 19329 12679 19363
rect 12621 19323 12679 19329
rect 13357 19363 13415 19369
rect 13357 19329 13369 19363
rect 13403 19329 13415 19363
rect 13357 19323 13415 19329
rect 14185 19363 14243 19369
rect 14185 19329 14197 19363
rect 14231 19329 14243 19363
rect 14185 19323 14243 19329
rect 14369 19363 14427 19369
rect 14369 19329 14381 19363
rect 14415 19360 14427 19363
rect 14458 19360 14464 19372
rect 14415 19332 14464 19360
rect 14415 19329 14427 19332
rect 14369 19323 14427 19329
rect 14458 19320 14464 19332
rect 14516 19320 14522 19372
rect 16301 19363 16359 19369
rect 16301 19329 16313 19363
rect 16347 19360 16359 19363
rect 17696 19360 17724 19400
rect 16347 19332 17724 19360
rect 16347 19329 16359 19332
rect 16301 19323 16359 19329
rect 17770 19320 17776 19372
rect 17828 19360 17834 19372
rect 17828 19332 18092 19360
rect 17828 19320 17834 19332
rect 13538 19252 13544 19304
rect 13596 19252 13602 19304
rect 15286 19252 15292 19304
rect 15344 19252 15350 19304
rect 15470 19252 15476 19304
rect 15528 19252 15534 19304
rect 13814 19184 13820 19236
rect 13872 19224 13878 19236
rect 18064 19233 18092 19332
rect 18230 19320 18236 19372
rect 18288 19320 18294 19372
rect 18782 19320 18788 19372
rect 18840 19360 18846 19372
rect 19352 19360 19380 19400
rect 19613 19397 19625 19431
rect 19659 19428 19671 19431
rect 24854 19428 24860 19440
rect 19659 19400 24860 19428
rect 19659 19397 19671 19400
rect 19613 19391 19671 19397
rect 24854 19388 24860 19400
rect 24912 19388 24918 19440
rect 26326 19428 26332 19440
rect 25898 19400 26332 19428
rect 26326 19388 26332 19400
rect 26384 19388 26390 19440
rect 26418 19388 26424 19440
rect 26476 19428 26482 19440
rect 27356 19428 27384 19468
rect 28905 19465 28917 19468
rect 28951 19465 28963 19499
rect 30742 19496 30748 19508
rect 28905 19459 28963 19465
rect 29012 19468 30748 19496
rect 26476 19400 27384 19428
rect 26476 19388 26482 19400
rect 27430 19388 27436 19440
rect 27488 19388 27494 19440
rect 28718 19428 28724 19440
rect 28658 19400 28724 19428
rect 28718 19388 28724 19400
rect 28776 19428 28782 19440
rect 29012 19428 29040 19468
rect 30742 19456 30748 19468
rect 30800 19456 30806 19508
rect 31478 19428 31484 19440
rect 28776 19400 29040 19428
rect 31234 19400 31484 19428
rect 28776 19388 28782 19400
rect 31478 19388 31484 19400
rect 31536 19388 31542 19440
rect 31662 19388 31668 19440
rect 31720 19428 31726 19440
rect 31757 19431 31815 19437
rect 31757 19428 31769 19431
rect 31720 19400 31769 19428
rect 31720 19388 31726 19400
rect 31757 19397 31769 19400
rect 31803 19397 31815 19431
rect 31757 19391 31815 19397
rect 20622 19360 20628 19372
rect 18840 19332 19288 19360
rect 19352 19332 20628 19360
rect 18840 19320 18846 19332
rect 19260 19233 19288 19332
rect 20622 19320 20628 19332
rect 20680 19320 20686 19372
rect 20901 19363 20959 19369
rect 20901 19329 20913 19363
rect 20947 19360 20959 19363
rect 21082 19360 21088 19372
rect 20947 19332 21088 19360
rect 20947 19329 20959 19332
rect 20901 19323 20959 19329
rect 21082 19320 21088 19332
rect 21140 19320 21146 19372
rect 21450 19320 21456 19372
rect 21508 19360 21514 19372
rect 22189 19363 22247 19369
rect 22189 19360 22201 19363
rect 21508 19332 22201 19360
rect 21508 19320 21514 19332
rect 22189 19329 22201 19332
rect 22235 19329 22247 19363
rect 22189 19323 22247 19329
rect 22296 19332 23612 19360
rect 19610 19252 19616 19304
rect 19668 19292 19674 19304
rect 19705 19295 19763 19301
rect 19705 19292 19717 19295
rect 19668 19264 19717 19292
rect 19668 19252 19674 19264
rect 19705 19261 19717 19264
rect 19751 19261 19763 19295
rect 19705 19255 19763 19261
rect 17037 19227 17095 19233
rect 17037 19224 17049 19227
rect 13872 19196 17049 19224
rect 13872 19184 13878 19196
rect 17037 19193 17049 19196
rect 17083 19193 17095 19227
rect 17037 19187 17095 19193
rect 18049 19227 18107 19233
rect 18049 19193 18061 19227
rect 18095 19193 18107 19227
rect 18049 19187 18107 19193
rect 19245 19227 19303 19233
rect 19245 19193 19257 19227
rect 19291 19193 19303 19227
rect 19245 19187 19303 19193
rect 19720 19156 19748 19255
rect 19886 19252 19892 19304
rect 19944 19252 19950 19304
rect 20993 19295 21051 19301
rect 20993 19261 21005 19295
rect 21039 19261 21051 19295
rect 20993 19255 21051 19261
rect 19904 19224 19932 19252
rect 21008 19224 21036 19255
rect 21174 19252 21180 19304
rect 21232 19292 21238 19304
rect 22296 19292 22324 19332
rect 21232 19264 22324 19292
rect 21232 19252 21238 19264
rect 23290 19252 23296 19304
rect 23348 19252 23354 19304
rect 23382 19252 23388 19304
rect 23440 19252 23446 19304
rect 23584 19301 23612 19332
rect 23658 19320 23664 19372
rect 23716 19360 23722 19372
rect 24118 19360 24124 19372
rect 23716 19332 24124 19360
rect 23716 19320 23722 19332
rect 24118 19320 24124 19332
rect 24176 19320 24182 19372
rect 24302 19320 24308 19372
rect 24360 19320 24366 19372
rect 23477 19295 23535 19301
rect 23477 19261 23489 19295
rect 23523 19261 23535 19295
rect 23477 19255 23535 19261
rect 23569 19295 23627 19301
rect 23569 19261 23581 19295
rect 23615 19292 23627 19295
rect 24857 19295 24915 19301
rect 24857 19292 24869 19295
rect 23615 19264 24869 19292
rect 23615 19261 23627 19264
rect 23569 19255 23627 19261
rect 24857 19261 24869 19264
rect 24903 19261 24915 19295
rect 24857 19255 24915 19261
rect 19904 19196 21036 19224
rect 23308 19156 23336 19252
rect 23492 19224 23520 19255
rect 26234 19252 26240 19304
rect 26292 19292 26298 19304
rect 26329 19295 26387 19301
rect 26329 19292 26341 19295
rect 26292 19264 26341 19292
rect 26292 19252 26298 19264
rect 26329 19261 26341 19264
rect 26375 19261 26387 19295
rect 26329 19255 26387 19261
rect 26605 19295 26663 19301
rect 26605 19261 26617 19295
rect 26651 19292 26663 19295
rect 27157 19295 27215 19301
rect 27157 19292 27169 19295
rect 26651 19264 27169 19292
rect 26651 19261 26663 19264
rect 26605 19255 26663 19261
rect 27157 19261 27169 19264
rect 27203 19261 27215 19295
rect 27157 19255 27215 19261
rect 29733 19295 29791 19301
rect 29733 19261 29745 19295
rect 29779 19292 29791 19295
rect 30009 19295 30067 19301
rect 29779 19264 29868 19292
rect 29779 19261 29791 19264
rect 29733 19255 29791 19261
rect 23658 19224 23664 19236
rect 23492 19196 23664 19224
rect 23658 19184 23664 19196
rect 23716 19184 23722 19236
rect 19720 19128 23336 19156
rect 23474 19116 23480 19168
rect 23532 19156 23538 19168
rect 24302 19156 24308 19168
rect 23532 19128 24308 19156
rect 23532 19116 23538 19128
rect 24302 19116 24308 19128
rect 24360 19116 24366 19168
rect 26326 19116 26332 19168
rect 26384 19156 26390 19168
rect 26510 19156 26516 19168
rect 26384 19128 26516 19156
rect 26384 19116 26390 19128
rect 26510 19116 26516 19128
rect 26568 19156 26574 19168
rect 26620 19156 26648 19255
rect 26568 19128 26648 19156
rect 29840 19156 29868 19264
rect 30009 19261 30021 19295
rect 30055 19292 30067 19295
rect 30098 19292 30104 19304
rect 30055 19264 30104 19292
rect 30055 19261 30067 19264
rect 30009 19255 30067 19261
rect 30098 19252 30104 19264
rect 30156 19252 30162 19304
rect 30006 19156 30012 19168
rect 29840 19128 30012 19156
rect 26568 19116 26574 19128
rect 30006 19116 30012 19128
rect 30064 19116 30070 19168
rect 1104 19066 32476 19088
rect 1104 19014 4871 19066
rect 4923 19014 4935 19066
rect 4987 19014 4999 19066
rect 5051 19014 5063 19066
rect 5115 19014 5127 19066
rect 5179 19014 12713 19066
rect 12765 19014 12777 19066
rect 12829 19014 12841 19066
rect 12893 19014 12905 19066
rect 12957 19014 12969 19066
rect 13021 19014 20555 19066
rect 20607 19014 20619 19066
rect 20671 19014 20683 19066
rect 20735 19014 20747 19066
rect 20799 19014 20811 19066
rect 20863 19014 28397 19066
rect 28449 19014 28461 19066
rect 28513 19014 28525 19066
rect 28577 19014 28589 19066
rect 28641 19014 28653 19066
rect 28705 19014 32476 19066
rect 1104 18992 32476 19014
rect 11054 18912 11060 18964
rect 11112 18952 11118 18964
rect 11517 18955 11575 18961
rect 11517 18952 11529 18955
rect 11112 18924 11529 18952
rect 11112 18912 11118 18924
rect 11517 18921 11529 18924
rect 11563 18921 11575 18955
rect 11517 18915 11575 18921
rect 13354 18912 13360 18964
rect 13412 18912 13418 18964
rect 15013 18955 15071 18961
rect 15013 18952 15025 18955
rect 13464 18924 15025 18952
rect 11146 18844 11152 18896
rect 11204 18884 11210 18896
rect 13464 18884 13492 18924
rect 15013 18921 15025 18924
rect 15059 18921 15071 18955
rect 15013 18915 15071 18921
rect 15838 18912 15844 18964
rect 15896 18912 15902 18964
rect 16574 18912 16580 18964
rect 16632 18952 16638 18964
rect 17129 18955 17187 18961
rect 17129 18952 17141 18955
rect 16632 18924 17141 18952
rect 16632 18912 16638 18924
rect 17129 18921 17141 18924
rect 17175 18921 17187 18955
rect 17129 18915 17187 18921
rect 19702 18912 19708 18964
rect 19760 18912 19766 18964
rect 20717 18955 20775 18961
rect 20717 18921 20729 18955
rect 20763 18952 20775 18955
rect 20990 18952 20996 18964
rect 20763 18924 20996 18952
rect 20763 18921 20775 18924
rect 20717 18915 20775 18921
rect 20990 18912 20996 18924
rect 21048 18912 21054 18964
rect 23017 18955 23075 18961
rect 23017 18921 23029 18955
rect 23063 18952 23075 18955
rect 30098 18952 30104 18964
rect 23063 18924 28304 18952
rect 23063 18921 23075 18924
rect 23017 18915 23075 18921
rect 11204 18856 13492 18884
rect 11204 18844 11210 18856
rect 13538 18844 13544 18896
rect 13596 18884 13602 18896
rect 15194 18884 15200 18896
rect 13596 18856 15200 18884
rect 13596 18844 13602 18856
rect 15194 18844 15200 18856
rect 15252 18884 15258 18896
rect 20254 18884 20260 18896
rect 15252 18856 20260 18884
rect 15252 18844 15258 18856
rect 20254 18844 20260 18856
rect 20312 18844 20318 18896
rect 21082 18844 21088 18896
rect 21140 18884 21146 18896
rect 22002 18884 22008 18896
rect 21140 18856 22008 18884
rect 21140 18844 21146 18856
rect 22002 18844 22008 18856
rect 22060 18884 22066 18896
rect 24029 18887 24087 18893
rect 22060 18856 23704 18884
rect 22060 18844 22066 18856
rect 15286 18816 15292 18828
rect 13556 18788 15292 18816
rect 11698 18708 11704 18760
rect 11756 18708 11762 18760
rect 13556 18757 13584 18788
rect 15286 18776 15292 18788
rect 15344 18816 15350 18828
rect 22741 18819 22799 18825
rect 15344 18788 22692 18816
rect 15344 18776 15350 18788
rect 13541 18751 13599 18757
rect 13541 18717 13553 18751
rect 13587 18717 13599 18751
rect 13541 18711 13599 18717
rect 13725 18751 13783 18757
rect 13725 18717 13737 18751
rect 13771 18748 13783 18751
rect 14458 18748 14464 18760
rect 13771 18720 14464 18748
rect 13771 18717 13783 18720
rect 13725 18711 13783 18717
rect 13446 18640 13452 18692
rect 13504 18680 13510 18692
rect 13740 18680 13768 18711
rect 14458 18708 14464 18720
rect 14516 18708 14522 18760
rect 15197 18751 15255 18757
rect 15197 18717 15209 18751
rect 15243 18717 15255 18751
rect 15197 18711 15255 18717
rect 15381 18751 15439 18757
rect 15381 18717 15393 18751
rect 15427 18748 15439 18751
rect 15470 18748 15476 18760
rect 15427 18720 15476 18748
rect 15427 18717 15439 18720
rect 15381 18711 15439 18717
rect 13504 18652 13768 18680
rect 13504 18640 13510 18652
rect 15212 18612 15240 18711
rect 15470 18708 15476 18720
rect 15528 18708 15534 18760
rect 16025 18751 16083 18757
rect 16025 18717 16037 18751
rect 16071 18717 16083 18751
rect 16025 18711 16083 18717
rect 16209 18751 16267 18757
rect 16209 18717 16221 18751
rect 16255 18748 16267 18751
rect 16390 18748 16396 18760
rect 16255 18720 16396 18748
rect 16255 18717 16267 18720
rect 16209 18711 16267 18717
rect 16040 18680 16068 18711
rect 16390 18708 16396 18720
rect 16448 18708 16454 18760
rect 17313 18751 17371 18757
rect 17313 18717 17325 18751
rect 17359 18748 17371 18751
rect 17954 18748 17960 18760
rect 17359 18720 17960 18748
rect 17359 18717 17371 18720
rect 17313 18711 17371 18717
rect 17954 18708 17960 18720
rect 18012 18708 18018 18760
rect 20088 18757 20116 18788
rect 20073 18751 20131 18757
rect 20073 18717 20085 18751
rect 20119 18717 20131 18751
rect 20073 18711 20131 18717
rect 20898 18708 20904 18760
rect 20956 18708 20962 18760
rect 22664 18757 22692 18788
rect 22741 18785 22753 18819
rect 22787 18816 22799 18819
rect 22830 18816 22836 18828
rect 22787 18788 22836 18816
rect 22787 18785 22799 18788
rect 22741 18779 22799 18785
rect 22830 18776 22836 18788
rect 22888 18816 22894 18828
rect 22888 18788 23336 18816
rect 22888 18776 22894 18788
rect 22649 18751 22707 18757
rect 22649 18717 22661 18751
rect 22695 18748 22707 18751
rect 22695 18720 23244 18748
rect 22695 18717 22707 18720
rect 22649 18711 22707 18717
rect 19702 18680 19708 18692
rect 16040 18652 19708 18680
rect 19702 18640 19708 18652
rect 19760 18640 19766 18692
rect 19981 18683 20039 18689
rect 19981 18680 19993 18683
rect 19812 18652 19993 18680
rect 19812 18612 19840 18652
rect 19981 18649 19993 18652
rect 20027 18649 20039 18683
rect 19981 18643 20039 18649
rect 15212 18584 19840 18612
rect 19886 18572 19892 18624
rect 19944 18572 19950 18624
rect 19996 18612 20024 18643
rect 20254 18640 20260 18692
rect 20312 18680 20318 18692
rect 23216 18680 23244 18720
rect 23308 18744 23336 18788
rect 23382 18776 23388 18828
rect 23440 18816 23446 18828
rect 23569 18819 23627 18825
rect 23569 18816 23581 18819
rect 23440 18788 23581 18816
rect 23440 18776 23446 18788
rect 23569 18785 23581 18788
rect 23615 18785 23627 18819
rect 23569 18779 23627 18785
rect 23676 18757 23704 18856
rect 24029 18853 24041 18887
rect 24075 18884 24087 18887
rect 25038 18884 25044 18896
rect 24075 18856 25044 18884
rect 24075 18853 24087 18856
rect 24029 18847 24087 18853
rect 25038 18844 25044 18856
rect 25096 18844 25102 18896
rect 25222 18844 25228 18896
rect 25280 18844 25286 18896
rect 24118 18776 24124 18828
rect 24176 18816 24182 18828
rect 24176 18788 24808 18816
rect 24176 18776 24182 18788
rect 23661 18751 23719 18757
rect 23308 18716 23428 18744
rect 23400 18680 23428 18716
rect 23661 18717 23673 18751
rect 23707 18748 23719 18751
rect 23750 18748 23756 18760
rect 23707 18720 23756 18748
rect 23707 18717 23719 18720
rect 23661 18711 23719 18717
rect 23750 18708 23756 18720
rect 23808 18708 23814 18760
rect 24780 18757 24808 18788
rect 25130 18776 25136 18828
rect 25188 18816 25194 18828
rect 25188 18788 28212 18816
rect 25188 18776 25194 18788
rect 24581 18751 24639 18757
rect 24581 18717 24593 18751
rect 24627 18717 24639 18751
rect 24581 18711 24639 18717
rect 24765 18751 24823 18757
rect 24765 18717 24777 18751
rect 24811 18717 24823 18751
rect 24765 18711 24823 18717
rect 24596 18680 24624 18711
rect 24854 18708 24860 18760
rect 24912 18748 24918 18760
rect 25409 18751 25467 18757
rect 25409 18748 25421 18751
rect 24912 18720 25421 18748
rect 24912 18708 24918 18720
rect 25409 18717 25421 18720
rect 25455 18717 25467 18751
rect 25409 18711 25467 18717
rect 26326 18708 26332 18760
rect 26384 18708 26390 18760
rect 27706 18708 27712 18760
rect 27764 18708 27770 18760
rect 20312 18652 22692 18680
rect 23216 18652 23336 18680
rect 23400 18652 24624 18680
rect 24673 18683 24731 18689
rect 20312 18640 20318 18652
rect 21082 18612 21088 18624
rect 19996 18584 21088 18612
rect 21082 18572 21088 18584
rect 21140 18572 21146 18624
rect 22664 18612 22692 18652
rect 23198 18612 23204 18624
rect 22664 18584 23204 18612
rect 23198 18572 23204 18584
rect 23256 18572 23262 18624
rect 23308 18612 23336 18652
rect 24673 18649 24685 18683
rect 24719 18680 24731 18683
rect 24719 18652 25452 18680
rect 24719 18649 24731 18652
rect 24673 18643 24731 18649
rect 25130 18612 25136 18624
rect 23308 18584 25136 18612
rect 25130 18572 25136 18584
rect 25188 18572 25194 18624
rect 25424 18612 25452 18652
rect 25498 18640 25504 18692
rect 25556 18680 25562 18692
rect 26605 18683 26663 18689
rect 26605 18680 26617 18683
rect 25556 18652 26617 18680
rect 25556 18640 25562 18652
rect 26605 18649 26617 18652
rect 26651 18649 26663 18683
rect 26605 18643 26663 18649
rect 27614 18612 27620 18624
rect 25424 18584 27620 18612
rect 27614 18572 27620 18584
rect 27672 18572 27678 18624
rect 28074 18572 28080 18624
rect 28132 18572 28138 18624
rect 28184 18612 28212 18788
rect 28276 18748 28304 18924
rect 29196 18924 30104 18952
rect 29196 18825 29224 18924
rect 30098 18912 30104 18924
rect 30156 18912 30162 18964
rect 29181 18819 29239 18825
rect 29181 18785 29193 18819
rect 29227 18785 29239 18819
rect 29181 18779 29239 18785
rect 28276 18720 29224 18748
rect 29196 18680 29224 18720
rect 30006 18708 30012 18760
rect 30064 18708 30070 18760
rect 30285 18683 30343 18689
rect 30285 18680 30297 18683
rect 29196 18652 30297 18680
rect 30285 18649 30297 18652
rect 30331 18649 30343 18683
rect 30285 18643 30343 18649
rect 30742 18640 30748 18692
rect 30800 18640 30806 18692
rect 31757 18615 31815 18621
rect 31757 18612 31769 18615
rect 28184 18584 31769 18612
rect 31757 18581 31769 18584
rect 31803 18581 31815 18615
rect 31757 18575 31815 18581
rect 1104 18522 32632 18544
rect 1104 18470 8792 18522
rect 8844 18470 8856 18522
rect 8908 18470 8920 18522
rect 8972 18470 8984 18522
rect 9036 18470 9048 18522
rect 9100 18470 16634 18522
rect 16686 18470 16698 18522
rect 16750 18470 16762 18522
rect 16814 18470 16826 18522
rect 16878 18470 16890 18522
rect 16942 18470 24476 18522
rect 24528 18470 24540 18522
rect 24592 18470 24604 18522
rect 24656 18470 24668 18522
rect 24720 18470 24732 18522
rect 24784 18470 32318 18522
rect 32370 18470 32382 18522
rect 32434 18470 32446 18522
rect 32498 18470 32510 18522
rect 32562 18470 32574 18522
rect 32626 18470 32632 18522
rect 1104 18448 32632 18470
rect 11698 18368 11704 18420
rect 11756 18408 11762 18420
rect 15657 18411 15715 18417
rect 15657 18408 15669 18411
rect 11756 18380 15669 18408
rect 11756 18368 11762 18380
rect 15657 18377 15669 18380
rect 15703 18377 15715 18411
rect 15657 18371 15715 18377
rect 19794 18368 19800 18420
rect 19852 18368 19858 18420
rect 19886 18368 19892 18420
rect 19944 18408 19950 18420
rect 19944 18380 20208 18408
rect 19944 18368 19950 18380
rect 19518 18300 19524 18352
rect 19576 18340 19582 18352
rect 19613 18343 19671 18349
rect 19613 18340 19625 18343
rect 19576 18312 19625 18340
rect 19576 18300 19582 18312
rect 19613 18309 19625 18312
rect 19659 18309 19671 18343
rect 19613 18303 19671 18309
rect 19702 18300 19708 18352
rect 19760 18340 19766 18352
rect 20180 18349 20208 18380
rect 22830 18368 22836 18420
rect 22888 18368 22894 18420
rect 23750 18368 23756 18420
rect 23808 18408 23814 18420
rect 24946 18408 24952 18420
rect 23808 18380 24952 18408
rect 23808 18368 23814 18380
rect 24946 18368 24952 18380
rect 25004 18368 25010 18420
rect 25133 18411 25191 18417
rect 25133 18377 25145 18411
rect 25179 18408 25191 18411
rect 25498 18408 25504 18420
rect 25179 18380 25504 18408
rect 25179 18377 25191 18380
rect 25133 18371 25191 18377
rect 25498 18368 25504 18380
rect 25556 18368 25562 18420
rect 27617 18411 27675 18417
rect 27617 18408 27629 18411
rect 26206 18380 27629 18408
rect 20165 18343 20223 18349
rect 19760 18312 19932 18340
rect 19760 18300 19766 18312
rect 15841 18275 15899 18281
rect 15841 18241 15853 18275
rect 15887 18241 15899 18275
rect 15841 18235 15899 18241
rect 16025 18275 16083 18281
rect 16025 18241 16037 18275
rect 16071 18272 16083 18275
rect 16390 18272 16396 18284
rect 16071 18244 16396 18272
rect 16071 18241 16083 18244
rect 16025 18235 16083 18241
rect 15856 18204 15884 18235
rect 16390 18232 16396 18244
rect 16448 18232 16454 18284
rect 19904 18281 19932 18312
rect 20165 18309 20177 18343
rect 20211 18340 20223 18343
rect 22186 18340 22192 18352
rect 20211 18312 22192 18340
rect 20211 18309 20223 18312
rect 20165 18303 20223 18309
rect 22186 18300 22192 18312
rect 22244 18340 22250 18352
rect 22985 18343 23043 18349
rect 22985 18340 22997 18343
rect 22244 18312 22997 18340
rect 22244 18300 22250 18312
rect 22985 18309 22997 18312
rect 23031 18340 23043 18343
rect 23031 18309 23060 18340
rect 22985 18303 23060 18309
rect 19889 18275 19947 18281
rect 19889 18241 19901 18275
rect 19935 18241 19947 18275
rect 19889 18235 19947 18241
rect 19981 18275 20039 18281
rect 19981 18241 19993 18275
rect 20027 18272 20039 18275
rect 21174 18272 21180 18284
rect 20027 18244 21180 18272
rect 20027 18241 20039 18244
rect 19981 18235 20039 18241
rect 19996 18204 20024 18235
rect 21174 18232 21180 18244
rect 21232 18232 21238 18284
rect 23032 18272 23060 18303
rect 23198 18300 23204 18352
rect 23256 18340 23262 18352
rect 23937 18343 23995 18349
rect 23937 18340 23949 18343
rect 23256 18312 23949 18340
rect 23256 18300 23262 18312
rect 23937 18309 23949 18312
rect 23983 18340 23995 18343
rect 26206 18340 26234 18380
rect 27617 18377 27629 18380
rect 27663 18377 27675 18411
rect 27617 18371 27675 18377
rect 27706 18368 27712 18420
rect 27764 18408 27770 18420
rect 28718 18408 28724 18420
rect 27764 18380 28724 18408
rect 27764 18368 27770 18380
rect 28718 18368 28724 18380
rect 28776 18368 28782 18420
rect 30006 18368 30012 18420
rect 30064 18408 30070 18420
rect 31297 18411 31355 18417
rect 31297 18408 31309 18411
rect 30064 18380 31309 18408
rect 30064 18368 30070 18380
rect 31297 18377 31309 18380
rect 31343 18377 31355 18411
rect 31297 18371 31355 18377
rect 28736 18340 28764 18368
rect 30024 18340 30052 18368
rect 23983 18312 26234 18340
rect 28658 18312 28764 18340
rect 29380 18312 30052 18340
rect 23983 18309 23995 18312
rect 23937 18303 23995 18309
rect 23382 18272 23388 18284
rect 23032 18244 23388 18272
rect 23382 18232 23388 18244
rect 23440 18272 23446 18284
rect 23661 18275 23719 18281
rect 23661 18272 23673 18275
rect 23440 18244 23673 18272
rect 23440 18232 23446 18244
rect 23661 18241 23673 18244
rect 23707 18241 23719 18275
rect 23661 18235 23719 18241
rect 24394 18232 24400 18284
rect 24452 18232 24458 18284
rect 29380 18281 29408 18312
rect 25041 18275 25099 18281
rect 25041 18241 25053 18275
rect 25087 18241 25099 18275
rect 25041 18235 25099 18241
rect 29365 18275 29423 18281
rect 29365 18241 29377 18275
rect 29411 18241 29423 18275
rect 29365 18235 29423 18241
rect 30009 18275 30067 18281
rect 30009 18241 30021 18275
rect 30055 18272 30067 18275
rect 30190 18272 30196 18284
rect 30055 18244 30196 18272
rect 30055 18241 30067 18244
rect 30009 18235 30067 18241
rect 23474 18204 23480 18216
rect 15856 18176 20024 18204
rect 20088 18176 23480 18204
rect 19794 18096 19800 18148
rect 19852 18136 19858 18148
rect 20088 18136 20116 18176
rect 23474 18164 23480 18176
rect 23532 18164 23538 18216
rect 25056 18204 25084 18235
rect 30190 18232 30196 18244
rect 30248 18232 30254 18284
rect 28074 18204 28080 18216
rect 23676 18176 28080 18204
rect 23676 18148 23704 18176
rect 28074 18164 28080 18176
rect 28132 18164 28138 18216
rect 23658 18136 23664 18148
rect 19852 18108 20116 18136
rect 20180 18108 23664 18136
rect 19852 18096 19858 18108
rect 19518 18028 19524 18080
rect 19576 18068 19582 18080
rect 20180 18068 20208 18108
rect 23658 18096 23664 18108
rect 23716 18096 23722 18148
rect 23937 18139 23995 18145
rect 23937 18105 23949 18139
rect 23983 18136 23995 18139
rect 24118 18136 24124 18148
rect 23983 18108 24124 18136
rect 23983 18105 23995 18108
rect 23937 18099 23995 18105
rect 24118 18096 24124 18108
rect 24176 18096 24182 18148
rect 24581 18139 24639 18145
rect 24581 18105 24593 18139
rect 24627 18136 24639 18139
rect 25590 18136 25596 18148
rect 24627 18108 25596 18136
rect 24627 18105 24639 18108
rect 24581 18099 24639 18105
rect 25590 18096 25596 18108
rect 25648 18096 25654 18148
rect 19576 18040 20208 18068
rect 19576 18028 19582 18040
rect 22002 18028 22008 18080
rect 22060 18068 22066 18080
rect 23017 18071 23075 18077
rect 23017 18068 23029 18071
rect 22060 18040 23029 18068
rect 22060 18028 22066 18040
rect 23017 18037 23029 18040
rect 23063 18037 23075 18071
rect 23017 18031 23075 18037
rect 27614 18028 27620 18080
rect 27672 18068 27678 18080
rect 29101 18071 29159 18077
rect 29101 18068 29113 18071
rect 27672 18040 29113 18068
rect 27672 18028 27678 18040
rect 29101 18037 29113 18040
rect 29147 18037 29159 18071
rect 29101 18031 29159 18037
rect 1104 17978 32476 18000
rect 1104 17926 4871 17978
rect 4923 17926 4935 17978
rect 4987 17926 4999 17978
rect 5051 17926 5063 17978
rect 5115 17926 5127 17978
rect 5179 17926 12713 17978
rect 12765 17926 12777 17978
rect 12829 17926 12841 17978
rect 12893 17926 12905 17978
rect 12957 17926 12969 17978
rect 13021 17926 20555 17978
rect 20607 17926 20619 17978
rect 20671 17926 20683 17978
rect 20735 17926 20747 17978
rect 20799 17926 20811 17978
rect 20863 17926 28397 17978
rect 28449 17926 28461 17978
rect 28513 17926 28525 17978
rect 28577 17926 28589 17978
rect 28641 17926 28653 17978
rect 28705 17926 32476 17978
rect 1104 17904 32476 17926
rect 26326 17824 26332 17876
rect 26384 17824 26390 17876
rect 30834 17824 30840 17876
rect 30892 17824 30898 17876
rect 31478 17824 31484 17876
rect 31536 17824 31542 17876
rect 27801 17663 27859 17669
rect 27801 17629 27813 17663
rect 27847 17660 27859 17663
rect 30190 17660 30196 17672
rect 27847 17632 30196 17660
rect 27847 17629 27859 17632
rect 27801 17623 27859 17629
rect 30190 17620 30196 17632
rect 30248 17620 30254 17672
rect 30282 17620 30288 17672
rect 30340 17660 30346 17672
rect 31021 17663 31079 17669
rect 31021 17660 31033 17663
rect 30340 17632 31033 17660
rect 30340 17620 30346 17632
rect 31021 17629 31033 17632
rect 31067 17629 31079 17663
rect 31021 17623 31079 17629
rect 31294 17620 31300 17672
rect 31352 17660 31358 17672
rect 31665 17663 31723 17669
rect 31665 17660 31677 17663
rect 31352 17632 31677 17660
rect 31352 17620 31358 17632
rect 31665 17629 31677 17632
rect 31711 17629 31723 17663
rect 31665 17623 31723 17629
rect 1104 17434 32632 17456
rect 1104 17382 8792 17434
rect 8844 17382 8856 17434
rect 8908 17382 8920 17434
rect 8972 17382 8984 17434
rect 9036 17382 9048 17434
rect 9100 17382 16634 17434
rect 16686 17382 16698 17434
rect 16750 17382 16762 17434
rect 16814 17382 16826 17434
rect 16878 17382 16890 17434
rect 16942 17382 24476 17434
rect 24528 17382 24540 17434
rect 24592 17382 24604 17434
rect 24656 17382 24668 17434
rect 24720 17382 24732 17434
rect 24784 17382 32318 17434
rect 32370 17382 32382 17434
rect 32434 17382 32446 17434
rect 32498 17382 32510 17434
rect 32562 17382 32574 17434
rect 32626 17382 32632 17434
rect 1104 17360 32632 17382
rect 1104 16890 32476 16912
rect 1104 16838 4871 16890
rect 4923 16838 4935 16890
rect 4987 16838 4999 16890
rect 5051 16838 5063 16890
rect 5115 16838 5127 16890
rect 5179 16838 12713 16890
rect 12765 16838 12777 16890
rect 12829 16838 12841 16890
rect 12893 16838 12905 16890
rect 12957 16838 12969 16890
rect 13021 16838 20555 16890
rect 20607 16838 20619 16890
rect 20671 16838 20683 16890
rect 20735 16838 20747 16890
rect 20799 16838 20811 16890
rect 20863 16838 28397 16890
rect 28449 16838 28461 16890
rect 28513 16838 28525 16890
rect 28577 16838 28589 16890
rect 28641 16838 28653 16890
rect 28705 16838 32476 16890
rect 1104 16816 32476 16838
rect 1104 16346 32632 16368
rect 1104 16294 8792 16346
rect 8844 16294 8856 16346
rect 8908 16294 8920 16346
rect 8972 16294 8984 16346
rect 9036 16294 9048 16346
rect 9100 16294 16634 16346
rect 16686 16294 16698 16346
rect 16750 16294 16762 16346
rect 16814 16294 16826 16346
rect 16878 16294 16890 16346
rect 16942 16294 24476 16346
rect 24528 16294 24540 16346
rect 24592 16294 24604 16346
rect 24656 16294 24668 16346
rect 24720 16294 24732 16346
rect 24784 16294 32318 16346
rect 32370 16294 32382 16346
rect 32434 16294 32446 16346
rect 32498 16294 32510 16346
rect 32562 16294 32574 16346
rect 32626 16294 32632 16346
rect 1104 16272 32632 16294
rect 1104 15802 32476 15824
rect 1104 15750 4871 15802
rect 4923 15750 4935 15802
rect 4987 15750 4999 15802
rect 5051 15750 5063 15802
rect 5115 15750 5127 15802
rect 5179 15750 12713 15802
rect 12765 15750 12777 15802
rect 12829 15750 12841 15802
rect 12893 15750 12905 15802
rect 12957 15750 12969 15802
rect 13021 15750 20555 15802
rect 20607 15750 20619 15802
rect 20671 15750 20683 15802
rect 20735 15750 20747 15802
rect 20799 15750 20811 15802
rect 20863 15750 28397 15802
rect 28449 15750 28461 15802
rect 28513 15750 28525 15802
rect 28577 15750 28589 15802
rect 28641 15750 28653 15802
rect 28705 15750 32476 15802
rect 1104 15728 32476 15750
rect 1104 15258 32632 15280
rect 1104 15206 8792 15258
rect 8844 15206 8856 15258
rect 8908 15206 8920 15258
rect 8972 15206 8984 15258
rect 9036 15206 9048 15258
rect 9100 15206 16634 15258
rect 16686 15206 16698 15258
rect 16750 15206 16762 15258
rect 16814 15206 16826 15258
rect 16878 15206 16890 15258
rect 16942 15206 24476 15258
rect 24528 15206 24540 15258
rect 24592 15206 24604 15258
rect 24656 15206 24668 15258
rect 24720 15206 24732 15258
rect 24784 15206 32318 15258
rect 32370 15206 32382 15258
rect 32434 15206 32446 15258
rect 32498 15206 32510 15258
rect 32562 15206 32574 15258
rect 32626 15206 32632 15258
rect 1104 15184 32632 15206
rect 1104 14714 32476 14736
rect 1104 14662 4871 14714
rect 4923 14662 4935 14714
rect 4987 14662 4999 14714
rect 5051 14662 5063 14714
rect 5115 14662 5127 14714
rect 5179 14662 12713 14714
rect 12765 14662 12777 14714
rect 12829 14662 12841 14714
rect 12893 14662 12905 14714
rect 12957 14662 12969 14714
rect 13021 14662 20555 14714
rect 20607 14662 20619 14714
rect 20671 14662 20683 14714
rect 20735 14662 20747 14714
rect 20799 14662 20811 14714
rect 20863 14662 28397 14714
rect 28449 14662 28461 14714
rect 28513 14662 28525 14714
rect 28577 14662 28589 14714
rect 28641 14662 28653 14714
rect 28705 14662 32476 14714
rect 1104 14640 32476 14662
rect 1104 14170 32632 14192
rect 1104 14118 8792 14170
rect 8844 14118 8856 14170
rect 8908 14118 8920 14170
rect 8972 14118 8984 14170
rect 9036 14118 9048 14170
rect 9100 14118 16634 14170
rect 16686 14118 16698 14170
rect 16750 14118 16762 14170
rect 16814 14118 16826 14170
rect 16878 14118 16890 14170
rect 16942 14118 24476 14170
rect 24528 14118 24540 14170
rect 24592 14118 24604 14170
rect 24656 14118 24668 14170
rect 24720 14118 24732 14170
rect 24784 14118 32318 14170
rect 32370 14118 32382 14170
rect 32434 14118 32446 14170
rect 32498 14118 32510 14170
rect 32562 14118 32574 14170
rect 32626 14118 32632 14170
rect 1104 14096 32632 14118
rect 1104 13626 32476 13648
rect 1104 13574 4871 13626
rect 4923 13574 4935 13626
rect 4987 13574 4999 13626
rect 5051 13574 5063 13626
rect 5115 13574 5127 13626
rect 5179 13574 12713 13626
rect 12765 13574 12777 13626
rect 12829 13574 12841 13626
rect 12893 13574 12905 13626
rect 12957 13574 12969 13626
rect 13021 13574 20555 13626
rect 20607 13574 20619 13626
rect 20671 13574 20683 13626
rect 20735 13574 20747 13626
rect 20799 13574 20811 13626
rect 20863 13574 28397 13626
rect 28449 13574 28461 13626
rect 28513 13574 28525 13626
rect 28577 13574 28589 13626
rect 28641 13574 28653 13626
rect 28705 13574 32476 13626
rect 1104 13552 32476 13574
rect 1104 13082 32632 13104
rect 1104 13030 8792 13082
rect 8844 13030 8856 13082
rect 8908 13030 8920 13082
rect 8972 13030 8984 13082
rect 9036 13030 9048 13082
rect 9100 13030 16634 13082
rect 16686 13030 16698 13082
rect 16750 13030 16762 13082
rect 16814 13030 16826 13082
rect 16878 13030 16890 13082
rect 16942 13030 24476 13082
rect 24528 13030 24540 13082
rect 24592 13030 24604 13082
rect 24656 13030 24668 13082
rect 24720 13030 24732 13082
rect 24784 13030 32318 13082
rect 32370 13030 32382 13082
rect 32434 13030 32446 13082
rect 32498 13030 32510 13082
rect 32562 13030 32574 13082
rect 32626 13030 32632 13082
rect 1104 13008 32632 13030
rect 1104 12538 32476 12560
rect 1104 12486 4871 12538
rect 4923 12486 4935 12538
rect 4987 12486 4999 12538
rect 5051 12486 5063 12538
rect 5115 12486 5127 12538
rect 5179 12486 12713 12538
rect 12765 12486 12777 12538
rect 12829 12486 12841 12538
rect 12893 12486 12905 12538
rect 12957 12486 12969 12538
rect 13021 12486 20555 12538
rect 20607 12486 20619 12538
rect 20671 12486 20683 12538
rect 20735 12486 20747 12538
rect 20799 12486 20811 12538
rect 20863 12486 28397 12538
rect 28449 12486 28461 12538
rect 28513 12486 28525 12538
rect 28577 12486 28589 12538
rect 28641 12486 28653 12538
rect 28705 12486 32476 12538
rect 1104 12464 32476 12486
rect 1104 11994 32632 12016
rect 1104 11942 8792 11994
rect 8844 11942 8856 11994
rect 8908 11942 8920 11994
rect 8972 11942 8984 11994
rect 9036 11942 9048 11994
rect 9100 11942 16634 11994
rect 16686 11942 16698 11994
rect 16750 11942 16762 11994
rect 16814 11942 16826 11994
rect 16878 11942 16890 11994
rect 16942 11942 24476 11994
rect 24528 11942 24540 11994
rect 24592 11942 24604 11994
rect 24656 11942 24668 11994
rect 24720 11942 24732 11994
rect 24784 11942 32318 11994
rect 32370 11942 32382 11994
rect 32434 11942 32446 11994
rect 32498 11942 32510 11994
rect 32562 11942 32574 11994
rect 32626 11942 32632 11994
rect 1104 11920 32632 11942
rect 1104 11450 32476 11472
rect 1104 11398 4871 11450
rect 4923 11398 4935 11450
rect 4987 11398 4999 11450
rect 5051 11398 5063 11450
rect 5115 11398 5127 11450
rect 5179 11398 12713 11450
rect 12765 11398 12777 11450
rect 12829 11398 12841 11450
rect 12893 11398 12905 11450
rect 12957 11398 12969 11450
rect 13021 11398 20555 11450
rect 20607 11398 20619 11450
rect 20671 11398 20683 11450
rect 20735 11398 20747 11450
rect 20799 11398 20811 11450
rect 20863 11398 28397 11450
rect 28449 11398 28461 11450
rect 28513 11398 28525 11450
rect 28577 11398 28589 11450
rect 28641 11398 28653 11450
rect 28705 11398 32476 11450
rect 1104 11376 32476 11398
rect 1104 10906 32632 10928
rect 1104 10854 8792 10906
rect 8844 10854 8856 10906
rect 8908 10854 8920 10906
rect 8972 10854 8984 10906
rect 9036 10854 9048 10906
rect 9100 10854 16634 10906
rect 16686 10854 16698 10906
rect 16750 10854 16762 10906
rect 16814 10854 16826 10906
rect 16878 10854 16890 10906
rect 16942 10854 24476 10906
rect 24528 10854 24540 10906
rect 24592 10854 24604 10906
rect 24656 10854 24668 10906
rect 24720 10854 24732 10906
rect 24784 10854 32318 10906
rect 32370 10854 32382 10906
rect 32434 10854 32446 10906
rect 32498 10854 32510 10906
rect 32562 10854 32574 10906
rect 32626 10854 32632 10906
rect 1104 10832 32632 10854
rect 1104 10362 32476 10384
rect 1104 10310 4871 10362
rect 4923 10310 4935 10362
rect 4987 10310 4999 10362
rect 5051 10310 5063 10362
rect 5115 10310 5127 10362
rect 5179 10310 12713 10362
rect 12765 10310 12777 10362
rect 12829 10310 12841 10362
rect 12893 10310 12905 10362
rect 12957 10310 12969 10362
rect 13021 10310 20555 10362
rect 20607 10310 20619 10362
rect 20671 10310 20683 10362
rect 20735 10310 20747 10362
rect 20799 10310 20811 10362
rect 20863 10310 28397 10362
rect 28449 10310 28461 10362
rect 28513 10310 28525 10362
rect 28577 10310 28589 10362
rect 28641 10310 28653 10362
rect 28705 10310 32476 10362
rect 1104 10288 32476 10310
rect 1104 9818 32632 9840
rect 1104 9766 8792 9818
rect 8844 9766 8856 9818
rect 8908 9766 8920 9818
rect 8972 9766 8984 9818
rect 9036 9766 9048 9818
rect 9100 9766 16634 9818
rect 16686 9766 16698 9818
rect 16750 9766 16762 9818
rect 16814 9766 16826 9818
rect 16878 9766 16890 9818
rect 16942 9766 24476 9818
rect 24528 9766 24540 9818
rect 24592 9766 24604 9818
rect 24656 9766 24668 9818
rect 24720 9766 24732 9818
rect 24784 9766 32318 9818
rect 32370 9766 32382 9818
rect 32434 9766 32446 9818
rect 32498 9766 32510 9818
rect 32562 9766 32574 9818
rect 32626 9766 32632 9818
rect 1104 9744 32632 9766
rect 1104 9274 32476 9296
rect 1104 9222 4871 9274
rect 4923 9222 4935 9274
rect 4987 9222 4999 9274
rect 5051 9222 5063 9274
rect 5115 9222 5127 9274
rect 5179 9222 12713 9274
rect 12765 9222 12777 9274
rect 12829 9222 12841 9274
rect 12893 9222 12905 9274
rect 12957 9222 12969 9274
rect 13021 9222 20555 9274
rect 20607 9222 20619 9274
rect 20671 9222 20683 9274
rect 20735 9222 20747 9274
rect 20799 9222 20811 9274
rect 20863 9222 28397 9274
rect 28449 9222 28461 9274
rect 28513 9222 28525 9274
rect 28577 9222 28589 9274
rect 28641 9222 28653 9274
rect 28705 9222 32476 9274
rect 1104 9200 32476 9222
rect 1104 8730 32632 8752
rect 1104 8678 8792 8730
rect 8844 8678 8856 8730
rect 8908 8678 8920 8730
rect 8972 8678 8984 8730
rect 9036 8678 9048 8730
rect 9100 8678 16634 8730
rect 16686 8678 16698 8730
rect 16750 8678 16762 8730
rect 16814 8678 16826 8730
rect 16878 8678 16890 8730
rect 16942 8678 24476 8730
rect 24528 8678 24540 8730
rect 24592 8678 24604 8730
rect 24656 8678 24668 8730
rect 24720 8678 24732 8730
rect 24784 8678 32318 8730
rect 32370 8678 32382 8730
rect 32434 8678 32446 8730
rect 32498 8678 32510 8730
rect 32562 8678 32574 8730
rect 32626 8678 32632 8730
rect 1104 8656 32632 8678
rect 1104 8186 32476 8208
rect 1104 8134 4871 8186
rect 4923 8134 4935 8186
rect 4987 8134 4999 8186
rect 5051 8134 5063 8186
rect 5115 8134 5127 8186
rect 5179 8134 12713 8186
rect 12765 8134 12777 8186
rect 12829 8134 12841 8186
rect 12893 8134 12905 8186
rect 12957 8134 12969 8186
rect 13021 8134 20555 8186
rect 20607 8134 20619 8186
rect 20671 8134 20683 8186
rect 20735 8134 20747 8186
rect 20799 8134 20811 8186
rect 20863 8134 28397 8186
rect 28449 8134 28461 8186
rect 28513 8134 28525 8186
rect 28577 8134 28589 8186
rect 28641 8134 28653 8186
rect 28705 8134 32476 8186
rect 1104 8112 32476 8134
rect 1104 7642 32632 7664
rect 1104 7590 8792 7642
rect 8844 7590 8856 7642
rect 8908 7590 8920 7642
rect 8972 7590 8984 7642
rect 9036 7590 9048 7642
rect 9100 7590 16634 7642
rect 16686 7590 16698 7642
rect 16750 7590 16762 7642
rect 16814 7590 16826 7642
rect 16878 7590 16890 7642
rect 16942 7590 24476 7642
rect 24528 7590 24540 7642
rect 24592 7590 24604 7642
rect 24656 7590 24668 7642
rect 24720 7590 24732 7642
rect 24784 7590 32318 7642
rect 32370 7590 32382 7642
rect 32434 7590 32446 7642
rect 32498 7590 32510 7642
rect 32562 7590 32574 7642
rect 32626 7590 32632 7642
rect 1104 7568 32632 7590
rect 1104 7098 32476 7120
rect 1104 7046 4871 7098
rect 4923 7046 4935 7098
rect 4987 7046 4999 7098
rect 5051 7046 5063 7098
rect 5115 7046 5127 7098
rect 5179 7046 12713 7098
rect 12765 7046 12777 7098
rect 12829 7046 12841 7098
rect 12893 7046 12905 7098
rect 12957 7046 12969 7098
rect 13021 7046 20555 7098
rect 20607 7046 20619 7098
rect 20671 7046 20683 7098
rect 20735 7046 20747 7098
rect 20799 7046 20811 7098
rect 20863 7046 28397 7098
rect 28449 7046 28461 7098
rect 28513 7046 28525 7098
rect 28577 7046 28589 7098
rect 28641 7046 28653 7098
rect 28705 7046 32476 7098
rect 1104 7024 32476 7046
rect 1104 6554 32632 6576
rect 1104 6502 8792 6554
rect 8844 6502 8856 6554
rect 8908 6502 8920 6554
rect 8972 6502 8984 6554
rect 9036 6502 9048 6554
rect 9100 6502 16634 6554
rect 16686 6502 16698 6554
rect 16750 6502 16762 6554
rect 16814 6502 16826 6554
rect 16878 6502 16890 6554
rect 16942 6502 24476 6554
rect 24528 6502 24540 6554
rect 24592 6502 24604 6554
rect 24656 6502 24668 6554
rect 24720 6502 24732 6554
rect 24784 6502 32318 6554
rect 32370 6502 32382 6554
rect 32434 6502 32446 6554
rect 32498 6502 32510 6554
rect 32562 6502 32574 6554
rect 32626 6502 32632 6554
rect 1104 6480 32632 6502
rect 1104 6010 32476 6032
rect 1104 5958 4871 6010
rect 4923 5958 4935 6010
rect 4987 5958 4999 6010
rect 5051 5958 5063 6010
rect 5115 5958 5127 6010
rect 5179 5958 12713 6010
rect 12765 5958 12777 6010
rect 12829 5958 12841 6010
rect 12893 5958 12905 6010
rect 12957 5958 12969 6010
rect 13021 5958 20555 6010
rect 20607 5958 20619 6010
rect 20671 5958 20683 6010
rect 20735 5958 20747 6010
rect 20799 5958 20811 6010
rect 20863 5958 28397 6010
rect 28449 5958 28461 6010
rect 28513 5958 28525 6010
rect 28577 5958 28589 6010
rect 28641 5958 28653 6010
rect 28705 5958 32476 6010
rect 1104 5936 32476 5958
rect 1104 5466 32632 5488
rect 1104 5414 8792 5466
rect 8844 5414 8856 5466
rect 8908 5414 8920 5466
rect 8972 5414 8984 5466
rect 9036 5414 9048 5466
rect 9100 5414 16634 5466
rect 16686 5414 16698 5466
rect 16750 5414 16762 5466
rect 16814 5414 16826 5466
rect 16878 5414 16890 5466
rect 16942 5414 24476 5466
rect 24528 5414 24540 5466
rect 24592 5414 24604 5466
rect 24656 5414 24668 5466
rect 24720 5414 24732 5466
rect 24784 5414 32318 5466
rect 32370 5414 32382 5466
rect 32434 5414 32446 5466
rect 32498 5414 32510 5466
rect 32562 5414 32574 5466
rect 32626 5414 32632 5466
rect 1104 5392 32632 5414
rect 1104 4922 32476 4944
rect 1104 4870 4871 4922
rect 4923 4870 4935 4922
rect 4987 4870 4999 4922
rect 5051 4870 5063 4922
rect 5115 4870 5127 4922
rect 5179 4870 12713 4922
rect 12765 4870 12777 4922
rect 12829 4870 12841 4922
rect 12893 4870 12905 4922
rect 12957 4870 12969 4922
rect 13021 4870 20555 4922
rect 20607 4870 20619 4922
rect 20671 4870 20683 4922
rect 20735 4870 20747 4922
rect 20799 4870 20811 4922
rect 20863 4870 28397 4922
rect 28449 4870 28461 4922
rect 28513 4870 28525 4922
rect 28577 4870 28589 4922
rect 28641 4870 28653 4922
rect 28705 4870 32476 4922
rect 1104 4848 32476 4870
rect 1104 4378 32632 4400
rect 1104 4326 8792 4378
rect 8844 4326 8856 4378
rect 8908 4326 8920 4378
rect 8972 4326 8984 4378
rect 9036 4326 9048 4378
rect 9100 4326 16634 4378
rect 16686 4326 16698 4378
rect 16750 4326 16762 4378
rect 16814 4326 16826 4378
rect 16878 4326 16890 4378
rect 16942 4326 24476 4378
rect 24528 4326 24540 4378
rect 24592 4326 24604 4378
rect 24656 4326 24668 4378
rect 24720 4326 24732 4378
rect 24784 4326 32318 4378
rect 32370 4326 32382 4378
rect 32434 4326 32446 4378
rect 32498 4326 32510 4378
rect 32562 4326 32574 4378
rect 32626 4326 32632 4378
rect 1104 4304 32632 4326
rect 1104 3834 32476 3856
rect 1104 3782 4871 3834
rect 4923 3782 4935 3834
rect 4987 3782 4999 3834
rect 5051 3782 5063 3834
rect 5115 3782 5127 3834
rect 5179 3782 12713 3834
rect 12765 3782 12777 3834
rect 12829 3782 12841 3834
rect 12893 3782 12905 3834
rect 12957 3782 12969 3834
rect 13021 3782 20555 3834
rect 20607 3782 20619 3834
rect 20671 3782 20683 3834
rect 20735 3782 20747 3834
rect 20799 3782 20811 3834
rect 20863 3782 28397 3834
rect 28449 3782 28461 3834
rect 28513 3782 28525 3834
rect 28577 3782 28589 3834
rect 28641 3782 28653 3834
rect 28705 3782 32476 3834
rect 1104 3760 32476 3782
rect 1104 3290 32632 3312
rect 1104 3238 8792 3290
rect 8844 3238 8856 3290
rect 8908 3238 8920 3290
rect 8972 3238 8984 3290
rect 9036 3238 9048 3290
rect 9100 3238 16634 3290
rect 16686 3238 16698 3290
rect 16750 3238 16762 3290
rect 16814 3238 16826 3290
rect 16878 3238 16890 3290
rect 16942 3238 24476 3290
rect 24528 3238 24540 3290
rect 24592 3238 24604 3290
rect 24656 3238 24668 3290
rect 24720 3238 24732 3290
rect 24784 3238 32318 3290
rect 32370 3238 32382 3290
rect 32434 3238 32446 3290
rect 32498 3238 32510 3290
rect 32562 3238 32574 3290
rect 32626 3238 32632 3290
rect 1104 3216 32632 3238
rect 1104 2746 32476 2768
rect 1104 2694 4871 2746
rect 4923 2694 4935 2746
rect 4987 2694 4999 2746
rect 5051 2694 5063 2746
rect 5115 2694 5127 2746
rect 5179 2694 12713 2746
rect 12765 2694 12777 2746
rect 12829 2694 12841 2746
rect 12893 2694 12905 2746
rect 12957 2694 12969 2746
rect 13021 2694 20555 2746
rect 20607 2694 20619 2746
rect 20671 2694 20683 2746
rect 20735 2694 20747 2746
rect 20799 2694 20811 2746
rect 20863 2694 28397 2746
rect 28449 2694 28461 2746
rect 28513 2694 28525 2746
rect 28577 2694 28589 2746
rect 28641 2694 28653 2746
rect 28705 2694 32476 2746
rect 1104 2672 32476 2694
rect 1104 2202 32632 2224
rect 1104 2150 8792 2202
rect 8844 2150 8856 2202
rect 8908 2150 8920 2202
rect 8972 2150 8984 2202
rect 9036 2150 9048 2202
rect 9100 2150 16634 2202
rect 16686 2150 16698 2202
rect 16750 2150 16762 2202
rect 16814 2150 16826 2202
rect 16878 2150 16890 2202
rect 16942 2150 24476 2202
rect 24528 2150 24540 2202
rect 24592 2150 24604 2202
rect 24656 2150 24668 2202
rect 24720 2150 24732 2202
rect 24784 2150 32318 2202
rect 32370 2150 32382 2202
rect 32434 2150 32446 2202
rect 32498 2150 32510 2202
rect 32562 2150 32574 2202
rect 32626 2150 32632 2202
rect 1104 2128 32632 2150
rect 1104 1658 32476 1680
rect 1104 1606 4871 1658
rect 4923 1606 4935 1658
rect 4987 1606 4999 1658
rect 5051 1606 5063 1658
rect 5115 1606 5127 1658
rect 5179 1606 12713 1658
rect 12765 1606 12777 1658
rect 12829 1606 12841 1658
rect 12893 1606 12905 1658
rect 12957 1606 12969 1658
rect 13021 1606 20555 1658
rect 20607 1606 20619 1658
rect 20671 1606 20683 1658
rect 20735 1606 20747 1658
rect 20799 1606 20811 1658
rect 20863 1606 28397 1658
rect 28449 1606 28461 1658
rect 28513 1606 28525 1658
rect 28577 1606 28589 1658
rect 28641 1606 28653 1658
rect 28705 1606 32476 1658
rect 1104 1584 32476 1606
rect 1104 1114 32632 1136
rect 1104 1062 8792 1114
rect 8844 1062 8856 1114
rect 8908 1062 8920 1114
rect 8972 1062 8984 1114
rect 9036 1062 9048 1114
rect 9100 1062 16634 1114
rect 16686 1062 16698 1114
rect 16750 1062 16762 1114
rect 16814 1062 16826 1114
rect 16878 1062 16890 1114
rect 16942 1062 24476 1114
rect 24528 1062 24540 1114
rect 24592 1062 24604 1114
rect 24656 1062 24668 1114
rect 24720 1062 24732 1114
rect 24784 1062 32318 1114
rect 32370 1062 32382 1114
rect 32434 1062 32446 1114
rect 32498 1062 32510 1114
rect 32562 1062 32574 1114
rect 32626 1062 32632 1114
rect 1104 1040 32632 1062
<< via1 >>
rect 23664 21020 23716 21072
rect 26056 21020 26108 21072
rect 20076 20952 20128 21004
rect 25228 20952 25280 21004
rect 18512 20884 18564 20936
rect 24860 20884 24912 20936
rect 18880 20816 18932 20868
rect 30196 20816 30248 20868
rect 21088 20748 21140 20800
rect 30840 20748 30892 20800
rect 8792 20646 8844 20698
rect 8856 20646 8908 20698
rect 8920 20646 8972 20698
rect 8984 20646 9036 20698
rect 9048 20646 9100 20698
rect 16634 20646 16686 20698
rect 16698 20646 16750 20698
rect 16762 20646 16814 20698
rect 16826 20646 16878 20698
rect 16890 20646 16942 20698
rect 24476 20646 24528 20698
rect 24540 20646 24592 20698
rect 24604 20646 24656 20698
rect 24668 20646 24720 20698
rect 24732 20646 24784 20698
rect 32318 20646 32370 20698
rect 32382 20646 32434 20698
rect 32446 20646 32498 20698
rect 32510 20646 32562 20698
rect 32574 20646 32626 20698
rect 11980 20587 12032 20596
rect 11980 20553 11989 20587
rect 11989 20553 12023 20587
rect 12023 20553 12032 20587
rect 11980 20544 12032 20553
rect 12716 20587 12768 20596
rect 12716 20553 12725 20587
rect 12725 20553 12759 20587
rect 12759 20553 12768 20587
rect 12716 20544 12768 20553
rect 14832 20544 14884 20596
rect 15568 20544 15620 20596
rect 15844 20476 15896 20528
rect 14372 20408 14424 20460
rect 14648 20451 14700 20460
rect 14648 20417 14657 20451
rect 14657 20417 14691 20451
rect 14691 20417 14700 20451
rect 14648 20408 14700 20417
rect 15292 20408 15344 20460
rect 14464 20315 14516 20324
rect 14464 20281 14473 20315
rect 14473 20281 14507 20315
rect 14507 20281 14516 20315
rect 14464 20272 14516 20281
rect 16948 20408 17000 20460
rect 16396 20340 16448 20392
rect 17776 20587 17828 20596
rect 17776 20553 17785 20587
rect 17785 20553 17819 20587
rect 17819 20553 17828 20587
rect 17776 20544 17828 20553
rect 18696 20587 18748 20596
rect 18696 20553 18705 20587
rect 18705 20553 18739 20587
rect 18739 20553 18748 20587
rect 18696 20544 18748 20553
rect 18788 20408 18840 20460
rect 20076 20587 20128 20596
rect 20076 20553 20085 20587
rect 20085 20553 20119 20587
rect 20119 20553 20128 20587
rect 20076 20544 20128 20553
rect 20168 20544 20220 20596
rect 22192 20544 22244 20596
rect 19984 20476 20036 20528
rect 19800 20408 19852 20460
rect 21088 20451 21140 20460
rect 21088 20417 21097 20451
rect 21097 20417 21131 20451
rect 21131 20417 21140 20451
rect 21088 20408 21140 20417
rect 22928 20408 22980 20460
rect 19524 20340 19576 20392
rect 24584 20408 24636 20460
rect 24860 20544 24912 20596
rect 26056 20451 26108 20460
rect 26056 20417 26065 20451
rect 26065 20417 26099 20451
rect 26099 20417 26108 20451
rect 26056 20408 26108 20417
rect 19800 20272 19852 20324
rect 19892 20272 19944 20324
rect 21088 20272 21140 20324
rect 25596 20340 25648 20392
rect 28724 20476 28776 20528
rect 30196 20519 30248 20528
rect 30196 20485 30205 20519
rect 30205 20485 30239 20519
rect 30239 20485 30248 20519
rect 30196 20476 30248 20485
rect 30748 20476 30800 20528
rect 26516 20340 26568 20392
rect 29920 20383 29972 20392
rect 29920 20349 29929 20383
rect 29929 20349 29963 20383
rect 29963 20349 29972 20383
rect 29920 20340 29972 20349
rect 14648 20204 14700 20256
rect 16212 20204 16264 20256
rect 17040 20204 17092 20256
rect 20168 20204 20220 20256
rect 23388 20272 23440 20324
rect 24400 20204 24452 20256
rect 24492 20204 24544 20256
rect 24860 20204 24912 20256
rect 25320 20204 25372 20256
rect 4871 20102 4923 20154
rect 4935 20102 4987 20154
rect 4999 20102 5051 20154
rect 5063 20102 5115 20154
rect 5127 20102 5179 20154
rect 12713 20102 12765 20154
rect 12777 20102 12829 20154
rect 12841 20102 12893 20154
rect 12905 20102 12957 20154
rect 12969 20102 13021 20154
rect 20555 20102 20607 20154
rect 20619 20102 20671 20154
rect 20683 20102 20735 20154
rect 20747 20102 20799 20154
rect 20811 20102 20863 20154
rect 28397 20102 28449 20154
rect 28461 20102 28513 20154
rect 28525 20102 28577 20154
rect 28589 20102 28641 20154
rect 28653 20102 28705 20154
rect 2228 20043 2280 20052
rect 2228 20009 2237 20043
rect 2237 20009 2271 20043
rect 2271 20009 2280 20043
rect 2228 20000 2280 20009
rect 3056 20043 3108 20052
rect 3056 20009 3065 20043
rect 3065 20009 3099 20043
rect 3099 20009 3108 20043
rect 3056 20000 3108 20009
rect 4344 20043 4396 20052
rect 4344 20009 4353 20043
rect 4353 20009 4387 20043
rect 4387 20009 4396 20043
rect 4344 20000 4396 20009
rect 5264 20000 5316 20052
rect 5816 20043 5868 20052
rect 5816 20009 5825 20043
rect 5825 20009 5859 20043
rect 5859 20009 5868 20043
rect 5816 20000 5868 20009
rect 6552 20043 6604 20052
rect 6552 20009 6561 20043
rect 6561 20009 6595 20043
rect 6595 20009 6604 20043
rect 6552 20000 6604 20009
rect 9128 20000 9180 20052
rect 11060 20000 11112 20052
rect 13728 20000 13780 20052
rect 14372 20043 14424 20052
rect 14372 20009 14381 20043
rect 14381 20009 14415 20043
rect 14415 20009 14424 20043
rect 14372 20000 14424 20009
rect 15292 20043 15344 20052
rect 15292 20009 15301 20043
rect 15301 20009 15335 20043
rect 15335 20009 15344 20043
rect 15292 20000 15344 20009
rect 16028 20000 16080 20052
rect 14648 19932 14700 19984
rect 18880 20043 18932 20052
rect 18880 20009 18889 20043
rect 18889 20009 18923 20043
rect 18923 20009 18932 20043
rect 18880 20000 18932 20009
rect 4068 19796 4120 19848
rect 11060 19864 11112 19916
rect 14464 19864 14516 19916
rect 15476 19864 15528 19916
rect 16396 19864 16448 19916
rect 19616 19932 19668 19984
rect 16948 19864 17000 19916
rect 13176 19796 13228 19848
rect 13728 19839 13780 19848
rect 13728 19805 13737 19839
rect 13737 19805 13771 19839
rect 13771 19805 13780 19839
rect 13728 19796 13780 19805
rect 15568 19796 15620 19848
rect 16212 19728 16264 19780
rect 17868 19839 17920 19848
rect 17868 19805 17877 19839
rect 17877 19805 17911 19839
rect 17911 19805 17920 19839
rect 17868 19796 17920 19805
rect 18512 19839 18564 19848
rect 18512 19805 18521 19839
rect 18521 19805 18555 19839
rect 18555 19805 18564 19839
rect 18512 19796 18564 19805
rect 19708 19796 19760 19848
rect 24492 20000 24544 20052
rect 24584 20043 24636 20052
rect 24584 20009 24593 20043
rect 24593 20009 24627 20043
rect 24627 20009 24636 20043
rect 24584 20000 24636 20009
rect 23112 19932 23164 19984
rect 27436 20000 27488 20052
rect 19892 19864 19944 19916
rect 23388 19907 23440 19916
rect 23388 19873 23397 19907
rect 23397 19873 23431 19907
rect 23431 19873 23440 19907
rect 23388 19864 23440 19873
rect 21088 19796 21140 19848
rect 23296 19839 23348 19848
rect 23296 19805 23305 19839
rect 23305 19805 23339 19839
rect 23339 19805 23348 19839
rect 25964 19864 26016 19916
rect 26516 19864 26568 19916
rect 26792 19864 26844 19916
rect 23296 19796 23348 19805
rect 13360 19660 13412 19712
rect 15200 19660 15252 19712
rect 17316 19660 17368 19712
rect 22192 19771 22244 19780
rect 22192 19737 22201 19771
rect 22201 19737 22235 19771
rect 22235 19737 22244 19771
rect 22192 19728 22244 19737
rect 18236 19660 18288 19712
rect 19616 19660 19668 19712
rect 19800 19660 19852 19712
rect 20628 19703 20680 19712
rect 20628 19669 20637 19703
rect 20637 19669 20671 19703
rect 20671 19669 20680 19703
rect 20628 19660 20680 19669
rect 20996 19660 21048 19712
rect 21180 19660 21232 19712
rect 24124 19728 24176 19780
rect 24308 19660 24360 19712
rect 25044 19728 25096 19780
rect 31668 19864 31720 19916
rect 31760 19796 31812 19848
rect 25320 19660 25372 19712
rect 26240 19660 26292 19712
rect 26332 19660 26384 19712
rect 26792 19660 26844 19712
rect 27068 19660 27120 19712
rect 28724 19660 28776 19712
rect 30196 19703 30248 19712
rect 30196 19669 30205 19703
rect 30205 19669 30239 19703
rect 30239 19669 30248 19703
rect 30196 19660 30248 19669
rect 8792 19558 8844 19610
rect 8856 19558 8908 19610
rect 8920 19558 8972 19610
rect 8984 19558 9036 19610
rect 9048 19558 9100 19610
rect 16634 19558 16686 19610
rect 16698 19558 16750 19610
rect 16762 19558 16814 19610
rect 16826 19558 16878 19610
rect 16890 19558 16942 19610
rect 24476 19558 24528 19610
rect 24540 19558 24592 19610
rect 24604 19558 24656 19610
rect 24668 19558 24720 19610
rect 24732 19558 24784 19610
rect 32318 19558 32370 19610
rect 32382 19558 32434 19610
rect 32446 19558 32498 19610
rect 32510 19558 32562 19610
rect 32574 19558 32626 19610
rect 2412 19499 2464 19508
rect 2412 19465 2421 19499
rect 2421 19465 2455 19499
rect 2455 19465 2464 19499
rect 2412 19456 2464 19465
rect 3884 19499 3936 19508
rect 3884 19465 3893 19499
rect 3893 19465 3927 19499
rect 3927 19465 3936 19499
rect 3884 19456 3936 19465
rect 10968 19499 11020 19508
rect 10968 19465 10977 19499
rect 10977 19465 11011 19499
rect 11011 19465 11020 19499
rect 10968 19456 11020 19465
rect 11888 19456 11940 19508
rect 13176 19499 13228 19508
rect 13176 19465 13185 19499
rect 13185 19465 13219 19499
rect 13219 19465 13228 19499
rect 13176 19456 13228 19465
rect 4068 19363 4120 19372
rect 4068 19329 4077 19363
rect 4077 19329 4111 19363
rect 4111 19329 4120 19363
rect 4068 19320 4120 19329
rect 11152 19363 11204 19372
rect 11152 19329 11161 19363
rect 11161 19329 11195 19363
rect 11195 19329 11204 19363
rect 11152 19320 11204 19329
rect 13452 19388 13504 19440
rect 13728 19456 13780 19508
rect 16028 19456 16080 19508
rect 16120 19499 16172 19508
rect 16120 19465 16129 19499
rect 16129 19465 16163 19499
rect 16163 19465 16172 19499
rect 16120 19456 16172 19465
rect 17960 19456 18012 19508
rect 23112 19499 23164 19508
rect 23112 19465 23121 19499
rect 23121 19465 23155 19499
rect 23155 19465 23164 19499
rect 23112 19456 23164 19465
rect 23388 19456 23440 19508
rect 24952 19456 25004 19508
rect 27068 19456 27120 19508
rect 17040 19388 17092 19440
rect 17316 19431 17368 19440
rect 17316 19397 17325 19431
rect 17325 19397 17359 19431
rect 17359 19397 17368 19431
rect 17316 19388 17368 19397
rect 14464 19320 14516 19372
rect 17776 19320 17828 19372
rect 13544 19295 13596 19304
rect 13544 19261 13553 19295
rect 13553 19261 13587 19295
rect 13587 19261 13596 19295
rect 13544 19252 13596 19261
rect 15292 19295 15344 19304
rect 15292 19261 15301 19295
rect 15301 19261 15335 19295
rect 15335 19261 15344 19295
rect 15292 19252 15344 19261
rect 15476 19295 15528 19304
rect 15476 19261 15485 19295
rect 15485 19261 15519 19295
rect 15519 19261 15528 19295
rect 15476 19252 15528 19261
rect 13820 19184 13872 19236
rect 18236 19363 18288 19372
rect 18236 19329 18245 19363
rect 18245 19329 18279 19363
rect 18279 19329 18288 19363
rect 18236 19320 18288 19329
rect 18788 19320 18840 19372
rect 24860 19388 24912 19440
rect 26332 19388 26384 19440
rect 26424 19388 26476 19440
rect 27436 19431 27488 19440
rect 27436 19397 27445 19431
rect 27445 19397 27479 19431
rect 27479 19397 27488 19431
rect 27436 19388 27488 19397
rect 28724 19388 28776 19440
rect 30748 19456 30800 19508
rect 31484 19388 31536 19440
rect 31668 19388 31720 19440
rect 20628 19320 20680 19372
rect 21088 19320 21140 19372
rect 21456 19320 21508 19372
rect 19616 19252 19668 19304
rect 19892 19295 19944 19304
rect 19892 19261 19901 19295
rect 19901 19261 19935 19295
rect 19935 19261 19944 19295
rect 19892 19252 19944 19261
rect 21180 19252 21232 19304
rect 23296 19295 23348 19304
rect 23296 19261 23305 19295
rect 23305 19261 23339 19295
rect 23339 19261 23348 19295
rect 23296 19252 23348 19261
rect 23388 19295 23440 19304
rect 23388 19261 23397 19295
rect 23397 19261 23431 19295
rect 23431 19261 23440 19295
rect 23388 19252 23440 19261
rect 23664 19320 23716 19372
rect 24124 19363 24176 19372
rect 24124 19329 24133 19363
rect 24133 19329 24167 19363
rect 24167 19329 24176 19363
rect 24124 19320 24176 19329
rect 24308 19363 24360 19372
rect 24308 19329 24317 19363
rect 24317 19329 24351 19363
rect 24351 19329 24360 19363
rect 24308 19320 24360 19329
rect 26240 19252 26292 19304
rect 23664 19184 23716 19236
rect 23480 19116 23532 19168
rect 24308 19116 24360 19168
rect 26332 19116 26384 19168
rect 26516 19116 26568 19168
rect 30104 19252 30156 19304
rect 30012 19116 30064 19168
rect 4871 19014 4923 19066
rect 4935 19014 4987 19066
rect 4999 19014 5051 19066
rect 5063 19014 5115 19066
rect 5127 19014 5179 19066
rect 12713 19014 12765 19066
rect 12777 19014 12829 19066
rect 12841 19014 12893 19066
rect 12905 19014 12957 19066
rect 12969 19014 13021 19066
rect 20555 19014 20607 19066
rect 20619 19014 20671 19066
rect 20683 19014 20735 19066
rect 20747 19014 20799 19066
rect 20811 19014 20863 19066
rect 28397 19014 28449 19066
rect 28461 19014 28513 19066
rect 28525 19014 28577 19066
rect 28589 19014 28641 19066
rect 28653 19014 28705 19066
rect 11060 18912 11112 18964
rect 13360 18955 13412 18964
rect 13360 18921 13369 18955
rect 13369 18921 13403 18955
rect 13403 18921 13412 18955
rect 13360 18912 13412 18921
rect 11152 18844 11204 18896
rect 15844 18955 15896 18964
rect 15844 18921 15853 18955
rect 15853 18921 15887 18955
rect 15887 18921 15896 18955
rect 15844 18912 15896 18921
rect 16580 18912 16632 18964
rect 19708 18955 19760 18964
rect 19708 18921 19717 18955
rect 19717 18921 19751 18955
rect 19751 18921 19760 18955
rect 19708 18912 19760 18921
rect 20996 18912 21048 18964
rect 13544 18844 13596 18896
rect 15200 18844 15252 18896
rect 20260 18887 20312 18896
rect 20260 18853 20269 18887
rect 20269 18853 20303 18887
rect 20303 18853 20312 18887
rect 20260 18844 20312 18853
rect 21088 18844 21140 18896
rect 22008 18844 22060 18896
rect 11704 18751 11756 18760
rect 11704 18717 11713 18751
rect 11713 18717 11747 18751
rect 11747 18717 11756 18751
rect 11704 18708 11756 18717
rect 15292 18776 15344 18828
rect 13452 18640 13504 18692
rect 14464 18708 14516 18760
rect 15476 18708 15528 18760
rect 16396 18708 16448 18760
rect 17960 18708 18012 18760
rect 20904 18751 20956 18760
rect 20904 18717 20913 18751
rect 20913 18717 20947 18751
rect 20947 18717 20956 18751
rect 20904 18708 20956 18717
rect 22836 18776 22888 18828
rect 19708 18640 19760 18692
rect 19892 18615 19944 18624
rect 19892 18581 19901 18615
rect 19901 18581 19935 18615
rect 19935 18581 19944 18615
rect 19892 18572 19944 18581
rect 20260 18640 20312 18692
rect 23388 18776 23440 18828
rect 25044 18844 25096 18896
rect 25228 18887 25280 18896
rect 25228 18853 25237 18887
rect 25237 18853 25271 18887
rect 25271 18853 25280 18887
rect 25228 18844 25280 18853
rect 24124 18776 24176 18828
rect 23756 18708 23808 18760
rect 25136 18776 25188 18828
rect 24860 18708 24912 18760
rect 26332 18751 26384 18760
rect 26332 18717 26341 18751
rect 26341 18717 26375 18751
rect 26375 18717 26384 18751
rect 26332 18708 26384 18717
rect 27712 18708 27764 18760
rect 21088 18572 21140 18624
rect 23204 18572 23256 18624
rect 25136 18572 25188 18624
rect 25504 18640 25556 18692
rect 27620 18572 27672 18624
rect 28080 18615 28132 18624
rect 28080 18581 28089 18615
rect 28089 18581 28123 18615
rect 28123 18581 28132 18615
rect 28080 18572 28132 18581
rect 30104 18912 30156 18964
rect 30012 18751 30064 18760
rect 30012 18717 30021 18751
rect 30021 18717 30055 18751
rect 30055 18717 30064 18751
rect 30012 18708 30064 18717
rect 30748 18640 30800 18692
rect 8792 18470 8844 18522
rect 8856 18470 8908 18522
rect 8920 18470 8972 18522
rect 8984 18470 9036 18522
rect 9048 18470 9100 18522
rect 16634 18470 16686 18522
rect 16698 18470 16750 18522
rect 16762 18470 16814 18522
rect 16826 18470 16878 18522
rect 16890 18470 16942 18522
rect 24476 18470 24528 18522
rect 24540 18470 24592 18522
rect 24604 18470 24656 18522
rect 24668 18470 24720 18522
rect 24732 18470 24784 18522
rect 32318 18470 32370 18522
rect 32382 18470 32434 18522
rect 32446 18470 32498 18522
rect 32510 18470 32562 18522
rect 32574 18470 32626 18522
rect 11704 18368 11756 18420
rect 19800 18411 19852 18420
rect 19800 18377 19809 18411
rect 19809 18377 19843 18411
rect 19843 18377 19852 18411
rect 19800 18368 19852 18377
rect 19892 18368 19944 18420
rect 19524 18300 19576 18352
rect 19708 18300 19760 18352
rect 22836 18411 22888 18420
rect 22836 18377 22845 18411
rect 22845 18377 22879 18411
rect 22879 18377 22888 18411
rect 22836 18368 22888 18377
rect 23756 18411 23808 18420
rect 23756 18377 23765 18411
rect 23765 18377 23799 18411
rect 23799 18377 23808 18411
rect 23756 18368 23808 18377
rect 24952 18368 25004 18420
rect 25504 18368 25556 18420
rect 16396 18232 16448 18284
rect 22192 18300 22244 18352
rect 21180 18232 21232 18284
rect 23204 18343 23256 18352
rect 23204 18309 23213 18343
rect 23213 18309 23247 18343
rect 23247 18309 23256 18343
rect 23204 18300 23256 18309
rect 27712 18368 27764 18420
rect 28724 18368 28776 18420
rect 30012 18368 30064 18420
rect 23388 18232 23440 18284
rect 24400 18275 24452 18284
rect 24400 18241 24409 18275
rect 24409 18241 24443 18275
rect 24443 18241 24452 18275
rect 24400 18232 24452 18241
rect 19800 18096 19852 18148
rect 23480 18164 23532 18216
rect 30196 18232 30248 18284
rect 28080 18164 28132 18216
rect 19524 18028 19576 18080
rect 23664 18096 23716 18148
rect 24124 18096 24176 18148
rect 25596 18096 25648 18148
rect 22008 18028 22060 18080
rect 27620 18028 27672 18080
rect 4871 17926 4923 17978
rect 4935 17926 4987 17978
rect 4999 17926 5051 17978
rect 5063 17926 5115 17978
rect 5127 17926 5179 17978
rect 12713 17926 12765 17978
rect 12777 17926 12829 17978
rect 12841 17926 12893 17978
rect 12905 17926 12957 17978
rect 12969 17926 13021 17978
rect 20555 17926 20607 17978
rect 20619 17926 20671 17978
rect 20683 17926 20735 17978
rect 20747 17926 20799 17978
rect 20811 17926 20863 17978
rect 28397 17926 28449 17978
rect 28461 17926 28513 17978
rect 28525 17926 28577 17978
rect 28589 17926 28641 17978
rect 28653 17926 28705 17978
rect 26332 17867 26384 17876
rect 26332 17833 26341 17867
rect 26341 17833 26375 17867
rect 26375 17833 26384 17867
rect 26332 17824 26384 17833
rect 30840 17867 30892 17876
rect 30840 17833 30849 17867
rect 30849 17833 30883 17867
rect 30883 17833 30892 17867
rect 30840 17824 30892 17833
rect 31484 17867 31536 17876
rect 31484 17833 31493 17867
rect 31493 17833 31527 17867
rect 31527 17833 31536 17867
rect 31484 17824 31536 17833
rect 30196 17620 30248 17672
rect 30288 17620 30340 17672
rect 31300 17620 31352 17672
rect 8792 17382 8844 17434
rect 8856 17382 8908 17434
rect 8920 17382 8972 17434
rect 8984 17382 9036 17434
rect 9048 17382 9100 17434
rect 16634 17382 16686 17434
rect 16698 17382 16750 17434
rect 16762 17382 16814 17434
rect 16826 17382 16878 17434
rect 16890 17382 16942 17434
rect 24476 17382 24528 17434
rect 24540 17382 24592 17434
rect 24604 17382 24656 17434
rect 24668 17382 24720 17434
rect 24732 17382 24784 17434
rect 32318 17382 32370 17434
rect 32382 17382 32434 17434
rect 32446 17382 32498 17434
rect 32510 17382 32562 17434
rect 32574 17382 32626 17434
rect 4871 16838 4923 16890
rect 4935 16838 4987 16890
rect 4999 16838 5051 16890
rect 5063 16838 5115 16890
rect 5127 16838 5179 16890
rect 12713 16838 12765 16890
rect 12777 16838 12829 16890
rect 12841 16838 12893 16890
rect 12905 16838 12957 16890
rect 12969 16838 13021 16890
rect 20555 16838 20607 16890
rect 20619 16838 20671 16890
rect 20683 16838 20735 16890
rect 20747 16838 20799 16890
rect 20811 16838 20863 16890
rect 28397 16838 28449 16890
rect 28461 16838 28513 16890
rect 28525 16838 28577 16890
rect 28589 16838 28641 16890
rect 28653 16838 28705 16890
rect 8792 16294 8844 16346
rect 8856 16294 8908 16346
rect 8920 16294 8972 16346
rect 8984 16294 9036 16346
rect 9048 16294 9100 16346
rect 16634 16294 16686 16346
rect 16698 16294 16750 16346
rect 16762 16294 16814 16346
rect 16826 16294 16878 16346
rect 16890 16294 16942 16346
rect 24476 16294 24528 16346
rect 24540 16294 24592 16346
rect 24604 16294 24656 16346
rect 24668 16294 24720 16346
rect 24732 16294 24784 16346
rect 32318 16294 32370 16346
rect 32382 16294 32434 16346
rect 32446 16294 32498 16346
rect 32510 16294 32562 16346
rect 32574 16294 32626 16346
rect 4871 15750 4923 15802
rect 4935 15750 4987 15802
rect 4999 15750 5051 15802
rect 5063 15750 5115 15802
rect 5127 15750 5179 15802
rect 12713 15750 12765 15802
rect 12777 15750 12829 15802
rect 12841 15750 12893 15802
rect 12905 15750 12957 15802
rect 12969 15750 13021 15802
rect 20555 15750 20607 15802
rect 20619 15750 20671 15802
rect 20683 15750 20735 15802
rect 20747 15750 20799 15802
rect 20811 15750 20863 15802
rect 28397 15750 28449 15802
rect 28461 15750 28513 15802
rect 28525 15750 28577 15802
rect 28589 15750 28641 15802
rect 28653 15750 28705 15802
rect 8792 15206 8844 15258
rect 8856 15206 8908 15258
rect 8920 15206 8972 15258
rect 8984 15206 9036 15258
rect 9048 15206 9100 15258
rect 16634 15206 16686 15258
rect 16698 15206 16750 15258
rect 16762 15206 16814 15258
rect 16826 15206 16878 15258
rect 16890 15206 16942 15258
rect 24476 15206 24528 15258
rect 24540 15206 24592 15258
rect 24604 15206 24656 15258
rect 24668 15206 24720 15258
rect 24732 15206 24784 15258
rect 32318 15206 32370 15258
rect 32382 15206 32434 15258
rect 32446 15206 32498 15258
rect 32510 15206 32562 15258
rect 32574 15206 32626 15258
rect 4871 14662 4923 14714
rect 4935 14662 4987 14714
rect 4999 14662 5051 14714
rect 5063 14662 5115 14714
rect 5127 14662 5179 14714
rect 12713 14662 12765 14714
rect 12777 14662 12829 14714
rect 12841 14662 12893 14714
rect 12905 14662 12957 14714
rect 12969 14662 13021 14714
rect 20555 14662 20607 14714
rect 20619 14662 20671 14714
rect 20683 14662 20735 14714
rect 20747 14662 20799 14714
rect 20811 14662 20863 14714
rect 28397 14662 28449 14714
rect 28461 14662 28513 14714
rect 28525 14662 28577 14714
rect 28589 14662 28641 14714
rect 28653 14662 28705 14714
rect 8792 14118 8844 14170
rect 8856 14118 8908 14170
rect 8920 14118 8972 14170
rect 8984 14118 9036 14170
rect 9048 14118 9100 14170
rect 16634 14118 16686 14170
rect 16698 14118 16750 14170
rect 16762 14118 16814 14170
rect 16826 14118 16878 14170
rect 16890 14118 16942 14170
rect 24476 14118 24528 14170
rect 24540 14118 24592 14170
rect 24604 14118 24656 14170
rect 24668 14118 24720 14170
rect 24732 14118 24784 14170
rect 32318 14118 32370 14170
rect 32382 14118 32434 14170
rect 32446 14118 32498 14170
rect 32510 14118 32562 14170
rect 32574 14118 32626 14170
rect 4871 13574 4923 13626
rect 4935 13574 4987 13626
rect 4999 13574 5051 13626
rect 5063 13574 5115 13626
rect 5127 13574 5179 13626
rect 12713 13574 12765 13626
rect 12777 13574 12829 13626
rect 12841 13574 12893 13626
rect 12905 13574 12957 13626
rect 12969 13574 13021 13626
rect 20555 13574 20607 13626
rect 20619 13574 20671 13626
rect 20683 13574 20735 13626
rect 20747 13574 20799 13626
rect 20811 13574 20863 13626
rect 28397 13574 28449 13626
rect 28461 13574 28513 13626
rect 28525 13574 28577 13626
rect 28589 13574 28641 13626
rect 28653 13574 28705 13626
rect 8792 13030 8844 13082
rect 8856 13030 8908 13082
rect 8920 13030 8972 13082
rect 8984 13030 9036 13082
rect 9048 13030 9100 13082
rect 16634 13030 16686 13082
rect 16698 13030 16750 13082
rect 16762 13030 16814 13082
rect 16826 13030 16878 13082
rect 16890 13030 16942 13082
rect 24476 13030 24528 13082
rect 24540 13030 24592 13082
rect 24604 13030 24656 13082
rect 24668 13030 24720 13082
rect 24732 13030 24784 13082
rect 32318 13030 32370 13082
rect 32382 13030 32434 13082
rect 32446 13030 32498 13082
rect 32510 13030 32562 13082
rect 32574 13030 32626 13082
rect 4871 12486 4923 12538
rect 4935 12486 4987 12538
rect 4999 12486 5051 12538
rect 5063 12486 5115 12538
rect 5127 12486 5179 12538
rect 12713 12486 12765 12538
rect 12777 12486 12829 12538
rect 12841 12486 12893 12538
rect 12905 12486 12957 12538
rect 12969 12486 13021 12538
rect 20555 12486 20607 12538
rect 20619 12486 20671 12538
rect 20683 12486 20735 12538
rect 20747 12486 20799 12538
rect 20811 12486 20863 12538
rect 28397 12486 28449 12538
rect 28461 12486 28513 12538
rect 28525 12486 28577 12538
rect 28589 12486 28641 12538
rect 28653 12486 28705 12538
rect 8792 11942 8844 11994
rect 8856 11942 8908 11994
rect 8920 11942 8972 11994
rect 8984 11942 9036 11994
rect 9048 11942 9100 11994
rect 16634 11942 16686 11994
rect 16698 11942 16750 11994
rect 16762 11942 16814 11994
rect 16826 11942 16878 11994
rect 16890 11942 16942 11994
rect 24476 11942 24528 11994
rect 24540 11942 24592 11994
rect 24604 11942 24656 11994
rect 24668 11942 24720 11994
rect 24732 11942 24784 11994
rect 32318 11942 32370 11994
rect 32382 11942 32434 11994
rect 32446 11942 32498 11994
rect 32510 11942 32562 11994
rect 32574 11942 32626 11994
rect 4871 11398 4923 11450
rect 4935 11398 4987 11450
rect 4999 11398 5051 11450
rect 5063 11398 5115 11450
rect 5127 11398 5179 11450
rect 12713 11398 12765 11450
rect 12777 11398 12829 11450
rect 12841 11398 12893 11450
rect 12905 11398 12957 11450
rect 12969 11398 13021 11450
rect 20555 11398 20607 11450
rect 20619 11398 20671 11450
rect 20683 11398 20735 11450
rect 20747 11398 20799 11450
rect 20811 11398 20863 11450
rect 28397 11398 28449 11450
rect 28461 11398 28513 11450
rect 28525 11398 28577 11450
rect 28589 11398 28641 11450
rect 28653 11398 28705 11450
rect 8792 10854 8844 10906
rect 8856 10854 8908 10906
rect 8920 10854 8972 10906
rect 8984 10854 9036 10906
rect 9048 10854 9100 10906
rect 16634 10854 16686 10906
rect 16698 10854 16750 10906
rect 16762 10854 16814 10906
rect 16826 10854 16878 10906
rect 16890 10854 16942 10906
rect 24476 10854 24528 10906
rect 24540 10854 24592 10906
rect 24604 10854 24656 10906
rect 24668 10854 24720 10906
rect 24732 10854 24784 10906
rect 32318 10854 32370 10906
rect 32382 10854 32434 10906
rect 32446 10854 32498 10906
rect 32510 10854 32562 10906
rect 32574 10854 32626 10906
rect 4871 10310 4923 10362
rect 4935 10310 4987 10362
rect 4999 10310 5051 10362
rect 5063 10310 5115 10362
rect 5127 10310 5179 10362
rect 12713 10310 12765 10362
rect 12777 10310 12829 10362
rect 12841 10310 12893 10362
rect 12905 10310 12957 10362
rect 12969 10310 13021 10362
rect 20555 10310 20607 10362
rect 20619 10310 20671 10362
rect 20683 10310 20735 10362
rect 20747 10310 20799 10362
rect 20811 10310 20863 10362
rect 28397 10310 28449 10362
rect 28461 10310 28513 10362
rect 28525 10310 28577 10362
rect 28589 10310 28641 10362
rect 28653 10310 28705 10362
rect 8792 9766 8844 9818
rect 8856 9766 8908 9818
rect 8920 9766 8972 9818
rect 8984 9766 9036 9818
rect 9048 9766 9100 9818
rect 16634 9766 16686 9818
rect 16698 9766 16750 9818
rect 16762 9766 16814 9818
rect 16826 9766 16878 9818
rect 16890 9766 16942 9818
rect 24476 9766 24528 9818
rect 24540 9766 24592 9818
rect 24604 9766 24656 9818
rect 24668 9766 24720 9818
rect 24732 9766 24784 9818
rect 32318 9766 32370 9818
rect 32382 9766 32434 9818
rect 32446 9766 32498 9818
rect 32510 9766 32562 9818
rect 32574 9766 32626 9818
rect 4871 9222 4923 9274
rect 4935 9222 4987 9274
rect 4999 9222 5051 9274
rect 5063 9222 5115 9274
rect 5127 9222 5179 9274
rect 12713 9222 12765 9274
rect 12777 9222 12829 9274
rect 12841 9222 12893 9274
rect 12905 9222 12957 9274
rect 12969 9222 13021 9274
rect 20555 9222 20607 9274
rect 20619 9222 20671 9274
rect 20683 9222 20735 9274
rect 20747 9222 20799 9274
rect 20811 9222 20863 9274
rect 28397 9222 28449 9274
rect 28461 9222 28513 9274
rect 28525 9222 28577 9274
rect 28589 9222 28641 9274
rect 28653 9222 28705 9274
rect 8792 8678 8844 8730
rect 8856 8678 8908 8730
rect 8920 8678 8972 8730
rect 8984 8678 9036 8730
rect 9048 8678 9100 8730
rect 16634 8678 16686 8730
rect 16698 8678 16750 8730
rect 16762 8678 16814 8730
rect 16826 8678 16878 8730
rect 16890 8678 16942 8730
rect 24476 8678 24528 8730
rect 24540 8678 24592 8730
rect 24604 8678 24656 8730
rect 24668 8678 24720 8730
rect 24732 8678 24784 8730
rect 32318 8678 32370 8730
rect 32382 8678 32434 8730
rect 32446 8678 32498 8730
rect 32510 8678 32562 8730
rect 32574 8678 32626 8730
rect 4871 8134 4923 8186
rect 4935 8134 4987 8186
rect 4999 8134 5051 8186
rect 5063 8134 5115 8186
rect 5127 8134 5179 8186
rect 12713 8134 12765 8186
rect 12777 8134 12829 8186
rect 12841 8134 12893 8186
rect 12905 8134 12957 8186
rect 12969 8134 13021 8186
rect 20555 8134 20607 8186
rect 20619 8134 20671 8186
rect 20683 8134 20735 8186
rect 20747 8134 20799 8186
rect 20811 8134 20863 8186
rect 28397 8134 28449 8186
rect 28461 8134 28513 8186
rect 28525 8134 28577 8186
rect 28589 8134 28641 8186
rect 28653 8134 28705 8186
rect 8792 7590 8844 7642
rect 8856 7590 8908 7642
rect 8920 7590 8972 7642
rect 8984 7590 9036 7642
rect 9048 7590 9100 7642
rect 16634 7590 16686 7642
rect 16698 7590 16750 7642
rect 16762 7590 16814 7642
rect 16826 7590 16878 7642
rect 16890 7590 16942 7642
rect 24476 7590 24528 7642
rect 24540 7590 24592 7642
rect 24604 7590 24656 7642
rect 24668 7590 24720 7642
rect 24732 7590 24784 7642
rect 32318 7590 32370 7642
rect 32382 7590 32434 7642
rect 32446 7590 32498 7642
rect 32510 7590 32562 7642
rect 32574 7590 32626 7642
rect 4871 7046 4923 7098
rect 4935 7046 4987 7098
rect 4999 7046 5051 7098
rect 5063 7046 5115 7098
rect 5127 7046 5179 7098
rect 12713 7046 12765 7098
rect 12777 7046 12829 7098
rect 12841 7046 12893 7098
rect 12905 7046 12957 7098
rect 12969 7046 13021 7098
rect 20555 7046 20607 7098
rect 20619 7046 20671 7098
rect 20683 7046 20735 7098
rect 20747 7046 20799 7098
rect 20811 7046 20863 7098
rect 28397 7046 28449 7098
rect 28461 7046 28513 7098
rect 28525 7046 28577 7098
rect 28589 7046 28641 7098
rect 28653 7046 28705 7098
rect 8792 6502 8844 6554
rect 8856 6502 8908 6554
rect 8920 6502 8972 6554
rect 8984 6502 9036 6554
rect 9048 6502 9100 6554
rect 16634 6502 16686 6554
rect 16698 6502 16750 6554
rect 16762 6502 16814 6554
rect 16826 6502 16878 6554
rect 16890 6502 16942 6554
rect 24476 6502 24528 6554
rect 24540 6502 24592 6554
rect 24604 6502 24656 6554
rect 24668 6502 24720 6554
rect 24732 6502 24784 6554
rect 32318 6502 32370 6554
rect 32382 6502 32434 6554
rect 32446 6502 32498 6554
rect 32510 6502 32562 6554
rect 32574 6502 32626 6554
rect 4871 5958 4923 6010
rect 4935 5958 4987 6010
rect 4999 5958 5051 6010
rect 5063 5958 5115 6010
rect 5127 5958 5179 6010
rect 12713 5958 12765 6010
rect 12777 5958 12829 6010
rect 12841 5958 12893 6010
rect 12905 5958 12957 6010
rect 12969 5958 13021 6010
rect 20555 5958 20607 6010
rect 20619 5958 20671 6010
rect 20683 5958 20735 6010
rect 20747 5958 20799 6010
rect 20811 5958 20863 6010
rect 28397 5958 28449 6010
rect 28461 5958 28513 6010
rect 28525 5958 28577 6010
rect 28589 5958 28641 6010
rect 28653 5958 28705 6010
rect 8792 5414 8844 5466
rect 8856 5414 8908 5466
rect 8920 5414 8972 5466
rect 8984 5414 9036 5466
rect 9048 5414 9100 5466
rect 16634 5414 16686 5466
rect 16698 5414 16750 5466
rect 16762 5414 16814 5466
rect 16826 5414 16878 5466
rect 16890 5414 16942 5466
rect 24476 5414 24528 5466
rect 24540 5414 24592 5466
rect 24604 5414 24656 5466
rect 24668 5414 24720 5466
rect 24732 5414 24784 5466
rect 32318 5414 32370 5466
rect 32382 5414 32434 5466
rect 32446 5414 32498 5466
rect 32510 5414 32562 5466
rect 32574 5414 32626 5466
rect 4871 4870 4923 4922
rect 4935 4870 4987 4922
rect 4999 4870 5051 4922
rect 5063 4870 5115 4922
rect 5127 4870 5179 4922
rect 12713 4870 12765 4922
rect 12777 4870 12829 4922
rect 12841 4870 12893 4922
rect 12905 4870 12957 4922
rect 12969 4870 13021 4922
rect 20555 4870 20607 4922
rect 20619 4870 20671 4922
rect 20683 4870 20735 4922
rect 20747 4870 20799 4922
rect 20811 4870 20863 4922
rect 28397 4870 28449 4922
rect 28461 4870 28513 4922
rect 28525 4870 28577 4922
rect 28589 4870 28641 4922
rect 28653 4870 28705 4922
rect 8792 4326 8844 4378
rect 8856 4326 8908 4378
rect 8920 4326 8972 4378
rect 8984 4326 9036 4378
rect 9048 4326 9100 4378
rect 16634 4326 16686 4378
rect 16698 4326 16750 4378
rect 16762 4326 16814 4378
rect 16826 4326 16878 4378
rect 16890 4326 16942 4378
rect 24476 4326 24528 4378
rect 24540 4326 24592 4378
rect 24604 4326 24656 4378
rect 24668 4326 24720 4378
rect 24732 4326 24784 4378
rect 32318 4326 32370 4378
rect 32382 4326 32434 4378
rect 32446 4326 32498 4378
rect 32510 4326 32562 4378
rect 32574 4326 32626 4378
rect 4871 3782 4923 3834
rect 4935 3782 4987 3834
rect 4999 3782 5051 3834
rect 5063 3782 5115 3834
rect 5127 3782 5179 3834
rect 12713 3782 12765 3834
rect 12777 3782 12829 3834
rect 12841 3782 12893 3834
rect 12905 3782 12957 3834
rect 12969 3782 13021 3834
rect 20555 3782 20607 3834
rect 20619 3782 20671 3834
rect 20683 3782 20735 3834
rect 20747 3782 20799 3834
rect 20811 3782 20863 3834
rect 28397 3782 28449 3834
rect 28461 3782 28513 3834
rect 28525 3782 28577 3834
rect 28589 3782 28641 3834
rect 28653 3782 28705 3834
rect 8792 3238 8844 3290
rect 8856 3238 8908 3290
rect 8920 3238 8972 3290
rect 8984 3238 9036 3290
rect 9048 3238 9100 3290
rect 16634 3238 16686 3290
rect 16698 3238 16750 3290
rect 16762 3238 16814 3290
rect 16826 3238 16878 3290
rect 16890 3238 16942 3290
rect 24476 3238 24528 3290
rect 24540 3238 24592 3290
rect 24604 3238 24656 3290
rect 24668 3238 24720 3290
rect 24732 3238 24784 3290
rect 32318 3238 32370 3290
rect 32382 3238 32434 3290
rect 32446 3238 32498 3290
rect 32510 3238 32562 3290
rect 32574 3238 32626 3290
rect 4871 2694 4923 2746
rect 4935 2694 4987 2746
rect 4999 2694 5051 2746
rect 5063 2694 5115 2746
rect 5127 2694 5179 2746
rect 12713 2694 12765 2746
rect 12777 2694 12829 2746
rect 12841 2694 12893 2746
rect 12905 2694 12957 2746
rect 12969 2694 13021 2746
rect 20555 2694 20607 2746
rect 20619 2694 20671 2746
rect 20683 2694 20735 2746
rect 20747 2694 20799 2746
rect 20811 2694 20863 2746
rect 28397 2694 28449 2746
rect 28461 2694 28513 2746
rect 28525 2694 28577 2746
rect 28589 2694 28641 2746
rect 28653 2694 28705 2746
rect 8792 2150 8844 2202
rect 8856 2150 8908 2202
rect 8920 2150 8972 2202
rect 8984 2150 9036 2202
rect 9048 2150 9100 2202
rect 16634 2150 16686 2202
rect 16698 2150 16750 2202
rect 16762 2150 16814 2202
rect 16826 2150 16878 2202
rect 16890 2150 16942 2202
rect 24476 2150 24528 2202
rect 24540 2150 24592 2202
rect 24604 2150 24656 2202
rect 24668 2150 24720 2202
rect 24732 2150 24784 2202
rect 32318 2150 32370 2202
rect 32382 2150 32434 2202
rect 32446 2150 32498 2202
rect 32510 2150 32562 2202
rect 32574 2150 32626 2202
rect 4871 1606 4923 1658
rect 4935 1606 4987 1658
rect 4999 1606 5051 1658
rect 5063 1606 5115 1658
rect 5127 1606 5179 1658
rect 12713 1606 12765 1658
rect 12777 1606 12829 1658
rect 12841 1606 12893 1658
rect 12905 1606 12957 1658
rect 12969 1606 13021 1658
rect 20555 1606 20607 1658
rect 20619 1606 20671 1658
rect 20683 1606 20735 1658
rect 20747 1606 20799 1658
rect 20811 1606 20863 1658
rect 28397 1606 28449 1658
rect 28461 1606 28513 1658
rect 28525 1606 28577 1658
rect 28589 1606 28641 1658
rect 28653 1606 28705 1658
rect 8792 1062 8844 1114
rect 8856 1062 8908 1114
rect 8920 1062 8972 1114
rect 8984 1062 9036 1114
rect 9048 1062 9100 1114
rect 16634 1062 16686 1114
rect 16698 1062 16750 1114
rect 16762 1062 16814 1114
rect 16826 1062 16878 1114
rect 16890 1062 16942 1114
rect 24476 1062 24528 1114
rect 24540 1062 24592 1114
rect 24604 1062 24656 1114
rect 24668 1062 24720 1114
rect 24732 1062 24784 1114
rect 32318 1062 32370 1114
rect 32382 1062 32434 1114
rect 32446 1062 32498 1114
rect 32510 1062 32562 1114
rect 32574 1062 32626 1114
<< metal2 >>
rect 19982 21176 20038 21185
rect 19982 21111 20038 21120
rect 23662 21176 23718 21185
rect 23662 21111 23718 21120
rect 18512 20936 18564 20942
rect 5262 20904 5318 20913
rect 5262 20839 5318 20848
rect 9126 20904 9182 20913
rect 9126 20839 9182 20848
rect 17774 20904 17830 20913
rect 18512 20878 18564 20884
rect 17774 20839 17830 20848
rect 4871 20156 5179 20165
rect 4871 20154 4877 20156
rect 4933 20154 4957 20156
rect 5013 20154 5037 20156
rect 5093 20154 5117 20156
rect 5173 20154 5179 20156
rect 4933 20102 4935 20154
rect 5115 20102 5117 20154
rect 4871 20100 4877 20102
rect 4933 20100 4957 20102
rect 5013 20100 5037 20102
rect 5093 20100 5117 20102
rect 5173 20100 5179 20102
rect 2226 20088 2282 20097
rect 2226 20023 2228 20032
rect 2280 20023 2282 20032
rect 3054 20088 3110 20097
rect 3054 20023 3056 20032
rect 2228 19994 2280 20000
rect 3108 20023 3110 20032
rect 4342 20088 4398 20097
rect 4871 20091 5179 20100
rect 5276 20058 5304 20839
rect 8792 20700 9100 20709
rect 8792 20698 8798 20700
rect 8854 20698 8878 20700
rect 8934 20698 8958 20700
rect 9014 20698 9038 20700
rect 9094 20698 9100 20700
rect 8854 20646 8856 20698
rect 9036 20646 9038 20698
rect 8792 20644 8798 20646
rect 8854 20644 8878 20646
rect 8934 20644 8958 20646
rect 9014 20644 9038 20646
rect 9094 20644 9100 20646
rect 8792 20635 9100 20644
rect 5814 20088 5870 20097
rect 4342 20023 4344 20032
rect 3056 19994 3108 20000
rect 4396 20023 4398 20032
rect 5264 20052 5316 20058
rect 4344 19994 4396 20000
rect 5814 20023 5816 20032
rect 5264 19994 5316 20000
rect 5868 20023 5870 20032
rect 6550 20088 6606 20097
rect 9140 20058 9168 20839
rect 16634 20700 16942 20709
rect 16634 20698 16640 20700
rect 16696 20698 16720 20700
rect 16776 20698 16800 20700
rect 16856 20698 16880 20700
rect 16936 20698 16942 20700
rect 16696 20646 16698 20698
rect 16878 20646 16880 20698
rect 16634 20644 16640 20646
rect 16696 20644 16720 20646
rect 16776 20644 16800 20646
rect 16856 20644 16880 20646
rect 16936 20644 16942 20646
rect 11978 20632 12034 20641
rect 11978 20567 11980 20576
rect 12032 20567 12034 20576
rect 12714 20632 12770 20641
rect 12714 20567 12716 20576
rect 11980 20538 12032 20544
rect 12768 20567 12770 20576
rect 14830 20632 14886 20641
rect 16634 20635 16942 20644
rect 17788 20602 17816 20839
rect 17866 20768 17922 20777
rect 17866 20703 17922 20712
rect 14830 20567 14832 20576
rect 12716 20538 12768 20544
rect 14884 20567 14886 20576
rect 15568 20596 15620 20602
rect 14832 20538 14884 20544
rect 15568 20538 15620 20544
rect 17776 20596 17828 20602
rect 17776 20538 17828 20544
rect 11058 20496 11114 20505
rect 11058 20431 11114 20440
rect 14372 20460 14424 20466
rect 11072 20058 11100 20431
rect 14372 20402 14424 20408
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 15292 20460 15344 20466
rect 15292 20402 15344 20408
rect 12713 20156 13021 20165
rect 12713 20154 12719 20156
rect 12775 20154 12799 20156
rect 12855 20154 12879 20156
rect 12935 20154 12959 20156
rect 13015 20154 13021 20156
rect 12775 20102 12777 20154
rect 12957 20102 12959 20154
rect 12713 20100 12719 20102
rect 12775 20100 12799 20102
rect 12855 20100 12879 20102
rect 12935 20100 12959 20102
rect 13015 20100 13021 20102
rect 12713 20091 13021 20100
rect 13726 20088 13782 20097
rect 6550 20023 6552 20032
rect 5816 19994 5868 20000
rect 6604 20023 6606 20032
rect 9128 20052 9180 20058
rect 6552 19994 6604 20000
rect 9128 19994 9180 20000
rect 11060 20052 11112 20058
rect 14384 20058 14412 20402
rect 14464 20324 14516 20330
rect 14464 20266 14516 20272
rect 13726 20023 13728 20032
rect 11060 19994 11112 20000
rect 13780 20023 13782 20032
rect 14372 20052 14424 20058
rect 13728 19994 13780 20000
rect 14372 19994 14424 20000
rect 11058 19952 11114 19961
rect 14476 19922 14504 20266
rect 14660 20262 14688 20402
rect 14648 20256 14700 20262
rect 14648 20198 14700 20204
rect 14660 19990 14688 20198
rect 15304 20058 15332 20402
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 14648 19984 14700 19990
rect 14648 19926 14700 19932
rect 11058 19887 11060 19896
rect 11112 19887 11114 19896
rect 14464 19916 14516 19922
rect 11060 19858 11112 19864
rect 14464 19858 14516 19864
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 4068 19848 4120 19854
rect 4068 19790 4120 19796
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 2410 19544 2466 19553
rect 2410 19479 2412 19488
rect 2464 19479 2466 19488
rect 3882 19544 3938 19553
rect 3882 19479 3884 19488
rect 2412 19450 2464 19456
rect 3936 19479 3938 19488
rect 3884 19450 3936 19456
rect 4080 19378 4108 19790
rect 8792 19612 9100 19621
rect 8792 19610 8798 19612
rect 8854 19610 8878 19612
rect 8934 19610 8958 19612
rect 9014 19610 9038 19612
rect 9094 19610 9100 19612
rect 8854 19558 8856 19610
rect 9036 19558 9038 19610
rect 8792 19556 8798 19558
rect 8854 19556 8878 19558
rect 8934 19556 8958 19558
rect 9014 19556 9038 19558
rect 9094 19556 9100 19558
rect 8792 19547 9100 19556
rect 10966 19544 11022 19553
rect 10966 19479 10968 19488
rect 11020 19479 11022 19488
rect 11886 19544 11942 19553
rect 13188 19514 13216 19790
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 11886 19479 11888 19488
rect 10968 19450 11020 19456
rect 11940 19479 11942 19488
rect 13176 19508 13228 19514
rect 11888 19450 11940 19456
rect 13176 19450 13228 19456
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 11152 19372 11204 19378
rect 11152 19314 11204 19320
rect 4871 19068 5179 19077
rect 4871 19066 4877 19068
rect 4933 19066 4957 19068
rect 5013 19066 5037 19068
rect 5093 19066 5117 19068
rect 5173 19066 5179 19068
rect 4933 19014 4935 19066
rect 5115 19014 5117 19066
rect 4871 19012 4877 19014
rect 4933 19012 4957 19014
rect 5013 19012 5037 19014
rect 5093 19012 5117 19014
rect 5173 19012 5179 19014
rect 4871 19003 5179 19012
rect 11058 19000 11114 19009
rect 11058 18935 11060 18944
rect 11112 18935 11114 18944
rect 11060 18906 11112 18912
rect 11164 18902 11192 19314
rect 12713 19068 13021 19077
rect 12713 19066 12719 19068
rect 12775 19066 12799 19068
rect 12855 19066 12879 19068
rect 12935 19066 12959 19068
rect 13015 19066 13021 19068
rect 12775 19014 12777 19066
rect 12957 19014 12959 19066
rect 12713 19012 12719 19014
rect 12775 19012 12799 19014
rect 12855 19012 12879 19014
rect 12935 19012 12959 19014
rect 13015 19012 13021 19014
rect 12713 19003 13021 19012
rect 13372 18970 13400 19654
rect 13740 19514 13768 19790
rect 13728 19508 13780 19514
rect 13728 19450 13780 19456
rect 13452 19440 13504 19446
rect 13452 19382 13504 19388
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 11152 18896 11204 18902
rect 11152 18838 11204 18844
rect 11704 18760 11756 18766
rect 11704 18702 11756 18708
rect 8792 18524 9100 18533
rect 8792 18522 8798 18524
rect 8854 18522 8878 18524
rect 8934 18522 8958 18524
rect 9014 18522 9038 18524
rect 9094 18522 9100 18524
rect 8854 18470 8856 18522
rect 9036 18470 9038 18522
rect 8792 18468 8798 18470
rect 8854 18468 8878 18470
rect 8934 18468 8958 18470
rect 9014 18468 9038 18470
rect 9094 18468 9100 18470
rect 8792 18459 9100 18468
rect 11716 18426 11744 18702
rect 13464 18698 13492 19382
rect 14476 19378 14504 19858
rect 15200 19712 15252 19718
rect 15200 19654 15252 19660
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 13818 19272 13874 19281
rect 13556 18902 13584 19246
rect 13818 19207 13820 19216
rect 13872 19207 13874 19216
rect 13820 19178 13872 19184
rect 13544 18896 13596 18902
rect 13544 18838 13596 18844
rect 14476 18766 14504 19314
rect 15212 18902 15240 19654
rect 15488 19310 15516 19858
rect 15580 19854 15608 20538
rect 15844 20528 15896 20534
rect 15844 20470 15896 20476
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 15200 18896 15252 18902
rect 15200 18838 15252 18844
rect 15304 18834 15332 19246
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 15488 18766 15516 19246
rect 15856 18970 15884 20470
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 16396 20392 16448 20398
rect 16396 20334 16448 20340
rect 16212 20256 16264 20262
rect 16212 20198 16264 20204
rect 16028 20052 16080 20058
rect 16028 19994 16080 20000
rect 16040 19514 16068 19994
rect 16224 19786 16252 20198
rect 16408 19922 16436 20334
rect 16960 19922 16988 20402
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 16212 19780 16264 19786
rect 16212 19722 16264 19728
rect 16118 19544 16174 19553
rect 16028 19508 16080 19514
rect 16118 19479 16120 19488
rect 16028 19450 16080 19456
rect 16172 19479 16174 19488
rect 16120 19450 16172 19456
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 16408 18766 16436 19858
rect 16634 19612 16942 19621
rect 16634 19610 16640 19612
rect 16696 19610 16720 19612
rect 16776 19610 16800 19612
rect 16856 19610 16880 19612
rect 16936 19610 16942 19612
rect 16696 19558 16698 19610
rect 16878 19558 16880 19610
rect 16634 19556 16640 19558
rect 16696 19556 16720 19558
rect 16776 19556 16800 19558
rect 16856 19556 16880 19558
rect 16936 19556 16942 19558
rect 16634 19547 16942 19556
rect 17052 19446 17080 20198
rect 17880 19854 17908 20703
rect 18524 19854 18552 20878
rect 18880 20868 18932 20874
rect 18880 20810 18932 20816
rect 18694 20632 18750 20641
rect 18694 20567 18696 20576
rect 18748 20567 18750 20576
rect 18696 20538 18748 20544
rect 18788 20460 18840 20466
rect 18788 20402 18840 20408
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 18512 19848 18564 19854
rect 18512 19790 18564 19796
rect 17316 19712 17368 19718
rect 17316 19654 17368 19660
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 17328 19446 17356 19654
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 17040 19440 17092 19446
rect 17040 19382 17092 19388
rect 17316 19440 17368 19446
rect 17316 19382 17368 19388
rect 17774 19408 17830 19417
rect 17774 19343 17776 19352
rect 17828 19343 17830 19352
rect 17776 19314 17828 19320
rect 16578 19000 16634 19009
rect 16578 18935 16580 18944
rect 16632 18935 16634 18944
rect 16580 18906 16632 18912
rect 17972 18766 18000 19450
rect 18248 19378 18276 19654
rect 18800 19378 18828 20402
rect 18892 20058 18920 20810
rect 19996 20534 20024 21111
rect 23676 21078 23704 21111
rect 23664 21072 23716 21078
rect 22190 21040 22246 21049
rect 20076 21004 20128 21010
rect 22190 20975 22246 20984
rect 22926 21040 22982 21049
rect 23664 21014 23716 21020
rect 26056 21072 26108 21078
rect 26056 21014 26108 21020
rect 22926 20975 22982 20984
rect 25228 21004 25280 21010
rect 20076 20946 20128 20952
rect 20088 20602 20116 20946
rect 20902 20904 20958 20913
rect 20902 20839 20958 20848
rect 20076 20596 20128 20602
rect 20076 20538 20128 20544
rect 20168 20596 20220 20602
rect 20168 20538 20220 20544
rect 19984 20528 20036 20534
rect 19984 20470 20036 20476
rect 19800 20460 19852 20466
rect 19800 20402 19852 20408
rect 19524 20392 19576 20398
rect 19524 20334 19576 20340
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 18236 19372 18288 19378
rect 18236 19314 18288 19320
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 13452 18692 13504 18698
rect 13452 18634 13504 18640
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 16408 18290 16436 18702
rect 16634 18524 16942 18533
rect 16634 18522 16640 18524
rect 16696 18522 16720 18524
rect 16776 18522 16800 18524
rect 16856 18522 16880 18524
rect 16936 18522 16942 18524
rect 16696 18470 16698 18522
rect 16878 18470 16880 18522
rect 16634 18468 16640 18470
rect 16696 18468 16720 18470
rect 16776 18468 16800 18470
rect 16856 18468 16880 18470
rect 16936 18468 16942 18470
rect 16634 18459 16942 18468
rect 19536 18358 19564 20334
rect 19812 20330 19840 20402
rect 19800 20324 19852 20330
rect 19800 20266 19852 20272
rect 19892 20324 19944 20330
rect 19892 20266 19944 20272
rect 19616 19984 19668 19990
rect 19616 19926 19668 19932
rect 19628 19718 19656 19926
rect 19904 19922 19932 20266
rect 20180 20262 20208 20538
rect 20168 20256 20220 20262
rect 20168 20198 20220 20204
rect 20555 20156 20863 20165
rect 20555 20154 20561 20156
rect 20617 20154 20641 20156
rect 20697 20154 20721 20156
rect 20777 20154 20801 20156
rect 20857 20154 20863 20156
rect 20617 20102 20619 20154
rect 20799 20102 20801 20154
rect 20555 20100 20561 20102
rect 20617 20100 20641 20102
rect 20697 20100 20721 20102
rect 20777 20100 20801 20102
rect 20857 20100 20863 20102
rect 20555 20091 20863 20100
rect 19892 19916 19944 19922
rect 19892 19858 19944 19864
rect 19708 19848 19760 19854
rect 19708 19790 19760 19796
rect 19616 19712 19668 19718
rect 19616 19654 19668 19660
rect 19616 19304 19668 19310
rect 19616 19246 19668 19252
rect 19628 18850 19656 19246
rect 19720 18970 19748 19790
rect 19800 19712 19852 19718
rect 19800 19654 19852 19660
rect 19708 18964 19760 18970
rect 19708 18906 19760 18912
rect 19628 18822 19748 18850
rect 19720 18698 19748 18822
rect 19708 18692 19760 18698
rect 19708 18634 19760 18640
rect 19720 18358 19748 18634
rect 19812 18426 19840 19654
rect 19904 19310 19932 19858
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20640 19378 20668 19654
rect 20628 19372 20680 19378
rect 20628 19314 20680 19320
rect 19892 19304 19944 19310
rect 19892 19246 19944 19252
rect 20555 19068 20863 19077
rect 20555 19066 20561 19068
rect 20617 19066 20641 19068
rect 20697 19066 20721 19068
rect 20777 19066 20801 19068
rect 20857 19066 20863 19068
rect 20617 19014 20619 19066
rect 20799 19014 20801 19066
rect 20555 19012 20561 19014
rect 20617 19012 20641 19014
rect 20697 19012 20721 19014
rect 20777 19012 20801 19014
rect 20857 19012 20863 19014
rect 20555 19003 20863 19012
rect 20260 18896 20312 18902
rect 20260 18838 20312 18844
rect 20272 18698 20300 18838
rect 20916 18766 20944 20839
rect 21088 20800 21140 20806
rect 21088 20742 21140 20748
rect 21100 20466 21128 20742
rect 22204 20602 22232 20975
rect 22192 20596 22244 20602
rect 22192 20538 22244 20544
rect 21454 20496 21510 20505
rect 21088 20460 21140 20466
rect 22940 20466 22968 20975
rect 25228 20946 25280 20952
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 24476 20700 24784 20709
rect 24476 20698 24482 20700
rect 24538 20698 24562 20700
rect 24618 20698 24642 20700
rect 24698 20698 24722 20700
rect 24778 20698 24784 20700
rect 24538 20646 24540 20698
rect 24720 20646 24722 20698
rect 24476 20644 24482 20646
rect 24538 20644 24562 20646
rect 24618 20644 24642 20646
rect 24698 20644 24722 20646
rect 24778 20644 24784 20646
rect 24476 20635 24784 20644
rect 24872 20602 24900 20878
rect 24860 20596 24912 20602
rect 24860 20538 24912 20544
rect 21454 20431 21510 20440
rect 22928 20460 22980 20466
rect 21088 20402 21140 20408
rect 21088 20324 21140 20330
rect 21088 20266 21140 20272
rect 21100 19854 21128 20266
rect 21088 19848 21140 19854
rect 21088 19790 21140 19796
rect 20996 19712 21048 19718
rect 20996 19654 21048 19660
rect 21180 19712 21232 19718
rect 21180 19654 21232 19660
rect 21008 18970 21036 19654
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 21100 18902 21128 19314
rect 21192 19310 21220 19654
rect 21468 19378 21496 20431
rect 22928 20402 22980 20408
rect 24584 20460 24636 20466
rect 24584 20402 24636 20408
rect 23388 20324 23440 20330
rect 23388 20266 23440 20272
rect 23112 19984 23164 19990
rect 23112 19926 23164 19932
rect 22192 19780 22244 19786
rect 22192 19722 22244 19728
rect 21456 19372 21508 19378
rect 21456 19314 21508 19320
rect 21180 19304 21232 19310
rect 21180 19246 21232 19252
rect 21088 18896 21140 18902
rect 21088 18838 21140 18844
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20260 18692 20312 18698
rect 20260 18634 20312 18640
rect 21100 18630 21128 18838
rect 19892 18624 19944 18630
rect 19892 18566 19944 18572
rect 21088 18624 21140 18630
rect 21088 18566 21140 18572
rect 19904 18426 19932 18566
rect 19800 18420 19852 18426
rect 19800 18362 19852 18368
rect 19892 18420 19944 18426
rect 19892 18362 19944 18368
rect 19524 18352 19576 18358
rect 19524 18294 19576 18300
rect 19708 18352 19760 18358
rect 19708 18294 19760 18300
rect 16396 18284 16448 18290
rect 16396 18226 16448 18232
rect 19536 18086 19564 18294
rect 19812 18154 19840 18362
rect 21192 18290 21220 19246
rect 22008 18896 22060 18902
rect 22008 18838 22060 18844
rect 21180 18284 21232 18290
rect 21180 18226 21232 18232
rect 19800 18148 19852 18154
rect 19800 18090 19852 18096
rect 22020 18086 22048 18838
rect 22204 18358 22232 19722
rect 23124 19514 23152 19926
rect 23400 19922 23428 20266
rect 24400 20256 24452 20262
rect 24400 20198 24452 20204
rect 24492 20256 24544 20262
rect 24492 20198 24544 20204
rect 23388 19916 23440 19922
rect 23388 19858 23440 19864
rect 23296 19848 23348 19854
rect 23296 19790 23348 19796
rect 23112 19508 23164 19514
rect 23112 19450 23164 19456
rect 23308 19310 23336 19790
rect 23400 19514 23428 19858
rect 24124 19780 24176 19786
rect 24124 19722 24176 19728
rect 23388 19508 23440 19514
rect 23388 19450 23440 19456
rect 24136 19378 24164 19722
rect 24308 19712 24360 19718
rect 24308 19654 24360 19660
rect 24320 19378 24348 19654
rect 23664 19372 23716 19378
rect 23664 19314 23716 19320
rect 24124 19372 24176 19378
rect 24124 19314 24176 19320
rect 24308 19372 24360 19378
rect 24308 19314 24360 19320
rect 23296 19304 23348 19310
rect 23296 19246 23348 19252
rect 23388 19304 23440 19310
rect 23440 19264 23520 19292
rect 23388 19246 23440 19252
rect 23492 19174 23520 19264
rect 23676 19242 23704 19314
rect 23664 19236 23716 19242
rect 23664 19178 23716 19184
rect 23480 19168 23532 19174
rect 23480 19110 23532 19116
rect 22836 18828 22888 18834
rect 22836 18770 22888 18776
rect 23388 18828 23440 18834
rect 23388 18770 23440 18776
rect 22848 18426 22876 18770
rect 23204 18624 23256 18630
rect 23204 18566 23256 18572
rect 22836 18420 22888 18426
rect 22836 18362 22888 18368
rect 23216 18358 23244 18566
rect 22192 18352 22244 18358
rect 22192 18294 22244 18300
rect 23204 18352 23256 18358
rect 23204 18294 23256 18300
rect 23400 18290 23428 18770
rect 23388 18284 23440 18290
rect 23388 18226 23440 18232
rect 23492 18222 23520 19110
rect 23480 18216 23532 18222
rect 23480 18158 23532 18164
rect 23676 18154 23704 19178
rect 24320 19174 24348 19314
rect 24308 19168 24360 19174
rect 24308 19110 24360 19116
rect 24124 18828 24176 18834
rect 24124 18770 24176 18776
rect 23756 18760 23808 18766
rect 23756 18702 23808 18708
rect 23768 18426 23796 18702
rect 23756 18420 23808 18426
rect 23756 18362 23808 18368
rect 24136 18154 24164 18770
rect 24412 18290 24440 20198
rect 24504 20058 24532 20198
rect 24596 20058 24624 20402
rect 24860 20256 24912 20262
rect 24860 20198 24912 20204
rect 24492 20052 24544 20058
rect 24492 19994 24544 20000
rect 24584 20052 24636 20058
rect 24584 19994 24636 20000
rect 24476 19612 24784 19621
rect 24476 19610 24482 19612
rect 24538 19610 24562 19612
rect 24618 19610 24642 19612
rect 24698 19610 24722 19612
rect 24778 19610 24784 19612
rect 24538 19558 24540 19610
rect 24720 19558 24722 19610
rect 24476 19556 24482 19558
rect 24538 19556 24562 19558
rect 24618 19556 24642 19558
rect 24698 19556 24722 19558
rect 24778 19556 24784 19558
rect 24476 19547 24784 19556
rect 24872 19446 24900 20198
rect 25044 19780 25096 19786
rect 25044 19722 25096 19728
rect 24952 19508 25004 19514
rect 24952 19450 25004 19456
rect 24860 19440 24912 19446
rect 24860 19382 24912 19388
rect 24858 19272 24914 19281
rect 24858 19207 24914 19216
rect 24872 18766 24900 19207
rect 24860 18760 24912 18766
rect 24860 18702 24912 18708
rect 24476 18524 24784 18533
rect 24476 18522 24482 18524
rect 24538 18522 24562 18524
rect 24618 18522 24642 18524
rect 24698 18522 24722 18524
rect 24778 18522 24784 18524
rect 24538 18470 24540 18522
rect 24720 18470 24722 18522
rect 24476 18468 24482 18470
rect 24538 18468 24562 18470
rect 24618 18468 24642 18470
rect 24698 18468 24722 18470
rect 24778 18468 24784 18470
rect 24476 18459 24784 18468
rect 24964 18426 24992 19450
rect 25056 18902 25084 19722
rect 25240 18902 25268 20946
rect 26068 20466 26096 21014
rect 30196 20868 30248 20874
rect 30196 20810 30248 20816
rect 30208 20534 30236 20810
rect 30840 20800 30892 20806
rect 30840 20742 30892 20748
rect 31758 20768 31814 20777
rect 28724 20528 28776 20534
rect 28724 20470 28776 20476
rect 30196 20528 30248 20534
rect 30196 20470 30248 20476
rect 30748 20528 30800 20534
rect 30748 20470 30800 20476
rect 26056 20460 26108 20466
rect 26056 20402 26108 20408
rect 25596 20392 25648 20398
rect 25596 20334 25648 20340
rect 26516 20392 26568 20398
rect 26516 20334 26568 20340
rect 25320 20256 25372 20262
rect 25320 20198 25372 20204
rect 25332 19718 25360 20198
rect 25320 19712 25372 19718
rect 25320 19654 25372 19660
rect 25044 18896 25096 18902
rect 25044 18838 25096 18844
rect 25228 18896 25280 18902
rect 25228 18838 25280 18844
rect 25136 18828 25188 18834
rect 25136 18770 25188 18776
rect 25148 18630 25176 18770
rect 25504 18692 25556 18698
rect 25504 18634 25556 18640
rect 25136 18624 25188 18630
rect 25136 18566 25188 18572
rect 25516 18426 25544 18634
rect 24952 18420 25004 18426
rect 24952 18362 25004 18368
rect 25504 18420 25556 18426
rect 25504 18362 25556 18368
rect 24400 18284 24452 18290
rect 24400 18226 24452 18232
rect 25608 18154 25636 20334
rect 26528 19922 26556 20334
rect 28397 20156 28705 20165
rect 28397 20154 28403 20156
rect 28459 20154 28483 20156
rect 28539 20154 28563 20156
rect 28619 20154 28643 20156
rect 28699 20154 28705 20156
rect 28459 20102 28461 20154
rect 28641 20102 28643 20154
rect 28397 20100 28403 20102
rect 28459 20100 28483 20102
rect 28539 20100 28563 20102
rect 28619 20100 28643 20102
rect 28699 20100 28705 20102
rect 28397 20091 28705 20100
rect 27436 20052 27488 20058
rect 27436 19994 27488 20000
rect 25964 19916 26016 19922
rect 25964 19858 26016 19864
rect 26516 19916 26568 19922
rect 26516 19858 26568 19864
rect 26792 19916 26844 19922
rect 26792 19858 26844 19864
rect 25976 19802 26004 19858
rect 25976 19774 26464 19802
rect 26240 19712 26292 19718
rect 26240 19654 26292 19660
rect 26332 19712 26384 19718
rect 26332 19654 26384 19660
rect 26252 19310 26280 19654
rect 26344 19446 26372 19654
rect 26436 19446 26464 19774
rect 26332 19440 26384 19446
rect 26332 19382 26384 19388
rect 26424 19440 26476 19446
rect 26424 19382 26476 19388
rect 26240 19304 26292 19310
rect 26240 19246 26292 19252
rect 26528 19174 26556 19858
rect 26804 19718 26832 19858
rect 26792 19712 26844 19718
rect 26792 19654 26844 19660
rect 27068 19712 27120 19718
rect 27068 19654 27120 19660
rect 27080 19514 27108 19654
rect 27068 19508 27120 19514
rect 27068 19450 27120 19456
rect 27448 19446 27476 19994
rect 28736 19718 28764 20470
rect 29920 20392 29972 20398
rect 29920 20334 29972 20340
rect 28724 19712 28776 19718
rect 28724 19654 28776 19660
rect 28736 19446 28764 19654
rect 27436 19440 27488 19446
rect 27436 19382 27488 19388
rect 28724 19440 28776 19446
rect 28724 19382 28776 19388
rect 26332 19168 26384 19174
rect 26332 19110 26384 19116
rect 26516 19168 26568 19174
rect 26516 19110 26568 19116
rect 26344 18766 26372 19110
rect 28397 19068 28705 19077
rect 28397 19066 28403 19068
rect 28459 19066 28483 19068
rect 28539 19066 28563 19068
rect 28619 19066 28643 19068
rect 28699 19066 28705 19068
rect 28459 19014 28461 19066
rect 28641 19014 28643 19066
rect 28397 19012 28403 19014
rect 28459 19012 28483 19014
rect 28539 19012 28563 19014
rect 28619 19012 28643 19014
rect 28699 19012 28705 19014
rect 28397 19003 28705 19012
rect 26332 18760 26384 18766
rect 26332 18702 26384 18708
rect 27712 18760 27764 18766
rect 27712 18702 27764 18708
rect 23664 18148 23716 18154
rect 23664 18090 23716 18096
rect 24124 18148 24176 18154
rect 24124 18090 24176 18096
rect 25596 18148 25648 18154
rect 25596 18090 25648 18096
rect 19524 18080 19576 18086
rect 19524 18022 19576 18028
rect 22008 18080 22060 18086
rect 22008 18022 22060 18028
rect 4871 17980 5179 17989
rect 4871 17978 4877 17980
rect 4933 17978 4957 17980
rect 5013 17978 5037 17980
rect 5093 17978 5117 17980
rect 5173 17978 5179 17980
rect 4933 17926 4935 17978
rect 5115 17926 5117 17978
rect 4871 17924 4877 17926
rect 4933 17924 4957 17926
rect 5013 17924 5037 17926
rect 5093 17924 5117 17926
rect 5173 17924 5179 17926
rect 4871 17915 5179 17924
rect 12713 17980 13021 17989
rect 12713 17978 12719 17980
rect 12775 17978 12799 17980
rect 12855 17978 12879 17980
rect 12935 17978 12959 17980
rect 13015 17978 13021 17980
rect 12775 17926 12777 17978
rect 12957 17926 12959 17978
rect 12713 17924 12719 17926
rect 12775 17924 12799 17926
rect 12855 17924 12879 17926
rect 12935 17924 12959 17926
rect 13015 17924 13021 17926
rect 12713 17915 13021 17924
rect 20555 17980 20863 17989
rect 20555 17978 20561 17980
rect 20617 17978 20641 17980
rect 20697 17978 20721 17980
rect 20777 17978 20801 17980
rect 20857 17978 20863 17980
rect 20617 17926 20619 17978
rect 20799 17926 20801 17978
rect 20555 17924 20561 17926
rect 20617 17924 20641 17926
rect 20697 17924 20721 17926
rect 20777 17924 20801 17926
rect 20857 17924 20863 17926
rect 20555 17915 20863 17924
rect 26344 17882 26372 18702
rect 27620 18624 27672 18630
rect 27620 18566 27672 18572
rect 27632 18086 27660 18566
rect 27724 18426 27752 18702
rect 28080 18624 28132 18630
rect 28080 18566 28132 18572
rect 27712 18420 27764 18426
rect 27712 18362 27764 18368
rect 28092 18222 28120 18566
rect 28736 18426 28764 19382
rect 29932 19258 29960 20334
rect 30196 19712 30248 19718
rect 30196 19654 30248 19660
rect 30104 19304 30156 19310
rect 29932 19230 30052 19258
rect 30104 19246 30156 19252
rect 30024 19174 30052 19230
rect 30012 19168 30064 19174
rect 30012 19110 30064 19116
rect 30024 18766 30052 19110
rect 30116 18970 30144 19246
rect 30104 18964 30156 18970
rect 30104 18906 30156 18912
rect 30012 18760 30064 18766
rect 30012 18702 30064 18708
rect 30024 18426 30052 18702
rect 28724 18420 28776 18426
rect 28724 18362 28776 18368
rect 30012 18420 30064 18426
rect 30012 18362 30064 18368
rect 30208 18290 30236 19654
rect 30760 19514 30788 20470
rect 30748 19508 30800 19514
rect 30748 19450 30800 19456
rect 30760 18698 30788 19450
rect 30748 18692 30800 18698
rect 30748 18634 30800 18640
rect 30196 18284 30248 18290
rect 30196 18226 30248 18232
rect 28080 18216 28132 18222
rect 28080 18158 28132 18164
rect 27620 18080 27672 18086
rect 27620 18022 27672 18028
rect 28397 17980 28705 17989
rect 28397 17978 28403 17980
rect 28459 17978 28483 17980
rect 28539 17978 28563 17980
rect 28619 17978 28643 17980
rect 28699 17978 28705 17980
rect 28459 17926 28461 17978
rect 28641 17926 28643 17978
rect 28397 17924 28403 17926
rect 28459 17924 28483 17926
rect 28539 17924 28563 17926
rect 28619 17924 28643 17926
rect 28699 17924 28705 17926
rect 28397 17915 28705 17924
rect 26332 17876 26384 17882
rect 26332 17818 26384 17824
rect 30208 17678 30236 18226
rect 30286 17912 30342 17921
rect 30852 17882 30880 20742
rect 31758 20703 31814 20712
rect 31668 19916 31720 19922
rect 31668 19858 31720 19864
rect 31298 19680 31354 19689
rect 31298 19615 31354 19624
rect 30286 17847 30342 17856
rect 30840 17876 30892 17882
rect 30300 17678 30328 17847
rect 30840 17818 30892 17824
rect 31312 17678 31340 19615
rect 31680 19446 31708 19858
rect 31772 19854 31800 20703
rect 32318 20700 32626 20709
rect 32318 20698 32324 20700
rect 32380 20698 32404 20700
rect 32460 20698 32484 20700
rect 32540 20698 32564 20700
rect 32620 20698 32626 20700
rect 32380 20646 32382 20698
rect 32562 20646 32564 20698
rect 32318 20644 32324 20646
rect 32380 20644 32404 20646
rect 32460 20644 32484 20646
rect 32540 20644 32564 20646
rect 32620 20644 32626 20646
rect 32318 20635 32626 20644
rect 31760 19848 31812 19854
rect 31760 19790 31812 19796
rect 32318 19612 32626 19621
rect 32318 19610 32324 19612
rect 32380 19610 32404 19612
rect 32460 19610 32484 19612
rect 32540 19610 32564 19612
rect 32620 19610 32626 19612
rect 32380 19558 32382 19610
rect 32562 19558 32564 19610
rect 32318 19556 32324 19558
rect 32380 19556 32404 19558
rect 32460 19556 32484 19558
rect 32540 19556 32564 19558
rect 32620 19556 32626 19558
rect 32318 19547 32626 19556
rect 31484 19440 31536 19446
rect 31484 19382 31536 19388
rect 31668 19440 31720 19446
rect 31668 19382 31720 19388
rect 31496 17882 31524 19382
rect 32318 18524 32626 18533
rect 32318 18522 32324 18524
rect 32380 18522 32404 18524
rect 32460 18522 32484 18524
rect 32540 18522 32564 18524
rect 32620 18522 32626 18524
rect 32380 18470 32382 18522
rect 32562 18470 32564 18522
rect 32318 18468 32324 18470
rect 32380 18468 32404 18470
rect 32460 18468 32484 18470
rect 32540 18468 32564 18470
rect 32620 18468 32626 18470
rect 32318 18459 32626 18468
rect 31484 17876 31536 17882
rect 31484 17818 31536 17824
rect 30196 17672 30248 17678
rect 30196 17614 30248 17620
rect 30288 17672 30340 17678
rect 30288 17614 30340 17620
rect 31300 17672 31352 17678
rect 31300 17614 31352 17620
rect 8792 17436 9100 17445
rect 8792 17434 8798 17436
rect 8854 17434 8878 17436
rect 8934 17434 8958 17436
rect 9014 17434 9038 17436
rect 9094 17434 9100 17436
rect 8854 17382 8856 17434
rect 9036 17382 9038 17434
rect 8792 17380 8798 17382
rect 8854 17380 8878 17382
rect 8934 17380 8958 17382
rect 9014 17380 9038 17382
rect 9094 17380 9100 17382
rect 8792 17371 9100 17380
rect 16634 17436 16942 17445
rect 16634 17434 16640 17436
rect 16696 17434 16720 17436
rect 16776 17434 16800 17436
rect 16856 17434 16880 17436
rect 16936 17434 16942 17436
rect 16696 17382 16698 17434
rect 16878 17382 16880 17434
rect 16634 17380 16640 17382
rect 16696 17380 16720 17382
rect 16776 17380 16800 17382
rect 16856 17380 16880 17382
rect 16936 17380 16942 17382
rect 16634 17371 16942 17380
rect 24476 17436 24784 17445
rect 24476 17434 24482 17436
rect 24538 17434 24562 17436
rect 24618 17434 24642 17436
rect 24698 17434 24722 17436
rect 24778 17434 24784 17436
rect 24538 17382 24540 17434
rect 24720 17382 24722 17434
rect 24476 17380 24482 17382
rect 24538 17380 24562 17382
rect 24618 17380 24642 17382
rect 24698 17380 24722 17382
rect 24778 17380 24784 17382
rect 24476 17371 24784 17380
rect 32318 17436 32626 17445
rect 32318 17434 32324 17436
rect 32380 17434 32404 17436
rect 32460 17434 32484 17436
rect 32540 17434 32564 17436
rect 32620 17434 32626 17436
rect 32380 17382 32382 17434
rect 32562 17382 32564 17434
rect 32318 17380 32324 17382
rect 32380 17380 32404 17382
rect 32460 17380 32484 17382
rect 32540 17380 32564 17382
rect 32620 17380 32626 17382
rect 32318 17371 32626 17380
rect 4871 16892 5179 16901
rect 4871 16890 4877 16892
rect 4933 16890 4957 16892
rect 5013 16890 5037 16892
rect 5093 16890 5117 16892
rect 5173 16890 5179 16892
rect 4933 16838 4935 16890
rect 5115 16838 5117 16890
rect 4871 16836 4877 16838
rect 4933 16836 4957 16838
rect 5013 16836 5037 16838
rect 5093 16836 5117 16838
rect 5173 16836 5179 16838
rect 4871 16827 5179 16836
rect 12713 16892 13021 16901
rect 12713 16890 12719 16892
rect 12775 16890 12799 16892
rect 12855 16890 12879 16892
rect 12935 16890 12959 16892
rect 13015 16890 13021 16892
rect 12775 16838 12777 16890
rect 12957 16838 12959 16890
rect 12713 16836 12719 16838
rect 12775 16836 12799 16838
rect 12855 16836 12879 16838
rect 12935 16836 12959 16838
rect 13015 16836 13021 16838
rect 12713 16827 13021 16836
rect 20555 16892 20863 16901
rect 20555 16890 20561 16892
rect 20617 16890 20641 16892
rect 20697 16890 20721 16892
rect 20777 16890 20801 16892
rect 20857 16890 20863 16892
rect 20617 16838 20619 16890
rect 20799 16838 20801 16890
rect 20555 16836 20561 16838
rect 20617 16836 20641 16838
rect 20697 16836 20721 16838
rect 20777 16836 20801 16838
rect 20857 16836 20863 16838
rect 20555 16827 20863 16836
rect 28397 16892 28705 16901
rect 28397 16890 28403 16892
rect 28459 16890 28483 16892
rect 28539 16890 28563 16892
rect 28619 16890 28643 16892
rect 28699 16890 28705 16892
rect 28459 16838 28461 16890
rect 28641 16838 28643 16890
rect 28397 16836 28403 16838
rect 28459 16836 28483 16838
rect 28539 16836 28563 16838
rect 28619 16836 28643 16838
rect 28699 16836 28705 16838
rect 28397 16827 28705 16836
rect 8792 16348 9100 16357
rect 8792 16346 8798 16348
rect 8854 16346 8878 16348
rect 8934 16346 8958 16348
rect 9014 16346 9038 16348
rect 9094 16346 9100 16348
rect 8854 16294 8856 16346
rect 9036 16294 9038 16346
rect 8792 16292 8798 16294
rect 8854 16292 8878 16294
rect 8934 16292 8958 16294
rect 9014 16292 9038 16294
rect 9094 16292 9100 16294
rect 8792 16283 9100 16292
rect 16634 16348 16942 16357
rect 16634 16346 16640 16348
rect 16696 16346 16720 16348
rect 16776 16346 16800 16348
rect 16856 16346 16880 16348
rect 16936 16346 16942 16348
rect 16696 16294 16698 16346
rect 16878 16294 16880 16346
rect 16634 16292 16640 16294
rect 16696 16292 16720 16294
rect 16776 16292 16800 16294
rect 16856 16292 16880 16294
rect 16936 16292 16942 16294
rect 16634 16283 16942 16292
rect 24476 16348 24784 16357
rect 24476 16346 24482 16348
rect 24538 16346 24562 16348
rect 24618 16346 24642 16348
rect 24698 16346 24722 16348
rect 24778 16346 24784 16348
rect 24538 16294 24540 16346
rect 24720 16294 24722 16346
rect 24476 16292 24482 16294
rect 24538 16292 24562 16294
rect 24618 16292 24642 16294
rect 24698 16292 24722 16294
rect 24778 16292 24784 16294
rect 24476 16283 24784 16292
rect 32318 16348 32626 16357
rect 32318 16346 32324 16348
rect 32380 16346 32404 16348
rect 32460 16346 32484 16348
rect 32540 16346 32564 16348
rect 32620 16346 32626 16348
rect 32380 16294 32382 16346
rect 32562 16294 32564 16346
rect 32318 16292 32324 16294
rect 32380 16292 32404 16294
rect 32460 16292 32484 16294
rect 32540 16292 32564 16294
rect 32620 16292 32626 16294
rect 32318 16283 32626 16292
rect 4871 15804 5179 15813
rect 4871 15802 4877 15804
rect 4933 15802 4957 15804
rect 5013 15802 5037 15804
rect 5093 15802 5117 15804
rect 5173 15802 5179 15804
rect 4933 15750 4935 15802
rect 5115 15750 5117 15802
rect 4871 15748 4877 15750
rect 4933 15748 4957 15750
rect 5013 15748 5037 15750
rect 5093 15748 5117 15750
rect 5173 15748 5179 15750
rect 4871 15739 5179 15748
rect 12713 15804 13021 15813
rect 12713 15802 12719 15804
rect 12775 15802 12799 15804
rect 12855 15802 12879 15804
rect 12935 15802 12959 15804
rect 13015 15802 13021 15804
rect 12775 15750 12777 15802
rect 12957 15750 12959 15802
rect 12713 15748 12719 15750
rect 12775 15748 12799 15750
rect 12855 15748 12879 15750
rect 12935 15748 12959 15750
rect 13015 15748 13021 15750
rect 12713 15739 13021 15748
rect 20555 15804 20863 15813
rect 20555 15802 20561 15804
rect 20617 15802 20641 15804
rect 20697 15802 20721 15804
rect 20777 15802 20801 15804
rect 20857 15802 20863 15804
rect 20617 15750 20619 15802
rect 20799 15750 20801 15802
rect 20555 15748 20561 15750
rect 20617 15748 20641 15750
rect 20697 15748 20721 15750
rect 20777 15748 20801 15750
rect 20857 15748 20863 15750
rect 20555 15739 20863 15748
rect 28397 15804 28705 15813
rect 28397 15802 28403 15804
rect 28459 15802 28483 15804
rect 28539 15802 28563 15804
rect 28619 15802 28643 15804
rect 28699 15802 28705 15804
rect 28459 15750 28461 15802
rect 28641 15750 28643 15802
rect 28397 15748 28403 15750
rect 28459 15748 28483 15750
rect 28539 15748 28563 15750
rect 28619 15748 28643 15750
rect 28699 15748 28705 15750
rect 28397 15739 28705 15748
rect 8792 15260 9100 15269
rect 8792 15258 8798 15260
rect 8854 15258 8878 15260
rect 8934 15258 8958 15260
rect 9014 15258 9038 15260
rect 9094 15258 9100 15260
rect 8854 15206 8856 15258
rect 9036 15206 9038 15258
rect 8792 15204 8798 15206
rect 8854 15204 8878 15206
rect 8934 15204 8958 15206
rect 9014 15204 9038 15206
rect 9094 15204 9100 15206
rect 8792 15195 9100 15204
rect 16634 15260 16942 15269
rect 16634 15258 16640 15260
rect 16696 15258 16720 15260
rect 16776 15258 16800 15260
rect 16856 15258 16880 15260
rect 16936 15258 16942 15260
rect 16696 15206 16698 15258
rect 16878 15206 16880 15258
rect 16634 15204 16640 15206
rect 16696 15204 16720 15206
rect 16776 15204 16800 15206
rect 16856 15204 16880 15206
rect 16936 15204 16942 15206
rect 16634 15195 16942 15204
rect 24476 15260 24784 15269
rect 24476 15258 24482 15260
rect 24538 15258 24562 15260
rect 24618 15258 24642 15260
rect 24698 15258 24722 15260
rect 24778 15258 24784 15260
rect 24538 15206 24540 15258
rect 24720 15206 24722 15258
rect 24476 15204 24482 15206
rect 24538 15204 24562 15206
rect 24618 15204 24642 15206
rect 24698 15204 24722 15206
rect 24778 15204 24784 15206
rect 24476 15195 24784 15204
rect 32318 15260 32626 15269
rect 32318 15258 32324 15260
rect 32380 15258 32404 15260
rect 32460 15258 32484 15260
rect 32540 15258 32564 15260
rect 32620 15258 32626 15260
rect 32380 15206 32382 15258
rect 32562 15206 32564 15258
rect 32318 15204 32324 15206
rect 32380 15204 32404 15206
rect 32460 15204 32484 15206
rect 32540 15204 32564 15206
rect 32620 15204 32626 15206
rect 32318 15195 32626 15204
rect 4871 14716 5179 14725
rect 4871 14714 4877 14716
rect 4933 14714 4957 14716
rect 5013 14714 5037 14716
rect 5093 14714 5117 14716
rect 5173 14714 5179 14716
rect 4933 14662 4935 14714
rect 5115 14662 5117 14714
rect 4871 14660 4877 14662
rect 4933 14660 4957 14662
rect 5013 14660 5037 14662
rect 5093 14660 5117 14662
rect 5173 14660 5179 14662
rect 4871 14651 5179 14660
rect 12713 14716 13021 14725
rect 12713 14714 12719 14716
rect 12775 14714 12799 14716
rect 12855 14714 12879 14716
rect 12935 14714 12959 14716
rect 13015 14714 13021 14716
rect 12775 14662 12777 14714
rect 12957 14662 12959 14714
rect 12713 14660 12719 14662
rect 12775 14660 12799 14662
rect 12855 14660 12879 14662
rect 12935 14660 12959 14662
rect 13015 14660 13021 14662
rect 12713 14651 13021 14660
rect 20555 14716 20863 14725
rect 20555 14714 20561 14716
rect 20617 14714 20641 14716
rect 20697 14714 20721 14716
rect 20777 14714 20801 14716
rect 20857 14714 20863 14716
rect 20617 14662 20619 14714
rect 20799 14662 20801 14714
rect 20555 14660 20561 14662
rect 20617 14660 20641 14662
rect 20697 14660 20721 14662
rect 20777 14660 20801 14662
rect 20857 14660 20863 14662
rect 20555 14651 20863 14660
rect 28397 14716 28705 14725
rect 28397 14714 28403 14716
rect 28459 14714 28483 14716
rect 28539 14714 28563 14716
rect 28619 14714 28643 14716
rect 28699 14714 28705 14716
rect 28459 14662 28461 14714
rect 28641 14662 28643 14714
rect 28397 14660 28403 14662
rect 28459 14660 28483 14662
rect 28539 14660 28563 14662
rect 28619 14660 28643 14662
rect 28699 14660 28705 14662
rect 28397 14651 28705 14660
rect 8792 14172 9100 14181
rect 8792 14170 8798 14172
rect 8854 14170 8878 14172
rect 8934 14170 8958 14172
rect 9014 14170 9038 14172
rect 9094 14170 9100 14172
rect 8854 14118 8856 14170
rect 9036 14118 9038 14170
rect 8792 14116 8798 14118
rect 8854 14116 8878 14118
rect 8934 14116 8958 14118
rect 9014 14116 9038 14118
rect 9094 14116 9100 14118
rect 8792 14107 9100 14116
rect 16634 14172 16942 14181
rect 16634 14170 16640 14172
rect 16696 14170 16720 14172
rect 16776 14170 16800 14172
rect 16856 14170 16880 14172
rect 16936 14170 16942 14172
rect 16696 14118 16698 14170
rect 16878 14118 16880 14170
rect 16634 14116 16640 14118
rect 16696 14116 16720 14118
rect 16776 14116 16800 14118
rect 16856 14116 16880 14118
rect 16936 14116 16942 14118
rect 16634 14107 16942 14116
rect 24476 14172 24784 14181
rect 24476 14170 24482 14172
rect 24538 14170 24562 14172
rect 24618 14170 24642 14172
rect 24698 14170 24722 14172
rect 24778 14170 24784 14172
rect 24538 14118 24540 14170
rect 24720 14118 24722 14170
rect 24476 14116 24482 14118
rect 24538 14116 24562 14118
rect 24618 14116 24642 14118
rect 24698 14116 24722 14118
rect 24778 14116 24784 14118
rect 24476 14107 24784 14116
rect 32318 14172 32626 14181
rect 32318 14170 32324 14172
rect 32380 14170 32404 14172
rect 32460 14170 32484 14172
rect 32540 14170 32564 14172
rect 32620 14170 32626 14172
rect 32380 14118 32382 14170
rect 32562 14118 32564 14170
rect 32318 14116 32324 14118
rect 32380 14116 32404 14118
rect 32460 14116 32484 14118
rect 32540 14116 32564 14118
rect 32620 14116 32626 14118
rect 32318 14107 32626 14116
rect 4871 13628 5179 13637
rect 4871 13626 4877 13628
rect 4933 13626 4957 13628
rect 5013 13626 5037 13628
rect 5093 13626 5117 13628
rect 5173 13626 5179 13628
rect 4933 13574 4935 13626
rect 5115 13574 5117 13626
rect 4871 13572 4877 13574
rect 4933 13572 4957 13574
rect 5013 13572 5037 13574
rect 5093 13572 5117 13574
rect 5173 13572 5179 13574
rect 4871 13563 5179 13572
rect 12713 13628 13021 13637
rect 12713 13626 12719 13628
rect 12775 13626 12799 13628
rect 12855 13626 12879 13628
rect 12935 13626 12959 13628
rect 13015 13626 13021 13628
rect 12775 13574 12777 13626
rect 12957 13574 12959 13626
rect 12713 13572 12719 13574
rect 12775 13572 12799 13574
rect 12855 13572 12879 13574
rect 12935 13572 12959 13574
rect 13015 13572 13021 13574
rect 12713 13563 13021 13572
rect 20555 13628 20863 13637
rect 20555 13626 20561 13628
rect 20617 13626 20641 13628
rect 20697 13626 20721 13628
rect 20777 13626 20801 13628
rect 20857 13626 20863 13628
rect 20617 13574 20619 13626
rect 20799 13574 20801 13626
rect 20555 13572 20561 13574
rect 20617 13572 20641 13574
rect 20697 13572 20721 13574
rect 20777 13572 20801 13574
rect 20857 13572 20863 13574
rect 20555 13563 20863 13572
rect 28397 13628 28705 13637
rect 28397 13626 28403 13628
rect 28459 13626 28483 13628
rect 28539 13626 28563 13628
rect 28619 13626 28643 13628
rect 28699 13626 28705 13628
rect 28459 13574 28461 13626
rect 28641 13574 28643 13626
rect 28397 13572 28403 13574
rect 28459 13572 28483 13574
rect 28539 13572 28563 13574
rect 28619 13572 28643 13574
rect 28699 13572 28705 13574
rect 28397 13563 28705 13572
rect 8792 13084 9100 13093
rect 8792 13082 8798 13084
rect 8854 13082 8878 13084
rect 8934 13082 8958 13084
rect 9014 13082 9038 13084
rect 9094 13082 9100 13084
rect 8854 13030 8856 13082
rect 9036 13030 9038 13082
rect 8792 13028 8798 13030
rect 8854 13028 8878 13030
rect 8934 13028 8958 13030
rect 9014 13028 9038 13030
rect 9094 13028 9100 13030
rect 8792 13019 9100 13028
rect 16634 13084 16942 13093
rect 16634 13082 16640 13084
rect 16696 13082 16720 13084
rect 16776 13082 16800 13084
rect 16856 13082 16880 13084
rect 16936 13082 16942 13084
rect 16696 13030 16698 13082
rect 16878 13030 16880 13082
rect 16634 13028 16640 13030
rect 16696 13028 16720 13030
rect 16776 13028 16800 13030
rect 16856 13028 16880 13030
rect 16936 13028 16942 13030
rect 16634 13019 16942 13028
rect 24476 13084 24784 13093
rect 24476 13082 24482 13084
rect 24538 13082 24562 13084
rect 24618 13082 24642 13084
rect 24698 13082 24722 13084
rect 24778 13082 24784 13084
rect 24538 13030 24540 13082
rect 24720 13030 24722 13082
rect 24476 13028 24482 13030
rect 24538 13028 24562 13030
rect 24618 13028 24642 13030
rect 24698 13028 24722 13030
rect 24778 13028 24784 13030
rect 24476 13019 24784 13028
rect 32318 13084 32626 13093
rect 32318 13082 32324 13084
rect 32380 13082 32404 13084
rect 32460 13082 32484 13084
rect 32540 13082 32564 13084
rect 32620 13082 32626 13084
rect 32380 13030 32382 13082
rect 32562 13030 32564 13082
rect 32318 13028 32324 13030
rect 32380 13028 32404 13030
rect 32460 13028 32484 13030
rect 32540 13028 32564 13030
rect 32620 13028 32626 13030
rect 32318 13019 32626 13028
rect 4871 12540 5179 12549
rect 4871 12538 4877 12540
rect 4933 12538 4957 12540
rect 5013 12538 5037 12540
rect 5093 12538 5117 12540
rect 5173 12538 5179 12540
rect 4933 12486 4935 12538
rect 5115 12486 5117 12538
rect 4871 12484 4877 12486
rect 4933 12484 4957 12486
rect 5013 12484 5037 12486
rect 5093 12484 5117 12486
rect 5173 12484 5179 12486
rect 4871 12475 5179 12484
rect 12713 12540 13021 12549
rect 12713 12538 12719 12540
rect 12775 12538 12799 12540
rect 12855 12538 12879 12540
rect 12935 12538 12959 12540
rect 13015 12538 13021 12540
rect 12775 12486 12777 12538
rect 12957 12486 12959 12538
rect 12713 12484 12719 12486
rect 12775 12484 12799 12486
rect 12855 12484 12879 12486
rect 12935 12484 12959 12486
rect 13015 12484 13021 12486
rect 12713 12475 13021 12484
rect 20555 12540 20863 12549
rect 20555 12538 20561 12540
rect 20617 12538 20641 12540
rect 20697 12538 20721 12540
rect 20777 12538 20801 12540
rect 20857 12538 20863 12540
rect 20617 12486 20619 12538
rect 20799 12486 20801 12538
rect 20555 12484 20561 12486
rect 20617 12484 20641 12486
rect 20697 12484 20721 12486
rect 20777 12484 20801 12486
rect 20857 12484 20863 12486
rect 20555 12475 20863 12484
rect 28397 12540 28705 12549
rect 28397 12538 28403 12540
rect 28459 12538 28483 12540
rect 28539 12538 28563 12540
rect 28619 12538 28643 12540
rect 28699 12538 28705 12540
rect 28459 12486 28461 12538
rect 28641 12486 28643 12538
rect 28397 12484 28403 12486
rect 28459 12484 28483 12486
rect 28539 12484 28563 12486
rect 28619 12484 28643 12486
rect 28699 12484 28705 12486
rect 28397 12475 28705 12484
rect 8792 11996 9100 12005
rect 8792 11994 8798 11996
rect 8854 11994 8878 11996
rect 8934 11994 8958 11996
rect 9014 11994 9038 11996
rect 9094 11994 9100 11996
rect 8854 11942 8856 11994
rect 9036 11942 9038 11994
rect 8792 11940 8798 11942
rect 8854 11940 8878 11942
rect 8934 11940 8958 11942
rect 9014 11940 9038 11942
rect 9094 11940 9100 11942
rect 8792 11931 9100 11940
rect 16634 11996 16942 12005
rect 16634 11994 16640 11996
rect 16696 11994 16720 11996
rect 16776 11994 16800 11996
rect 16856 11994 16880 11996
rect 16936 11994 16942 11996
rect 16696 11942 16698 11994
rect 16878 11942 16880 11994
rect 16634 11940 16640 11942
rect 16696 11940 16720 11942
rect 16776 11940 16800 11942
rect 16856 11940 16880 11942
rect 16936 11940 16942 11942
rect 16634 11931 16942 11940
rect 24476 11996 24784 12005
rect 24476 11994 24482 11996
rect 24538 11994 24562 11996
rect 24618 11994 24642 11996
rect 24698 11994 24722 11996
rect 24778 11994 24784 11996
rect 24538 11942 24540 11994
rect 24720 11942 24722 11994
rect 24476 11940 24482 11942
rect 24538 11940 24562 11942
rect 24618 11940 24642 11942
rect 24698 11940 24722 11942
rect 24778 11940 24784 11942
rect 24476 11931 24784 11940
rect 32318 11996 32626 12005
rect 32318 11994 32324 11996
rect 32380 11994 32404 11996
rect 32460 11994 32484 11996
rect 32540 11994 32564 11996
rect 32620 11994 32626 11996
rect 32380 11942 32382 11994
rect 32562 11942 32564 11994
rect 32318 11940 32324 11942
rect 32380 11940 32404 11942
rect 32460 11940 32484 11942
rect 32540 11940 32564 11942
rect 32620 11940 32626 11942
rect 32318 11931 32626 11940
rect 4871 11452 5179 11461
rect 4871 11450 4877 11452
rect 4933 11450 4957 11452
rect 5013 11450 5037 11452
rect 5093 11450 5117 11452
rect 5173 11450 5179 11452
rect 4933 11398 4935 11450
rect 5115 11398 5117 11450
rect 4871 11396 4877 11398
rect 4933 11396 4957 11398
rect 5013 11396 5037 11398
rect 5093 11396 5117 11398
rect 5173 11396 5179 11398
rect 4871 11387 5179 11396
rect 12713 11452 13021 11461
rect 12713 11450 12719 11452
rect 12775 11450 12799 11452
rect 12855 11450 12879 11452
rect 12935 11450 12959 11452
rect 13015 11450 13021 11452
rect 12775 11398 12777 11450
rect 12957 11398 12959 11450
rect 12713 11396 12719 11398
rect 12775 11396 12799 11398
rect 12855 11396 12879 11398
rect 12935 11396 12959 11398
rect 13015 11396 13021 11398
rect 12713 11387 13021 11396
rect 20555 11452 20863 11461
rect 20555 11450 20561 11452
rect 20617 11450 20641 11452
rect 20697 11450 20721 11452
rect 20777 11450 20801 11452
rect 20857 11450 20863 11452
rect 20617 11398 20619 11450
rect 20799 11398 20801 11450
rect 20555 11396 20561 11398
rect 20617 11396 20641 11398
rect 20697 11396 20721 11398
rect 20777 11396 20801 11398
rect 20857 11396 20863 11398
rect 20555 11387 20863 11396
rect 28397 11452 28705 11461
rect 28397 11450 28403 11452
rect 28459 11450 28483 11452
rect 28539 11450 28563 11452
rect 28619 11450 28643 11452
rect 28699 11450 28705 11452
rect 28459 11398 28461 11450
rect 28641 11398 28643 11450
rect 28397 11396 28403 11398
rect 28459 11396 28483 11398
rect 28539 11396 28563 11398
rect 28619 11396 28643 11398
rect 28699 11396 28705 11398
rect 28397 11387 28705 11396
rect 8792 10908 9100 10917
rect 8792 10906 8798 10908
rect 8854 10906 8878 10908
rect 8934 10906 8958 10908
rect 9014 10906 9038 10908
rect 9094 10906 9100 10908
rect 8854 10854 8856 10906
rect 9036 10854 9038 10906
rect 8792 10852 8798 10854
rect 8854 10852 8878 10854
rect 8934 10852 8958 10854
rect 9014 10852 9038 10854
rect 9094 10852 9100 10854
rect 8792 10843 9100 10852
rect 16634 10908 16942 10917
rect 16634 10906 16640 10908
rect 16696 10906 16720 10908
rect 16776 10906 16800 10908
rect 16856 10906 16880 10908
rect 16936 10906 16942 10908
rect 16696 10854 16698 10906
rect 16878 10854 16880 10906
rect 16634 10852 16640 10854
rect 16696 10852 16720 10854
rect 16776 10852 16800 10854
rect 16856 10852 16880 10854
rect 16936 10852 16942 10854
rect 16634 10843 16942 10852
rect 24476 10908 24784 10917
rect 24476 10906 24482 10908
rect 24538 10906 24562 10908
rect 24618 10906 24642 10908
rect 24698 10906 24722 10908
rect 24778 10906 24784 10908
rect 24538 10854 24540 10906
rect 24720 10854 24722 10906
rect 24476 10852 24482 10854
rect 24538 10852 24562 10854
rect 24618 10852 24642 10854
rect 24698 10852 24722 10854
rect 24778 10852 24784 10854
rect 24476 10843 24784 10852
rect 32318 10908 32626 10917
rect 32318 10906 32324 10908
rect 32380 10906 32404 10908
rect 32460 10906 32484 10908
rect 32540 10906 32564 10908
rect 32620 10906 32626 10908
rect 32380 10854 32382 10906
rect 32562 10854 32564 10906
rect 32318 10852 32324 10854
rect 32380 10852 32404 10854
rect 32460 10852 32484 10854
rect 32540 10852 32564 10854
rect 32620 10852 32626 10854
rect 32318 10843 32626 10852
rect 4871 10364 5179 10373
rect 4871 10362 4877 10364
rect 4933 10362 4957 10364
rect 5013 10362 5037 10364
rect 5093 10362 5117 10364
rect 5173 10362 5179 10364
rect 4933 10310 4935 10362
rect 5115 10310 5117 10362
rect 4871 10308 4877 10310
rect 4933 10308 4957 10310
rect 5013 10308 5037 10310
rect 5093 10308 5117 10310
rect 5173 10308 5179 10310
rect 4871 10299 5179 10308
rect 12713 10364 13021 10373
rect 12713 10362 12719 10364
rect 12775 10362 12799 10364
rect 12855 10362 12879 10364
rect 12935 10362 12959 10364
rect 13015 10362 13021 10364
rect 12775 10310 12777 10362
rect 12957 10310 12959 10362
rect 12713 10308 12719 10310
rect 12775 10308 12799 10310
rect 12855 10308 12879 10310
rect 12935 10308 12959 10310
rect 13015 10308 13021 10310
rect 12713 10299 13021 10308
rect 20555 10364 20863 10373
rect 20555 10362 20561 10364
rect 20617 10362 20641 10364
rect 20697 10362 20721 10364
rect 20777 10362 20801 10364
rect 20857 10362 20863 10364
rect 20617 10310 20619 10362
rect 20799 10310 20801 10362
rect 20555 10308 20561 10310
rect 20617 10308 20641 10310
rect 20697 10308 20721 10310
rect 20777 10308 20801 10310
rect 20857 10308 20863 10310
rect 20555 10299 20863 10308
rect 28397 10364 28705 10373
rect 28397 10362 28403 10364
rect 28459 10362 28483 10364
rect 28539 10362 28563 10364
rect 28619 10362 28643 10364
rect 28699 10362 28705 10364
rect 28459 10310 28461 10362
rect 28641 10310 28643 10362
rect 28397 10308 28403 10310
rect 28459 10308 28483 10310
rect 28539 10308 28563 10310
rect 28619 10308 28643 10310
rect 28699 10308 28705 10310
rect 28397 10299 28705 10308
rect 8792 9820 9100 9829
rect 8792 9818 8798 9820
rect 8854 9818 8878 9820
rect 8934 9818 8958 9820
rect 9014 9818 9038 9820
rect 9094 9818 9100 9820
rect 8854 9766 8856 9818
rect 9036 9766 9038 9818
rect 8792 9764 8798 9766
rect 8854 9764 8878 9766
rect 8934 9764 8958 9766
rect 9014 9764 9038 9766
rect 9094 9764 9100 9766
rect 8792 9755 9100 9764
rect 16634 9820 16942 9829
rect 16634 9818 16640 9820
rect 16696 9818 16720 9820
rect 16776 9818 16800 9820
rect 16856 9818 16880 9820
rect 16936 9818 16942 9820
rect 16696 9766 16698 9818
rect 16878 9766 16880 9818
rect 16634 9764 16640 9766
rect 16696 9764 16720 9766
rect 16776 9764 16800 9766
rect 16856 9764 16880 9766
rect 16936 9764 16942 9766
rect 16634 9755 16942 9764
rect 24476 9820 24784 9829
rect 24476 9818 24482 9820
rect 24538 9818 24562 9820
rect 24618 9818 24642 9820
rect 24698 9818 24722 9820
rect 24778 9818 24784 9820
rect 24538 9766 24540 9818
rect 24720 9766 24722 9818
rect 24476 9764 24482 9766
rect 24538 9764 24562 9766
rect 24618 9764 24642 9766
rect 24698 9764 24722 9766
rect 24778 9764 24784 9766
rect 24476 9755 24784 9764
rect 32318 9820 32626 9829
rect 32318 9818 32324 9820
rect 32380 9818 32404 9820
rect 32460 9818 32484 9820
rect 32540 9818 32564 9820
rect 32620 9818 32626 9820
rect 32380 9766 32382 9818
rect 32562 9766 32564 9818
rect 32318 9764 32324 9766
rect 32380 9764 32404 9766
rect 32460 9764 32484 9766
rect 32540 9764 32564 9766
rect 32620 9764 32626 9766
rect 32318 9755 32626 9764
rect 4871 9276 5179 9285
rect 4871 9274 4877 9276
rect 4933 9274 4957 9276
rect 5013 9274 5037 9276
rect 5093 9274 5117 9276
rect 5173 9274 5179 9276
rect 4933 9222 4935 9274
rect 5115 9222 5117 9274
rect 4871 9220 4877 9222
rect 4933 9220 4957 9222
rect 5013 9220 5037 9222
rect 5093 9220 5117 9222
rect 5173 9220 5179 9222
rect 4871 9211 5179 9220
rect 12713 9276 13021 9285
rect 12713 9274 12719 9276
rect 12775 9274 12799 9276
rect 12855 9274 12879 9276
rect 12935 9274 12959 9276
rect 13015 9274 13021 9276
rect 12775 9222 12777 9274
rect 12957 9222 12959 9274
rect 12713 9220 12719 9222
rect 12775 9220 12799 9222
rect 12855 9220 12879 9222
rect 12935 9220 12959 9222
rect 13015 9220 13021 9222
rect 12713 9211 13021 9220
rect 20555 9276 20863 9285
rect 20555 9274 20561 9276
rect 20617 9274 20641 9276
rect 20697 9274 20721 9276
rect 20777 9274 20801 9276
rect 20857 9274 20863 9276
rect 20617 9222 20619 9274
rect 20799 9222 20801 9274
rect 20555 9220 20561 9222
rect 20617 9220 20641 9222
rect 20697 9220 20721 9222
rect 20777 9220 20801 9222
rect 20857 9220 20863 9222
rect 20555 9211 20863 9220
rect 28397 9276 28705 9285
rect 28397 9274 28403 9276
rect 28459 9274 28483 9276
rect 28539 9274 28563 9276
rect 28619 9274 28643 9276
rect 28699 9274 28705 9276
rect 28459 9222 28461 9274
rect 28641 9222 28643 9274
rect 28397 9220 28403 9222
rect 28459 9220 28483 9222
rect 28539 9220 28563 9222
rect 28619 9220 28643 9222
rect 28699 9220 28705 9222
rect 28397 9211 28705 9220
rect 8792 8732 9100 8741
rect 8792 8730 8798 8732
rect 8854 8730 8878 8732
rect 8934 8730 8958 8732
rect 9014 8730 9038 8732
rect 9094 8730 9100 8732
rect 8854 8678 8856 8730
rect 9036 8678 9038 8730
rect 8792 8676 8798 8678
rect 8854 8676 8878 8678
rect 8934 8676 8958 8678
rect 9014 8676 9038 8678
rect 9094 8676 9100 8678
rect 8792 8667 9100 8676
rect 16634 8732 16942 8741
rect 16634 8730 16640 8732
rect 16696 8730 16720 8732
rect 16776 8730 16800 8732
rect 16856 8730 16880 8732
rect 16936 8730 16942 8732
rect 16696 8678 16698 8730
rect 16878 8678 16880 8730
rect 16634 8676 16640 8678
rect 16696 8676 16720 8678
rect 16776 8676 16800 8678
rect 16856 8676 16880 8678
rect 16936 8676 16942 8678
rect 16634 8667 16942 8676
rect 24476 8732 24784 8741
rect 24476 8730 24482 8732
rect 24538 8730 24562 8732
rect 24618 8730 24642 8732
rect 24698 8730 24722 8732
rect 24778 8730 24784 8732
rect 24538 8678 24540 8730
rect 24720 8678 24722 8730
rect 24476 8676 24482 8678
rect 24538 8676 24562 8678
rect 24618 8676 24642 8678
rect 24698 8676 24722 8678
rect 24778 8676 24784 8678
rect 24476 8667 24784 8676
rect 32318 8732 32626 8741
rect 32318 8730 32324 8732
rect 32380 8730 32404 8732
rect 32460 8730 32484 8732
rect 32540 8730 32564 8732
rect 32620 8730 32626 8732
rect 32380 8678 32382 8730
rect 32562 8678 32564 8730
rect 32318 8676 32324 8678
rect 32380 8676 32404 8678
rect 32460 8676 32484 8678
rect 32540 8676 32564 8678
rect 32620 8676 32626 8678
rect 32318 8667 32626 8676
rect 4871 8188 5179 8197
rect 4871 8186 4877 8188
rect 4933 8186 4957 8188
rect 5013 8186 5037 8188
rect 5093 8186 5117 8188
rect 5173 8186 5179 8188
rect 4933 8134 4935 8186
rect 5115 8134 5117 8186
rect 4871 8132 4877 8134
rect 4933 8132 4957 8134
rect 5013 8132 5037 8134
rect 5093 8132 5117 8134
rect 5173 8132 5179 8134
rect 4871 8123 5179 8132
rect 12713 8188 13021 8197
rect 12713 8186 12719 8188
rect 12775 8186 12799 8188
rect 12855 8186 12879 8188
rect 12935 8186 12959 8188
rect 13015 8186 13021 8188
rect 12775 8134 12777 8186
rect 12957 8134 12959 8186
rect 12713 8132 12719 8134
rect 12775 8132 12799 8134
rect 12855 8132 12879 8134
rect 12935 8132 12959 8134
rect 13015 8132 13021 8134
rect 12713 8123 13021 8132
rect 20555 8188 20863 8197
rect 20555 8186 20561 8188
rect 20617 8186 20641 8188
rect 20697 8186 20721 8188
rect 20777 8186 20801 8188
rect 20857 8186 20863 8188
rect 20617 8134 20619 8186
rect 20799 8134 20801 8186
rect 20555 8132 20561 8134
rect 20617 8132 20641 8134
rect 20697 8132 20721 8134
rect 20777 8132 20801 8134
rect 20857 8132 20863 8134
rect 20555 8123 20863 8132
rect 28397 8188 28705 8197
rect 28397 8186 28403 8188
rect 28459 8186 28483 8188
rect 28539 8186 28563 8188
rect 28619 8186 28643 8188
rect 28699 8186 28705 8188
rect 28459 8134 28461 8186
rect 28641 8134 28643 8186
rect 28397 8132 28403 8134
rect 28459 8132 28483 8134
rect 28539 8132 28563 8134
rect 28619 8132 28643 8134
rect 28699 8132 28705 8134
rect 28397 8123 28705 8132
rect 8792 7644 9100 7653
rect 8792 7642 8798 7644
rect 8854 7642 8878 7644
rect 8934 7642 8958 7644
rect 9014 7642 9038 7644
rect 9094 7642 9100 7644
rect 8854 7590 8856 7642
rect 9036 7590 9038 7642
rect 8792 7588 8798 7590
rect 8854 7588 8878 7590
rect 8934 7588 8958 7590
rect 9014 7588 9038 7590
rect 9094 7588 9100 7590
rect 8792 7579 9100 7588
rect 16634 7644 16942 7653
rect 16634 7642 16640 7644
rect 16696 7642 16720 7644
rect 16776 7642 16800 7644
rect 16856 7642 16880 7644
rect 16936 7642 16942 7644
rect 16696 7590 16698 7642
rect 16878 7590 16880 7642
rect 16634 7588 16640 7590
rect 16696 7588 16720 7590
rect 16776 7588 16800 7590
rect 16856 7588 16880 7590
rect 16936 7588 16942 7590
rect 16634 7579 16942 7588
rect 24476 7644 24784 7653
rect 24476 7642 24482 7644
rect 24538 7642 24562 7644
rect 24618 7642 24642 7644
rect 24698 7642 24722 7644
rect 24778 7642 24784 7644
rect 24538 7590 24540 7642
rect 24720 7590 24722 7642
rect 24476 7588 24482 7590
rect 24538 7588 24562 7590
rect 24618 7588 24642 7590
rect 24698 7588 24722 7590
rect 24778 7588 24784 7590
rect 24476 7579 24784 7588
rect 32318 7644 32626 7653
rect 32318 7642 32324 7644
rect 32380 7642 32404 7644
rect 32460 7642 32484 7644
rect 32540 7642 32564 7644
rect 32620 7642 32626 7644
rect 32380 7590 32382 7642
rect 32562 7590 32564 7642
rect 32318 7588 32324 7590
rect 32380 7588 32404 7590
rect 32460 7588 32484 7590
rect 32540 7588 32564 7590
rect 32620 7588 32626 7590
rect 32318 7579 32626 7588
rect 4871 7100 5179 7109
rect 4871 7098 4877 7100
rect 4933 7098 4957 7100
rect 5013 7098 5037 7100
rect 5093 7098 5117 7100
rect 5173 7098 5179 7100
rect 4933 7046 4935 7098
rect 5115 7046 5117 7098
rect 4871 7044 4877 7046
rect 4933 7044 4957 7046
rect 5013 7044 5037 7046
rect 5093 7044 5117 7046
rect 5173 7044 5179 7046
rect 4871 7035 5179 7044
rect 12713 7100 13021 7109
rect 12713 7098 12719 7100
rect 12775 7098 12799 7100
rect 12855 7098 12879 7100
rect 12935 7098 12959 7100
rect 13015 7098 13021 7100
rect 12775 7046 12777 7098
rect 12957 7046 12959 7098
rect 12713 7044 12719 7046
rect 12775 7044 12799 7046
rect 12855 7044 12879 7046
rect 12935 7044 12959 7046
rect 13015 7044 13021 7046
rect 12713 7035 13021 7044
rect 20555 7100 20863 7109
rect 20555 7098 20561 7100
rect 20617 7098 20641 7100
rect 20697 7098 20721 7100
rect 20777 7098 20801 7100
rect 20857 7098 20863 7100
rect 20617 7046 20619 7098
rect 20799 7046 20801 7098
rect 20555 7044 20561 7046
rect 20617 7044 20641 7046
rect 20697 7044 20721 7046
rect 20777 7044 20801 7046
rect 20857 7044 20863 7046
rect 20555 7035 20863 7044
rect 28397 7100 28705 7109
rect 28397 7098 28403 7100
rect 28459 7098 28483 7100
rect 28539 7098 28563 7100
rect 28619 7098 28643 7100
rect 28699 7098 28705 7100
rect 28459 7046 28461 7098
rect 28641 7046 28643 7098
rect 28397 7044 28403 7046
rect 28459 7044 28483 7046
rect 28539 7044 28563 7046
rect 28619 7044 28643 7046
rect 28699 7044 28705 7046
rect 28397 7035 28705 7044
rect 8792 6556 9100 6565
rect 8792 6554 8798 6556
rect 8854 6554 8878 6556
rect 8934 6554 8958 6556
rect 9014 6554 9038 6556
rect 9094 6554 9100 6556
rect 8854 6502 8856 6554
rect 9036 6502 9038 6554
rect 8792 6500 8798 6502
rect 8854 6500 8878 6502
rect 8934 6500 8958 6502
rect 9014 6500 9038 6502
rect 9094 6500 9100 6502
rect 8792 6491 9100 6500
rect 16634 6556 16942 6565
rect 16634 6554 16640 6556
rect 16696 6554 16720 6556
rect 16776 6554 16800 6556
rect 16856 6554 16880 6556
rect 16936 6554 16942 6556
rect 16696 6502 16698 6554
rect 16878 6502 16880 6554
rect 16634 6500 16640 6502
rect 16696 6500 16720 6502
rect 16776 6500 16800 6502
rect 16856 6500 16880 6502
rect 16936 6500 16942 6502
rect 16634 6491 16942 6500
rect 24476 6556 24784 6565
rect 24476 6554 24482 6556
rect 24538 6554 24562 6556
rect 24618 6554 24642 6556
rect 24698 6554 24722 6556
rect 24778 6554 24784 6556
rect 24538 6502 24540 6554
rect 24720 6502 24722 6554
rect 24476 6500 24482 6502
rect 24538 6500 24562 6502
rect 24618 6500 24642 6502
rect 24698 6500 24722 6502
rect 24778 6500 24784 6502
rect 24476 6491 24784 6500
rect 32318 6556 32626 6565
rect 32318 6554 32324 6556
rect 32380 6554 32404 6556
rect 32460 6554 32484 6556
rect 32540 6554 32564 6556
rect 32620 6554 32626 6556
rect 32380 6502 32382 6554
rect 32562 6502 32564 6554
rect 32318 6500 32324 6502
rect 32380 6500 32404 6502
rect 32460 6500 32484 6502
rect 32540 6500 32564 6502
rect 32620 6500 32626 6502
rect 32318 6491 32626 6500
rect 4871 6012 5179 6021
rect 4871 6010 4877 6012
rect 4933 6010 4957 6012
rect 5013 6010 5037 6012
rect 5093 6010 5117 6012
rect 5173 6010 5179 6012
rect 4933 5958 4935 6010
rect 5115 5958 5117 6010
rect 4871 5956 4877 5958
rect 4933 5956 4957 5958
rect 5013 5956 5037 5958
rect 5093 5956 5117 5958
rect 5173 5956 5179 5958
rect 4871 5947 5179 5956
rect 12713 6012 13021 6021
rect 12713 6010 12719 6012
rect 12775 6010 12799 6012
rect 12855 6010 12879 6012
rect 12935 6010 12959 6012
rect 13015 6010 13021 6012
rect 12775 5958 12777 6010
rect 12957 5958 12959 6010
rect 12713 5956 12719 5958
rect 12775 5956 12799 5958
rect 12855 5956 12879 5958
rect 12935 5956 12959 5958
rect 13015 5956 13021 5958
rect 12713 5947 13021 5956
rect 20555 6012 20863 6021
rect 20555 6010 20561 6012
rect 20617 6010 20641 6012
rect 20697 6010 20721 6012
rect 20777 6010 20801 6012
rect 20857 6010 20863 6012
rect 20617 5958 20619 6010
rect 20799 5958 20801 6010
rect 20555 5956 20561 5958
rect 20617 5956 20641 5958
rect 20697 5956 20721 5958
rect 20777 5956 20801 5958
rect 20857 5956 20863 5958
rect 20555 5947 20863 5956
rect 28397 6012 28705 6021
rect 28397 6010 28403 6012
rect 28459 6010 28483 6012
rect 28539 6010 28563 6012
rect 28619 6010 28643 6012
rect 28699 6010 28705 6012
rect 28459 5958 28461 6010
rect 28641 5958 28643 6010
rect 28397 5956 28403 5958
rect 28459 5956 28483 5958
rect 28539 5956 28563 5958
rect 28619 5956 28643 5958
rect 28699 5956 28705 5958
rect 28397 5947 28705 5956
rect 8792 5468 9100 5477
rect 8792 5466 8798 5468
rect 8854 5466 8878 5468
rect 8934 5466 8958 5468
rect 9014 5466 9038 5468
rect 9094 5466 9100 5468
rect 8854 5414 8856 5466
rect 9036 5414 9038 5466
rect 8792 5412 8798 5414
rect 8854 5412 8878 5414
rect 8934 5412 8958 5414
rect 9014 5412 9038 5414
rect 9094 5412 9100 5414
rect 8792 5403 9100 5412
rect 16634 5468 16942 5477
rect 16634 5466 16640 5468
rect 16696 5466 16720 5468
rect 16776 5466 16800 5468
rect 16856 5466 16880 5468
rect 16936 5466 16942 5468
rect 16696 5414 16698 5466
rect 16878 5414 16880 5466
rect 16634 5412 16640 5414
rect 16696 5412 16720 5414
rect 16776 5412 16800 5414
rect 16856 5412 16880 5414
rect 16936 5412 16942 5414
rect 16634 5403 16942 5412
rect 24476 5468 24784 5477
rect 24476 5466 24482 5468
rect 24538 5466 24562 5468
rect 24618 5466 24642 5468
rect 24698 5466 24722 5468
rect 24778 5466 24784 5468
rect 24538 5414 24540 5466
rect 24720 5414 24722 5466
rect 24476 5412 24482 5414
rect 24538 5412 24562 5414
rect 24618 5412 24642 5414
rect 24698 5412 24722 5414
rect 24778 5412 24784 5414
rect 24476 5403 24784 5412
rect 32318 5468 32626 5477
rect 32318 5466 32324 5468
rect 32380 5466 32404 5468
rect 32460 5466 32484 5468
rect 32540 5466 32564 5468
rect 32620 5466 32626 5468
rect 32380 5414 32382 5466
rect 32562 5414 32564 5466
rect 32318 5412 32324 5414
rect 32380 5412 32404 5414
rect 32460 5412 32484 5414
rect 32540 5412 32564 5414
rect 32620 5412 32626 5414
rect 32318 5403 32626 5412
rect 4871 4924 5179 4933
rect 4871 4922 4877 4924
rect 4933 4922 4957 4924
rect 5013 4922 5037 4924
rect 5093 4922 5117 4924
rect 5173 4922 5179 4924
rect 4933 4870 4935 4922
rect 5115 4870 5117 4922
rect 4871 4868 4877 4870
rect 4933 4868 4957 4870
rect 5013 4868 5037 4870
rect 5093 4868 5117 4870
rect 5173 4868 5179 4870
rect 4871 4859 5179 4868
rect 12713 4924 13021 4933
rect 12713 4922 12719 4924
rect 12775 4922 12799 4924
rect 12855 4922 12879 4924
rect 12935 4922 12959 4924
rect 13015 4922 13021 4924
rect 12775 4870 12777 4922
rect 12957 4870 12959 4922
rect 12713 4868 12719 4870
rect 12775 4868 12799 4870
rect 12855 4868 12879 4870
rect 12935 4868 12959 4870
rect 13015 4868 13021 4870
rect 12713 4859 13021 4868
rect 20555 4924 20863 4933
rect 20555 4922 20561 4924
rect 20617 4922 20641 4924
rect 20697 4922 20721 4924
rect 20777 4922 20801 4924
rect 20857 4922 20863 4924
rect 20617 4870 20619 4922
rect 20799 4870 20801 4922
rect 20555 4868 20561 4870
rect 20617 4868 20641 4870
rect 20697 4868 20721 4870
rect 20777 4868 20801 4870
rect 20857 4868 20863 4870
rect 20555 4859 20863 4868
rect 28397 4924 28705 4933
rect 28397 4922 28403 4924
rect 28459 4922 28483 4924
rect 28539 4922 28563 4924
rect 28619 4922 28643 4924
rect 28699 4922 28705 4924
rect 28459 4870 28461 4922
rect 28641 4870 28643 4922
rect 28397 4868 28403 4870
rect 28459 4868 28483 4870
rect 28539 4868 28563 4870
rect 28619 4868 28643 4870
rect 28699 4868 28705 4870
rect 28397 4859 28705 4868
rect 8792 4380 9100 4389
rect 8792 4378 8798 4380
rect 8854 4378 8878 4380
rect 8934 4378 8958 4380
rect 9014 4378 9038 4380
rect 9094 4378 9100 4380
rect 8854 4326 8856 4378
rect 9036 4326 9038 4378
rect 8792 4324 8798 4326
rect 8854 4324 8878 4326
rect 8934 4324 8958 4326
rect 9014 4324 9038 4326
rect 9094 4324 9100 4326
rect 8792 4315 9100 4324
rect 16634 4380 16942 4389
rect 16634 4378 16640 4380
rect 16696 4378 16720 4380
rect 16776 4378 16800 4380
rect 16856 4378 16880 4380
rect 16936 4378 16942 4380
rect 16696 4326 16698 4378
rect 16878 4326 16880 4378
rect 16634 4324 16640 4326
rect 16696 4324 16720 4326
rect 16776 4324 16800 4326
rect 16856 4324 16880 4326
rect 16936 4324 16942 4326
rect 16634 4315 16942 4324
rect 24476 4380 24784 4389
rect 24476 4378 24482 4380
rect 24538 4378 24562 4380
rect 24618 4378 24642 4380
rect 24698 4378 24722 4380
rect 24778 4378 24784 4380
rect 24538 4326 24540 4378
rect 24720 4326 24722 4378
rect 24476 4324 24482 4326
rect 24538 4324 24562 4326
rect 24618 4324 24642 4326
rect 24698 4324 24722 4326
rect 24778 4324 24784 4326
rect 24476 4315 24784 4324
rect 32318 4380 32626 4389
rect 32318 4378 32324 4380
rect 32380 4378 32404 4380
rect 32460 4378 32484 4380
rect 32540 4378 32564 4380
rect 32620 4378 32626 4380
rect 32380 4326 32382 4378
rect 32562 4326 32564 4378
rect 32318 4324 32324 4326
rect 32380 4324 32404 4326
rect 32460 4324 32484 4326
rect 32540 4324 32564 4326
rect 32620 4324 32626 4326
rect 32318 4315 32626 4324
rect 4871 3836 5179 3845
rect 4871 3834 4877 3836
rect 4933 3834 4957 3836
rect 5013 3834 5037 3836
rect 5093 3834 5117 3836
rect 5173 3834 5179 3836
rect 4933 3782 4935 3834
rect 5115 3782 5117 3834
rect 4871 3780 4877 3782
rect 4933 3780 4957 3782
rect 5013 3780 5037 3782
rect 5093 3780 5117 3782
rect 5173 3780 5179 3782
rect 4871 3771 5179 3780
rect 12713 3836 13021 3845
rect 12713 3834 12719 3836
rect 12775 3834 12799 3836
rect 12855 3834 12879 3836
rect 12935 3834 12959 3836
rect 13015 3834 13021 3836
rect 12775 3782 12777 3834
rect 12957 3782 12959 3834
rect 12713 3780 12719 3782
rect 12775 3780 12799 3782
rect 12855 3780 12879 3782
rect 12935 3780 12959 3782
rect 13015 3780 13021 3782
rect 12713 3771 13021 3780
rect 20555 3836 20863 3845
rect 20555 3834 20561 3836
rect 20617 3834 20641 3836
rect 20697 3834 20721 3836
rect 20777 3834 20801 3836
rect 20857 3834 20863 3836
rect 20617 3782 20619 3834
rect 20799 3782 20801 3834
rect 20555 3780 20561 3782
rect 20617 3780 20641 3782
rect 20697 3780 20721 3782
rect 20777 3780 20801 3782
rect 20857 3780 20863 3782
rect 20555 3771 20863 3780
rect 28397 3836 28705 3845
rect 28397 3834 28403 3836
rect 28459 3834 28483 3836
rect 28539 3834 28563 3836
rect 28619 3834 28643 3836
rect 28699 3834 28705 3836
rect 28459 3782 28461 3834
rect 28641 3782 28643 3834
rect 28397 3780 28403 3782
rect 28459 3780 28483 3782
rect 28539 3780 28563 3782
rect 28619 3780 28643 3782
rect 28699 3780 28705 3782
rect 28397 3771 28705 3780
rect 8792 3292 9100 3301
rect 8792 3290 8798 3292
rect 8854 3290 8878 3292
rect 8934 3290 8958 3292
rect 9014 3290 9038 3292
rect 9094 3290 9100 3292
rect 8854 3238 8856 3290
rect 9036 3238 9038 3290
rect 8792 3236 8798 3238
rect 8854 3236 8878 3238
rect 8934 3236 8958 3238
rect 9014 3236 9038 3238
rect 9094 3236 9100 3238
rect 8792 3227 9100 3236
rect 16634 3292 16942 3301
rect 16634 3290 16640 3292
rect 16696 3290 16720 3292
rect 16776 3290 16800 3292
rect 16856 3290 16880 3292
rect 16936 3290 16942 3292
rect 16696 3238 16698 3290
rect 16878 3238 16880 3290
rect 16634 3236 16640 3238
rect 16696 3236 16720 3238
rect 16776 3236 16800 3238
rect 16856 3236 16880 3238
rect 16936 3236 16942 3238
rect 16634 3227 16942 3236
rect 24476 3292 24784 3301
rect 24476 3290 24482 3292
rect 24538 3290 24562 3292
rect 24618 3290 24642 3292
rect 24698 3290 24722 3292
rect 24778 3290 24784 3292
rect 24538 3238 24540 3290
rect 24720 3238 24722 3290
rect 24476 3236 24482 3238
rect 24538 3236 24562 3238
rect 24618 3236 24642 3238
rect 24698 3236 24722 3238
rect 24778 3236 24784 3238
rect 24476 3227 24784 3236
rect 32318 3292 32626 3301
rect 32318 3290 32324 3292
rect 32380 3290 32404 3292
rect 32460 3290 32484 3292
rect 32540 3290 32564 3292
rect 32620 3290 32626 3292
rect 32380 3238 32382 3290
rect 32562 3238 32564 3290
rect 32318 3236 32324 3238
rect 32380 3236 32404 3238
rect 32460 3236 32484 3238
rect 32540 3236 32564 3238
rect 32620 3236 32626 3238
rect 32318 3227 32626 3236
rect 4871 2748 5179 2757
rect 4871 2746 4877 2748
rect 4933 2746 4957 2748
rect 5013 2746 5037 2748
rect 5093 2746 5117 2748
rect 5173 2746 5179 2748
rect 4933 2694 4935 2746
rect 5115 2694 5117 2746
rect 4871 2692 4877 2694
rect 4933 2692 4957 2694
rect 5013 2692 5037 2694
rect 5093 2692 5117 2694
rect 5173 2692 5179 2694
rect 4871 2683 5179 2692
rect 12713 2748 13021 2757
rect 12713 2746 12719 2748
rect 12775 2746 12799 2748
rect 12855 2746 12879 2748
rect 12935 2746 12959 2748
rect 13015 2746 13021 2748
rect 12775 2694 12777 2746
rect 12957 2694 12959 2746
rect 12713 2692 12719 2694
rect 12775 2692 12799 2694
rect 12855 2692 12879 2694
rect 12935 2692 12959 2694
rect 13015 2692 13021 2694
rect 12713 2683 13021 2692
rect 20555 2748 20863 2757
rect 20555 2746 20561 2748
rect 20617 2746 20641 2748
rect 20697 2746 20721 2748
rect 20777 2746 20801 2748
rect 20857 2746 20863 2748
rect 20617 2694 20619 2746
rect 20799 2694 20801 2746
rect 20555 2692 20561 2694
rect 20617 2692 20641 2694
rect 20697 2692 20721 2694
rect 20777 2692 20801 2694
rect 20857 2692 20863 2694
rect 20555 2683 20863 2692
rect 28397 2748 28705 2757
rect 28397 2746 28403 2748
rect 28459 2746 28483 2748
rect 28539 2746 28563 2748
rect 28619 2746 28643 2748
rect 28699 2746 28705 2748
rect 28459 2694 28461 2746
rect 28641 2694 28643 2746
rect 28397 2692 28403 2694
rect 28459 2692 28483 2694
rect 28539 2692 28563 2694
rect 28619 2692 28643 2694
rect 28699 2692 28705 2694
rect 28397 2683 28705 2692
rect 8792 2204 9100 2213
rect 8792 2202 8798 2204
rect 8854 2202 8878 2204
rect 8934 2202 8958 2204
rect 9014 2202 9038 2204
rect 9094 2202 9100 2204
rect 8854 2150 8856 2202
rect 9036 2150 9038 2202
rect 8792 2148 8798 2150
rect 8854 2148 8878 2150
rect 8934 2148 8958 2150
rect 9014 2148 9038 2150
rect 9094 2148 9100 2150
rect 8792 2139 9100 2148
rect 16634 2204 16942 2213
rect 16634 2202 16640 2204
rect 16696 2202 16720 2204
rect 16776 2202 16800 2204
rect 16856 2202 16880 2204
rect 16936 2202 16942 2204
rect 16696 2150 16698 2202
rect 16878 2150 16880 2202
rect 16634 2148 16640 2150
rect 16696 2148 16720 2150
rect 16776 2148 16800 2150
rect 16856 2148 16880 2150
rect 16936 2148 16942 2150
rect 16634 2139 16942 2148
rect 24476 2204 24784 2213
rect 24476 2202 24482 2204
rect 24538 2202 24562 2204
rect 24618 2202 24642 2204
rect 24698 2202 24722 2204
rect 24778 2202 24784 2204
rect 24538 2150 24540 2202
rect 24720 2150 24722 2202
rect 24476 2148 24482 2150
rect 24538 2148 24562 2150
rect 24618 2148 24642 2150
rect 24698 2148 24722 2150
rect 24778 2148 24784 2150
rect 24476 2139 24784 2148
rect 32318 2204 32626 2213
rect 32318 2202 32324 2204
rect 32380 2202 32404 2204
rect 32460 2202 32484 2204
rect 32540 2202 32564 2204
rect 32620 2202 32626 2204
rect 32380 2150 32382 2202
rect 32562 2150 32564 2202
rect 32318 2148 32324 2150
rect 32380 2148 32404 2150
rect 32460 2148 32484 2150
rect 32540 2148 32564 2150
rect 32620 2148 32626 2150
rect 32318 2139 32626 2148
rect 4871 1660 5179 1669
rect 4871 1658 4877 1660
rect 4933 1658 4957 1660
rect 5013 1658 5037 1660
rect 5093 1658 5117 1660
rect 5173 1658 5179 1660
rect 4933 1606 4935 1658
rect 5115 1606 5117 1658
rect 4871 1604 4877 1606
rect 4933 1604 4957 1606
rect 5013 1604 5037 1606
rect 5093 1604 5117 1606
rect 5173 1604 5179 1606
rect 4871 1595 5179 1604
rect 12713 1660 13021 1669
rect 12713 1658 12719 1660
rect 12775 1658 12799 1660
rect 12855 1658 12879 1660
rect 12935 1658 12959 1660
rect 13015 1658 13021 1660
rect 12775 1606 12777 1658
rect 12957 1606 12959 1658
rect 12713 1604 12719 1606
rect 12775 1604 12799 1606
rect 12855 1604 12879 1606
rect 12935 1604 12959 1606
rect 13015 1604 13021 1606
rect 12713 1595 13021 1604
rect 20555 1660 20863 1669
rect 20555 1658 20561 1660
rect 20617 1658 20641 1660
rect 20697 1658 20721 1660
rect 20777 1658 20801 1660
rect 20857 1658 20863 1660
rect 20617 1606 20619 1658
rect 20799 1606 20801 1658
rect 20555 1604 20561 1606
rect 20617 1604 20641 1606
rect 20697 1604 20721 1606
rect 20777 1604 20801 1606
rect 20857 1604 20863 1606
rect 20555 1595 20863 1604
rect 28397 1660 28705 1669
rect 28397 1658 28403 1660
rect 28459 1658 28483 1660
rect 28539 1658 28563 1660
rect 28619 1658 28643 1660
rect 28699 1658 28705 1660
rect 28459 1606 28461 1658
rect 28641 1606 28643 1658
rect 28397 1604 28403 1606
rect 28459 1604 28483 1606
rect 28539 1604 28563 1606
rect 28619 1604 28643 1606
rect 28699 1604 28705 1606
rect 28397 1595 28705 1604
rect 8792 1116 9100 1125
rect 8792 1114 8798 1116
rect 8854 1114 8878 1116
rect 8934 1114 8958 1116
rect 9014 1114 9038 1116
rect 9094 1114 9100 1116
rect 8854 1062 8856 1114
rect 9036 1062 9038 1114
rect 8792 1060 8798 1062
rect 8854 1060 8878 1062
rect 8934 1060 8958 1062
rect 9014 1060 9038 1062
rect 9094 1060 9100 1062
rect 8792 1051 9100 1060
rect 16634 1116 16942 1125
rect 16634 1114 16640 1116
rect 16696 1114 16720 1116
rect 16776 1114 16800 1116
rect 16856 1114 16880 1116
rect 16936 1114 16942 1116
rect 16696 1062 16698 1114
rect 16878 1062 16880 1114
rect 16634 1060 16640 1062
rect 16696 1060 16720 1062
rect 16776 1060 16800 1062
rect 16856 1060 16880 1062
rect 16936 1060 16942 1062
rect 16634 1051 16942 1060
rect 24476 1116 24784 1125
rect 24476 1114 24482 1116
rect 24538 1114 24562 1116
rect 24618 1114 24642 1116
rect 24698 1114 24722 1116
rect 24778 1114 24784 1116
rect 24538 1062 24540 1114
rect 24720 1062 24722 1114
rect 24476 1060 24482 1062
rect 24538 1060 24562 1062
rect 24618 1060 24642 1062
rect 24698 1060 24722 1062
rect 24778 1060 24784 1062
rect 24476 1051 24784 1060
rect 32318 1116 32626 1125
rect 32318 1114 32324 1116
rect 32380 1114 32404 1116
rect 32460 1114 32484 1116
rect 32540 1114 32564 1116
rect 32620 1114 32626 1116
rect 32380 1062 32382 1114
rect 32562 1062 32564 1114
rect 32318 1060 32324 1062
rect 32380 1060 32404 1062
rect 32460 1060 32484 1062
rect 32540 1060 32564 1062
rect 32620 1060 32626 1062
rect 32318 1051 32626 1060
<< via2 >>
rect 19982 21120 20038 21176
rect 23662 21120 23718 21176
rect 5262 20848 5318 20904
rect 9126 20848 9182 20904
rect 17774 20848 17830 20904
rect 4877 20154 4933 20156
rect 4957 20154 5013 20156
rect 5037 20154 5093 20156
rect 5117 20154 5173 20156
rect 4877 20102 4923 20154
rect 4923 20102 4933 20154
rect 4957 20102 4987 20154
rect 4987 20102 4999 20154
rect 4999 20102 5013 20154
rect 5037 20102 5051 20154
rect 5051 20102 5063 20154
rect 5063 20102 5093 20154
rect 5117 20102 5127 20154
rect 5127 20102 5173 20154
rect 4877 20100 4933 20102
rect 4957 20100 5013 20102
rect 5037 20100 5093 20102
rect 5117 20100 5173 20102
rect 2226 20052 2282 20088
rect 2226 20032 2228 20052
rect 2228 20032 2280 20052
rect 2280 20032 2282 20052
rect 3054 20052 3110 20088
rect 3054 20032 3056 20052
rect 3056 20032 3108 20052
rect 3108 20032 3110 20052
rect 4342 20052 4398 20088
rect 8798 20698 8854 20700
rect 8878 20698 8934 20700
rect 8958 20698 9014 20700
rect 9038 20698 9094 20700
rect 8798 20646 8844 20698
rect 8844 20646 8854 20698
rect 8878 20646 8908 20698
rect 8908 20646 8920 20698
rect 8920 20646 8934 20698
rect 8958 20646 8972 20698
rect 8972 20646 8984 20698
rect 8984 20646 9014 20698
rect 9038 20646 9048 20698
rect 9048 20646 9094 20698
rect 8798 20644 8854 20646
rect 8878 20644 8934 20646
rect 8958 20644 9014 20646
rect 9038 20644 9094 20646
rect 4342 20032 4344 20052
rect 4344 20032 4396 20052
rect 4396 20032 4398 20052
rect 5814 20052 5870 20088
rect 5814 20032 5816 20052
rect 5816 20032 5868 20052
rect 5868 20032 5870 20052
rect 6550 20052 6606 20088
rect 16640 20698 16696 20700
rect 16720 20698 16776 20700
rect 16800 20698 16856 20700
rect 16880 20698 16936 20700
rect 16640 20646 16686 20698
rect 16686 20646 16696 20698
rect 16720 20646 16750 20698
rect 16750 20646 16762 20698
rect 16762 20646 16776 20698
rect 16800 20646 16814 20698
rect 16814 20646 16826 20698
rect 16826 20646 16856 20698
rect 16880 20646 16890 20698
rect 16890 20646 16936 20698
rect 16640 20644 16696 20646
rect 16720 20644 16776 20646
rect 16800 20644 16856 20646
rect 16880 20644 16936 20646
rect 11978 20596 12034 20632
rect 11978 20576 11980 20596
rect 11980 20576 12032 20596
rect 12032 20576 12034 20596
rect 12714 20596 12770 20632
rect 12714 20576 12716 20596
rect 12716 20576 12768 20596
rect 12768 20576 12770 20596
rect 14830 20596 14886 20632
rect 17866 20712 17922 20768
rect 14830 20576 14832 20596
rect 14832 20576 14884 20596
rect 14884 20576 14886 20596
rect 11058 20440 11114 20496
rect 12719 20154 12775 20156
rect 12799 20154 12855 20156
rect 12879 20154 12935 20156
rect 12959 20154 13015 20156
rect 12719 20102 12765 20154
rect 12765 20102 12775 20154
rect 12799 20102 12829 20154
rect 12829 20102 12841 20154
rect 12841 20102 12855 20154
rect 12879 20102 12893 20154
rect 12893 20102 12905 20154
rect 12905 20102 12935 20154
rect 12959 20102 12969 20154
rect 12969 20102 13015 20154
rect 12719 20100 12775 20102
rect 12799 20100 12855 20102
rect 12879 20100 12935 20102
rect 12959 20100 13015 20102
rect 6550 20032 6552 20052
rect 6552 20032 6604 20052
rect 6604 20032 6606 20052
rect 13726 20052 13782 20088
rect 13726 20032 13728 20052
rect 13728 20032 13780 20052
rect 13780 20032 13782 20052
rect 11058 19916 11114 19952
rect 11058 19896 11060 19916
rect 11060 19896 11112 19916
rect 11112 19896 11114 19916
rect 2410 19508 2466 19544
rect 2410 19488 2412 19508
rect 2412 19488 2464 19508
rect 2464 19488 2466 19508
rect 3882 19508 3938 19544
rect 3882 19488 3884 19508
rect 3884 19488 3936 19508
rect 3936 19488 3938 19508
rect 8798 19610 8854 19612
rect 8878 19610 8934 19612
rect 8958 19610 9014 19612
rect 9038 19610 9094 19612
rect 8798 19558 8844 19610
rect 8844 19558 8854 19610
rect 8878 19558 8908 19610
rect 8908 19558 8920 19610
rect 8920 19558 8934 19610
rect 8958 19558 8972 19610
rect 8972 19558 8984 19610
rect 8984 19558 9014 19610
rect 9038 19558 9048 19610
rect 9048 19558 9094 19610
rect 8798 19556 8854 19558
rect 8878 19556 8934 19558
rect 8958 19556 9014 19558
rect 9038 19556 9094 19558
rect 10966 19508 11022 19544
rect 10966 19488 10968 19508
rect 10968 19488 11020 19508
rect 11020 19488 11022 19508
rect 11886 19508 11942 19544
rect 11886 19488 11888 19508
rect 11888 19488 11940 19508
rect 11940 19488 11942 19508
rect 4877 19066 4933 19068
rect 4957 19066 5013 19068
rect 5037 19066 5093 19068
rect 5117 19066 5173 19068
rect 4877 19014 4923 19066
rect 4923 19014 4933 19066
rect 4957 19014 4987 19066
rect 4987 19014 4999 19066
rect 4999 19014 5013 19066
rect 5037 19014 5051 19066
rect 5051 19014 5063 19066
rect 5063 19014 5093 19066
rect 5117 19014 5127 19066
rect 5127 19014 5173 19066
rect 4877 19012 4933 19014
rect 4957 19012 5013 19014
rect 5037 19012 5093 19014
rect 5117 19012 5173 19014
rect 11058 18964 11114 19000
rect 11058 18944 11060 18964
rect 11060 18944 11112 18964
rect 11112 18944 11114 18964
rect 12719 19066 12775 19068
rect 12799 19066 12855 19068
rect 12879 19066 12935 19068
rect 12959 19066 13015 19068
rect 12719 19014 12765 19066
rect 12765 19014 12775 19066
rect 12799 19014 12829 19066
rect 12829 19014 12841 19066
rect 12841 19014 12855 19066
rect 12879 19014 12893 19066
rect 12893 19014 12905 19066
rect 12905 19014 12935 19066
rect 12959 19014 12969 19066
rect 12969 19014 13015 19066
rect 12719 19012 12775 19014
rect 12799 19012 12855 19014
rect 12879 19012 12935 19014
rect 12959 19012 13015 19014
rect 8798 18522 8854 18524
rect 8878 18522 8934 18524
rect 8958 18522 9014 18524
rect 9038 18522 9094 18524
rect 8798 18470 8844 18522
rect 8844 18470 8854 18522
rect 8878 18470 8908 18522
rect 8908 18470 8920 18522
rect 8920 18470 8934 18522
rect 8958 18470 8972 18522
rect 8972 18470 8984 18522
rect 8984 18470 9014 18522
rect 9038 18470 9048 18522
rect 9048 18470 9094 18522
rect 8798 18468 8854 18470
rect 8878 18468 8934 18470
rect 8958 18468 9014 18470
rect 9038 18468 9094 18470
rect 13818 19236 13874 19272
rect 13818 19216 13820 19236
rect 13820 19216 13872 19236
rect 13872 19216 13874 19236
rect 16118 19508 16174 19544
rect 16118 19488 16120 19508
rect 16120 19488 16172 19508
rect 16172 19488 16174 19508
rect 16640 19610 16696 19612
rect 16720 19610 16776 19612
rect 16800 19610 16856 19612
rect 16880 19610 16936 19612
rect 16640 19558 16686 19610
rect 16686 19558 16696 19610
rect 16720 19558 16750 19610
rect 16750 19558 16762 19610
rect 16762 19558 16776 19610
rect 16800 19558 16814 19610
rect 16814 19558 16826 19610
rect 16826 19558 16856 19610
rect 16880 19558 16890 19610
rect 16890 19558 16936 19610
rect 16640 19556 16696 19558
rect 16720 19556 16776 19558
rect 16800 19556 16856 19558
rect 16880 19556 16936 19558
rect 18694 20596 18750 20632
rect 18694 20576 18696 20596
rect 18696 20576 18748 20596
rect 18748 20576 18750 20596
rect 17774 19372 17830 19408
rect 17774 19352 17776 19372
rect 17776 19352 17828 19372
rect 17828 19352 17830 19372
rect 16578 18964 16634 19000
rect 16578 18944 16580 18964
rect 16580 18944 16632 18964
rect 16632 18944 16634 18964
rect 22190 20984 22246 21040
rect 22926 20984 22982 21040
rect 20902 20848 20958 20904
rect 16640 18522 16696 18524
rect 16720 18522 16776 18524
rect 16800 18522 16856 18524
rect 16880 18522 16936 18524
rect 16640 18470 16686 18522
rect 16686 18470 16696 18522
rect 16720 18470 16750 18522
rect 16750 18470 16762 18522
rect 16762 18470 16776 18522
rect 16800 18470 16814 18522
rect 16814 18470 16826 18522
rect 16826 18470 16856 18522
rect 16880 18470 16890 18522
rect 16890 18470 16936 18522
rect 16640 18468 16696 18470
rect 16720 18468 16776 18470
rect 16800 18468 16856 18470
rect 16880 18468 16936 18470
rect 20561 20154 20617 20156
rect 20641 20154 20697 20156
rect 20721 20154 20777 20156
rect 20801 20154 20857 20156
rect 20561 20102 20607 20154
rect 20607 20102 20617 20154
rect 20641 20102 20671 20154
rect 20671 20102 20683 20154
rect 20683 20102 20697 20154
rect 20721 20102 20735 20154
rect 20735 20102 20747 20154
rect 20747 20102 20777 20154
rect 20801 20102 20811 20154
rect 20811 20102 20857 20154
rect 20561 20100 20617 20102
rect 20641 20100 20697 20102
rect 20721 20100 20777 20102
rect 20801 20100 20857 20102
rect 20561 19066 20617 19068
rect 20641 19066 20697 19068
rect 20721 19066 20777 19068
rect 20801 19066 20857 19068
rect 20561 19014 20607 19066
rect 20607 19014 20617 19066
rect 20641 19014 20671 19066
rect 20671 19014 20683 19066
rect 20683 19014 20697 19066
rect 20721 19014 20735 19066
rect 20735 19014 20747 19066
rect 20747 19014 20777 19066
rect 20801 19014 20811 19066
rect 20811 19014 20857 19066
rect 20561 19012 20617 19014
rect 20641 19012 20697 19014
rect 20721 19012 20777 19014
rect 20801 19012 20857 19014
rect 21454 20440 21510 20496
rect 24482 20698 24538 20700
rect 24562 20698 24618 20700
rect 24642 20698 24698 20700
rect 24722 20698 24778 20700
rect 24482 20646 24528 20698
rect 24528 20646 24538 20698
rect 24562 20646 24592 20698
rect 24592 20646 24604 20698
rect 24604 20646 24618 20698
rect 24642 20646 24656 20698
rect 24656 20646 24668 20698
rect 24668 20646 24698 20698
rect 24722 20646 24732 20698
rect 24732 20646 24778 20698
rect 24482 20644 24538 20646
rect 24562 20644 24618 20646
rect 24642 20644 24698 20646
rect 24722 20644 24778 20646
rect 24482 19610 24538 19612
rect 24562 19610 24618 19612
rect 24642 19610 24698 19612
rect 24722 19610 24778 19612
rect 24482 19558 24528 19610
rect 24528 19558 24538 19610
rect 24562 19558 24592 19610
rect 24592 19558 24604 19610
rect 24604 19558 24618 19610
rect 24642 19558 24656 19610
rect 24656 19558 24668 19610
rect 24668 19558 24698 19610
rect 24722 19558 24732 19610
rect 24732 19558 24778 19610
rect 24482 19556 24538 19558
rect 24562 19556 24618 19558
rect 24642 19556 24698 19558
rect 24722 19556 24778 19558
rect 24858 19216 24914 19272
rect 24482 18522 24538 18524
rect 24562 18522 24618 18524
rect 24642 18522 24698 18524
rect 24722 18522 24778 18524
rect 24482 18470 24528 18522
rect 24528 18470 24538 18522
rect 24562 18470 24592 18522
rect 24592 18470 24604 18522
rect 24604 18470 24618 18522
rect 24642 18470 24656 18522
rect 24656 18470 24668 18522
rect 24668 18470 24698 18522
rect 24722 18470 24732 18522
rect 24732 18470 24778 18522
rect 24482 18468 24538 18470
rect 24562 18468 24618 18470
rect 24642 18468 24698 18470
rect 24722 18468 24778 18470
rect 28403 20154 28459 20156
rect 28483 20154 28539 20156
rect 28563 20154 28619 20156
rect 28643 20154 28699 20156
rect 28403 20102 28449 20154
rect 28449 20102 28459 20154
rect 28483 20102 28513 20154
rect 28513 20102 28525 20154
rect 28525 20102 28539 20154
rect 28563 20102 28577 20154
rect 28577 20102 28589 20154
rect 28589 20102 28619 20154
rect 28643 20102 28653 20154
rect 28653 20102 28699 20154
rect 28403 20100 28459 20102
rect 28483 20100 28539 20102
rect 28563 20100 28619 20102
rect 28643 20100 28699 20102
rect 28403 19066 28459 19068
rect 28483 19066 28539 19068
rect 28563 19066 28619 19068
rect 28643 19066 28699 19068
rect 28403 19014 28449 19066
rect 28449 19014 28459 19066
rect 28483 19014 28513 19066
rect 28513 19014 28525 19066
rect 28525 19014 28539 19066
rect 28563 19014 28577 19066
rect 28577 19014 28589 19066
rect 28589 19014 28619 19066
rect 28643 19014 28653 19066
rect 28653 19014 28699 19066
rect 28403 19012 28459 19014
rect 28483 19012 28539 19014
rect 28563 19012 28619 19014
rect 28643 19012 28699 19014
rect 4877 17978 4933 17980
rect 4957 17978 5013 17980
rect 5037 17978 5093 17980
rect 5117 17978 5173 17980
rect 4877 17926 4923 17978
rect 4923 17926 4933 17978
rect 4957 17926 4987 17978
rect 4987 17926 4999 17978
rect 4999 17926 5013 17978
rect 5037 17926 5051 17978
rect 5051 17926 5063 17978
rect 5063 17926 5093 17978
rect 5117 17926 5127 17978
rect 5127 17926 5173 17978
rect 4877 17924 4933 17926
rect 4957 17924 5013 17926
rect 5037 17924 5093 17926
rect 5117 17924 5173 17926
rect 12719 17978 12775 17980
rect 12799 17978 12855 17980
rect 12879 17978 12935 17980
rect 12959 17978 13015 17980
rect 12719 17926 12765 17978
rect 12765 17926 12775 17978
rect 12799 17926 12829 17978
rect 12829 17926 12841 17978
rect 12841 17926 12855 17978
rect 12879 17926 12893 17978
rect 12893 17926 12905 17978
rect 12905 17926 12935 17978
rect 12959 17926 12969 17978
rect 12969 17926 13015 17978
rect 12719 17924 12775 17926
rect 12799 17924 12855 17926
rect 12879 17924 12935 17926
rect 12959 17924 13015 17926
rect 20561 17978 20617 17980
rect 20641 17978 20697 17980
rect 20721 17978 20777 17980
rect 20801 17978 20857 17980
rect 20561 17926 20607 17978
rect 20607 17926 20617 17978
rect 20641 17926 20671 17978
rect 20671 17926 20683 17978
rect 20683 17926 20697 17978
rect 20721 17926 20735 17978
rect 20735 17926 20747 17978
rect 20747 17926 20777 17978
rect 20801 17926 20811 17978
rect 20811 17926 20857 17978
rect 20561 17924 20617 17926
rect 20641 17924 20697 17926
rect 20721 17924 20777 17926
rect 20801 17924 20857 17926
rect 28403 17978 28459 17980
rect 28483 17978 28539 17980
rect 28563 17978 28619 17980
rect 28643 17978 28699 17980
rect 28403 17926 28449 17978
rect 28449 17926 28459 17978
rect 28483 17926 28513 17978
rect 28513 17926 28525 17978
rect 28525 17926 28539 17978
rect 28563 17926 28577 17978
rect 28577 17926 28589 17978
rect 28589 17926 28619 17978
rect 28643 17926 28653 17978
rect 28653 17926 28699 17978
rect 28403 17924 28459 17926
rect 28483 17924 28539 17926
rect 28563 17924 28619 17926
rect 28643 17924 28699 17926
rect 30286 17856 30342 17912
rect 31758 20712 31814 20768
rect 31298 19624 31354 19680
rect 32324 20698 32380 20700
rect 32404 20698 32460 20700
rect 32484 20698 32540 20700
rect 32564 20698 32620 20700
rect 32324 20646 32370 20698
rect 32370 20646 32380 20698
rect 32404 20646 32434 20698
rect 32434 20646 32446 20698
rect 32446 20646 32460 20698
rect 32484 20646 32498 20698
rect 32498 20646 32510 20698
rect 32510 20646 32540 20698
rect 32564 20646 32574 20698
rect 32574 20646 32620 20698
rect 32324 20644 32380 20646
rect 32404 20644 32460 20646
rect 32484 20644 32540 20646
rect 32564 20644 32620 20646
rect 32324 19610 32380 19612
rect 32404 19610 32460 19612
rect 32484 19610 32540 19612
rect 32564 19610 32620 19612
rect 32324 19558 32370 19610
rect 32370 19558 32380 19610
rect 32404 19558 32434 19610
rect 32434 19558 32446 19610
rect 32446 19558 32460 19610
rect 32484 19558 32498 19610
rect 32498 19558 32510 19610
rect 32510 19558 32540 19610
rect 32564 19558 32574 19610
rect 32574 19558 32620 19610
rect 32324 19556 32380 19558
rect 32404 19556 32460 19558
rect 32484 19556 32540 19558
rect 32564 19556 32620 19558
rect 32324 18522 32380 18524
rect 32404 18522 32460 18524
rect 32484 18522 32540 18524
rect 32564 18522 32620 18524
rect 32324 18470 32370 18522
rect 32370 18470 32380 18522
rect 32404 18470 32434 18522
rect 32434 18470 32446 18522
rect 32446 18470 32460 18522
rect 32484 18470 32498 18522
rect 32498 18470 32510 18522
rect 32510 18470 32540 18522
rect 32564 18470 32574 18522
rect 32574 18470 32620 18522
rect 32324 18468 32380 18470
rect 32404 18468 32460 18470
rect 32484 18468 32540 18470
rect 32564 18468 32620 18470
rect 8798 17434 8854 17436
rect 8878 17434 8934 17436
rect 8958 17434 9014 17436
rect 9038 17434 9094 17436
rect 8798 17382 8844 17434
rect 8844 17382 8854 17434
rect 8878 17382 8908 17434
rect 8908 17382 8920 17434
rect 8920 17382 8934 17434
rect 8958 17382 8972 17434
rect 8972 17382 8984 17434
rect 8984 17382 9014 17434
rect 9038 17382 9048 17434
rect 9048 17382 9094 17434
rect 8798 17380 8854 17382
rect 8878 17380 8934 17382
rect 8958 17380 9014 17382
rect 9038 17380 9094 17382
rect 16640 17434 16696 17436
rect 16720 17434 16776 17436
rect 16800 17434 16856 17436
rect 16880 17434 16936 17436
rect 16640 17382 16686 17434
rect 16686 17382 16696 17434
rect 16720 17382 16750 17434
rect 16750 17382 16762 17434
rect 16762 17382 16776 17434
rect 16800 17382 16814 17434
rect 16814 17382 16826 17434
rect 16826 17382 16856 17434
rect 16880 17382 16890 17434
rect 16890 17382 16936 17434
rect 16640 17380 16696 17382
rect 16720 17380 16776 17382
rect 16800 17380 16856 17382
rect 16880 17380 16936 17382
rect 24482 17434 24538 17436
rect 24562 17434 24618 17436
rect 24642 17434 24698 17436
rect 24722 17434 24778 17436
rect 24482 17382 24528 17434
rect 24528 17382 24538 17434
rect 24562 17382 24592 17434
rect 24592 17382 24604 17434
rect 24604 17382 24618 17434
rect 24642 17382 24656 17434
rect 24656 17382 24668 17434
rect 24668 17382 24698 17434
rect 24722 17382 24732 17434
rect 24732 17382 24778 17434
rect 24482 17380 24538 17382
rect 24562 17380 24618 17382
rect 24642 17380 24698 17382
rect 24722 17380 24778 17382
rect 32324 17434 32380 17436
rect 32404 17434 32460 17436
rect 32484 17434 32540 17436
rect 32564 17434 32620 17436
rect 32324 17382 32370 17434
rect 32370 17382 32380 17434
rect 32404 17382 32434 17434
rect 32434 17382 32446 17434
rect 32446 17382 32460 17434
rect 32484 17382 32498 17434
rect 32498 17382 32510 17434
rect 32510 17382 32540 17434
rect 32564 17382 32574 17434
rect 32574 17382 32620 17434
rect 32324 17380 32380 17382
rect 32404 17380 32460 17382
rect 32484 17380 32540 17382
rect 32564 17380 32620 17382
rect 4877 16890 4933 16892
rect 4957 16890 5013 16892
rect 5037 16890 5093 16892
rect 5117 16890 5173 16892
rect 4877 16838 4923 16890
rect 4923 16838 4933 16890
rect 4957 16838 4987 16890
rect 4987 16838 4999 16890
rect 4999 16838 5013 16890
rect 5037 16838 5051 16890
rect 5051 16838 5063 16890
rect 5063 16838 5093 16890
rect 5117 16838 5127 16890
rect 5127 16838 5173 16890
rect 4877 16836 4933 16838
rect 4957 16836 5013 16838
rect 5037 16836 5093 16838
rect 5117 16836 5173 16838
rect 12719 16890 12775 16892
rect 12799 16890 12855 16892
rect 12879 16890 12935 16892
rect 12959 16890 13015 16892
rect 12719 16838 12765 16890
rect 12765 16838 12775 16890
rect 12799 16838 12829 16890
rect 12829 16838 12841 16890
rect 12841 16838 12855 16890
rect 12879 16838 12893 16890
rect 12893 16838 12905 16890
rect 12905 16838 12935 16890
rect 12959 16838 12969 16890
rect 12969 16838 13015 16890
rect 12719 16836 12775 16838
rect 12799 16836 12855 16838
rect 12879 16836 12935 16838
rect 12959 16836 13015 16838
rect 20561 16890 20617 16892
rect 20641 16890 20697 16892
rect 20721 16890 20777 16892
rect 20801 16890 20857 16892
rect 20561 16838 20607 16890
rect 20607 16838 20617 16890
rect 20641 16838 20671 16890
rect 20671 16838 20683 16890
rect 20683 16838 20697 16890
rect 20721 16838 20735 16890
rect 20735 16838 20747 16890
rect 20747 16838 20777 16890
rect 20801 16838 20811 16890
rect 20811 16838 20857 16890
rect 20561 16836 20617 16838
rect 20641 16836 20697 16838
rect 20721 16836 20777 16838
rect 20801 16836 20857 16838
rect 28403 16890 28459 16892
rect 28483 16890 28539 16892
rect 28563 16890 28619 16892
rect 28643 16890 28699 16892
rect 28403 16838 28449 16890
rect 28449 16838 28459 16890
rect 28483 16838 28513 16890
rect 28513 16838 28525 16890
rect 28525 16838 28539 16890
rect 28563 16838 28577 16890
rect 28577 16838 28589 16890
rect 28589 16838 28619 16890
rect 28643 16838 28653 16890
rect 28653 16838 28699 16890
rect 28403 16836 28459 16838
rect 28483 16836 28539 16838
rect 28563 16836 28619 16838
rect 28643 16836 28699 16838
rect 8798 16346 8854 16348
rect 8878 16346 8934 16348
rect 8958 16346 9014 16348
rect 9038 16346 9094 16348
rect 8798 16294 8844 16346
rect 8844 16294 8854 16346
rect 8878 16294 8908 16346
rect 8908 16294 8920 16346
rect 8920 16294 8934 16346
rect 8958 16294 8972 16346
rect 8972 16294 8984 16346
rect 8984 16294 9014 16346
rect 9038 16294 9048 16346
rect 9048 16294 9094 16346
rect 8798 16292 8854 16294
rect 8878 16292 8934 16294
rect 8958 16292 9014 16294
rect 9038 16292 9094 16294
rect 16640 16346 16696 16348
rect 16720 16346 16776 16348
rect 16800 16346 16856 16348
rect 16880 16346 16936 16348
rect 16640 16294 16686 16346
rect 16686 16294 16696 16346
rect 16720 16294 16750 16346
rect 16750 16294 16762 16346
rect 16762 16294 16776 16346
rect 16800 16294 16814 16346
rect 16814 16294 16826 16346
rect 16826 16294 16856 16346
rect 16880 16294 16890 16346
rect 16890 16294 16936 16346
rect 16640 16292 16696 16294
rect 16720 16292 16776 16294
rect 16800 16292 16856 16294
rect 16880 16292 16936 16294
rect 24482 16346 24538 16348
rect 24562 16346 24618 16348
rect 24642 16346 24698 16348
rect 24722 16346 24778 16348
rect 24482 16294 24528 16346
rect 24528 16294 24538 16346
rect 24562 16294 24592 16346
rect 24592 16294 24604 16346
rect 24604 16294 24618 16346
rect 24642 16294 24656 16346
rect 24656 16294 24668 16346
rect 24668 16294 24698 16346
rect 24722 16294 24732 16346
rect 24732 16294 24778 16346
rect 24482 16292 24538 16294
rect 24562 16292 24618 16294
rect 24642 16292 24698 16294
rect 24722 16292 24778 16294
rect 32324 16346 32380 16348
rect 32404 16346 32460 16348
rect 32484 16346 32540 16348
rect 32564 16346 32620 16348
rect 32324 16294 32370 16346
rect 32370 16294 32380 16346
rect 32404 16294 32434 16346
rect 32434 16294 32446 16346
rect 32446 16294 32460 16346
rect 32484 16294 32498 16346
rect 32498 16294 32510 16346
rect 32510 16294 32540 16346
rect 32564 16294 32574 16346
rect 32574 16294 32620 16346
rect 32324 16292 32380 16294
rect 32404 16292 32460 16294
rect 32484 16292 32540 16294
rect 32564 16292 32620 16294
rect 4877 15802 4933 15804
rect 4957 15802 5013 15804
rect 5037 15802 5093 15804
rect 5117 15802 5173 15804
rect 4877 15750 4923 15802
rect 4923 15750 4933 15802
rect 4957 15750 4987 15802
rect 4987 15750 4999 15802
rect 4999 15750 5013 15802
rect 5037 15750 5051 15802
rect 5051 15750 5063 15802
rect 5063 15750 5093 15802
rect 5117 15750 5127 15802
rect 5127 15750 5173 15802
rect 4877 15748 4933 15750
rect 4957 15748 5013 15750
rect 5037 15748 5093 15750
rect 5117 15748 5173 15750
rect 12719 15802 12775 15804
rect 12799 15802 12855 15804
rect 12879 15802 12935 15804
rect 12959 15802 13015 15804
rect 12719 15750 12765 15802
rect 12765 15750 12775 15802
rect 12799 15750 12829 15802
rect 12829 15750 12841 15802
rect 12841 15750 12855 15802
rect 12879 15750 12893 15802
rect 12893 15750 12905 15802
rect 12905 15750 12935 15802
rect 12959 15750 12969 15802
rect 12969 15750 13015 15802
rect 12719 15748 12775 15750
rect 12799 15748 12855 15750
rect 12879 15748 12935 15750
rect 12959 15748 13015 15750
rect 20561 15802 20617 15804
rect 20641 15802 20697 15804
rect 20721 15802 20777 15804
rect 20801 15802 20857 15804
rect 20561 15750 20607 15802
rect 20607 15750 20617 15802
rect 20641 15750 20671 15802
rect 20671 15750 20683 15802
rect 20683 15750 20697 15802
rect 20721 15750 20735 15802
rect 20735 15750 20747 15802
rect 20747 15750 20777 15802
rect 20801 15750 20811 15802
rect 20811 15750 20857 15802
rect 20561 15748 20617 15750
rect 20641 15748 20697 15750
rect 20721 15748 20777 15750
rect 20801 15748 20857 15750
rect 28403 15802 28459 15804
rect 28483 15802 28539 15804
rect 28563 15802 28619 15804
rect 28643 15802 28699 15804
rect 28403 15750 28449 15802
rect 28449 15750 28459 15802
rect 28483 15750 28513 15802
rect 28513 15750 28525 15802
rect 28525 15750 28539 15802
rect 28563 15750 28577 15802
rect 28577 15750 28589 15802
rect 28589 15750 28619 15802
rect 28643 15750 28653 15802
rect 28653 15750 28699 15802
rect 28403 15748 28459 15750
rect 28483 15748 28539 15750
rect 28563 15748 28619 15750
rect 28643 15748 28699 15750
rect 8798 15258 8854 15260
rect 8878 15258 8934 15260
rect 8958 15258 9014 15260
rect 9038 15258 9094 15260
rect 8798 15206 8844 15258
rect 8844 15206 8854 15258
rect 8878 15206 8908 15258
rect 8908 15206 8920 15258
rect 8920 15206 8934 15258
rect 8958 15206 8972 15258
rect 8972 15206 8984 15258
rect 8984 15206 9014 15258
rect 9038 15206 9048 15258
rect 9048 15206 9094 15258
rect 8798 15204 8854 15206
rect 8878 15204 8934 15206
rect 8958 15204 9014 15206
rect 9038 15204 9094 15206
rect 16640 15258 16696 15260
rect 16720 15258 16776 15260
rect 16800 15258 16856 15260
rect 16880 15258 16936 15260
rect 16640 15206 16686 15258
rect 16686 15206 16696 15258
rect 16720 15206 16750 15258
rect 16750 15206 16762 15258
rect 16762 15206 16776 15258
rect 16800 15206 16814 15258
rect 16814 15206 16826 15258
rect 16826 15206 16856 15258
rect 16880 15206 16890 15258
rect 16890 15206 16936 15258
rect 16640 15204 16696 15206
rect 16720 15204 16776 15206
rect 16800 15204 16856 15206
rect 16880 15204 16936 15206
rect 24482 15258 24538 15260
rect 24562 15258 24618 15260
rect 24642 15258 24698 15260
rect 24722 15258 24778 15260
rect 24482 15206 24528 15258
rect 24528 15206 24538 15258
rect 24562 15206 24592 15258
rect 24592 15206 24604 15258
rect 24604 15206 24618 15258
rect 24642 15206 24656 15258
rect 24656 15206 24668 15258
rect 24668 15206 24698 15258
rect 24722 15206 24732 15258
rect 24732 15206 24778 15258
rect 24482 15204 24538 15206
rect 24562 15204 24618 15206
rect 24642 15204 24698 15206
rect 24722 15204 24778 15206
rect 32324 15258 32380 15260
rect 32404 15258 32460 15260
rect 32484 15258 32540 15260
rect 32564 15258 32620 15260
rect 32324 15206 32370 15258
rect 32370 15206 32380 15258
rect 32404 15206 32434 15258
rect 32434 15206 32446 15258
rect 32446 15206 32460 15258
rect 32484 15206 32498 15258
rect 32498 15206 32510 15258
rect 32510 15206 32540 15258
rect 32564 15206 32574 15258
rect 32574 15206 32620 15258
rect 32324 15204 32380 15206
rect 32404 15204 32460 15206
rect 32484 15204 32540 15206
rect 32564 15204 32620 15206
rect 4877 14714 4933 14716
rect 4957 14714 5013 14716
rect 5037 14714 5093 14716
rect 5117 14714 5173 14716
rect 4877 14662 4923 14714
rect 4923 14662 4933 14714
rect 4957 14662 4987 14714
rect 4987 14662 4999 14714
rect 4999 14662 5013 14714
rect 5037 14662 5051 14714
rect 5051 14662 5063 14714
rect 5063 14662 5093 14714
rect 5117 14662 5127 14714
rect 5127 14662 5173 14714
rect 4877 14660 4933 14662
rect 4957 14660 5013 14662
rect 5037 14660 5093 14662
rect 5117 14660 5173 14662
rect 12719 14714 12775 14716
rect 12799 14714 12855 14716
rect 12879 14714 12935 14716
rect 12959 14714 13015 14716
rect 12719 14662 12765 14714
rect 12765 14662 12775 14714
rect 12799 14662 12829 14714
rect 12829 14662 12841 14714
rect 12841 14662 12855 14714
rect 12879 14662 12893 14714
rect 12893 14662 12905 14714
rect 12905 14662 12935 14714
rect 12959 14662 12969 14714
rect 12969 14662 13015 14714
rect 12719 14660 12775 14662
rect 12799 14660 12855 14662
rect 12879 14660 12935 14662
rect 12959 14660 13015 14662
rect 20561 14714 20617 14716
rect 20641 14714 20697 14716
rect 20721 14714 20777 14716
rect 20801 14714 20857 14716
rect 20561 14662 20607 14714
rect 20607 14662 20617 14714
rect 20641 14662 20671 14714
rect 20671 14662 20683 14714
rect 20683 14662 20697 14714
rect 20721 14662 20735 14714
rect 20735 14662 20747 14714
rect 20747 14662 20777 14714
rect 20801 14662 20811 14714
rect 20811 14662 20857 14714
rect 20561 14660 20617 14662
rect 20641 14660 20697 14662
rect 20721 14660 20777 14662
rect 20801 14660 20857 14662
rect 28403 14714 28459 14716
rect 28483 14714 28539 14716
rect 28563 14714 28619 14716
rect 28643 14714 28699 14716
rect 28403 14662 28449 14714
rect 28449 14662 28459 14714
rect 28483 14662 28513 14714
rect 28513 14662 28525 14714
rect 28525 14662 28539 14714
rect 28563 14662 28577 14714
rect 28577 14662 28589 14714
rect 28589 14662 28619 14714
rect 28643 14662 28653 14714
rect 28653 14662 28699 14714
rect 28403 14660 28459 14662
rect 28483 14660 28539 14662
rect 28563 14660 28619 14662
rect 28643 14660 28699 14662
rect 8798 14170 8854 14172
rect 8878 14170 8934 14172
rect 8958 14170 9014 14172
rect 9038 14170 9094 14172
rect 8798 14118 8844 14170
rect 8844 14118 8854 14170
rect 8878 14118 8908 14170
rect 8908 14118 8920 14170
rect 8920 14118 8934 14170
rect 8958 14118 8972 14170
rect 8972 14118 8984 14170
rect 8984 14118 9014 14170
rect 9038 14118 9048 14170
rect 9048 14118 9094 14170
rect 8798 14116 8854 14118
rect 8878 14116 8934 14118
rect 8958 14116 9014 14118
rect 9038 14116 9094 14118
rect 16640 14170 16696 14172
rect 16720 14170 16776 14172
rect 16800 14170 16856 14172
rect 16880 14170 16936 14172
rect 16640 14118 16686 14170
rect 16686 14118 16696 14170
rect 16720 14118 16750 14170
rect 16750 14118 16762 14170
rect 16762 14118 16776 14170
rect 16800 14118 16814 14170
rect 16814 14118 16826 14170
rect 16826 14118 16856 14170
rect 16880 14118 16890 14170
rect 16890 14118 16936 14170
rect 16640 14116 16696 14118
rect 16720 14116 16776 14118
rect 16800 14116 16856 14118
rect 16880 14116 16936 14118
rect 24482 14170 24538 14172
rect 24562 14170 24618 14172
rect 24642 14170 24698 14172
rect 24722 14170 24778 14172
rect 24482 14118 24528 14170
rect 24528 14118 24538 14170
rect 24562 14118 24592 14170
rect 24592 14118 24604 14170
rect 24604 14118 24618 14170
rect 24642 14118 24656 14170
rect 24656 14118 24668 14170
rect 24668 14118 24698 14170
rect 24722 14118 24732 14170
rect 24732 14118 24778 14170
rect 24482 14116 24538 14118
rect 24562 14116 24618 14118
rect 24642 14116 24698 14118
rect 24722 14116 24778 14118
rect 32324 14170 32380 14172
rect 32404 14170 32460 14172
rect 32484 14170 32540 14172
rect 32564 14170 32620 14172
rect 32324 14118 32370 14170
rect 32370 14118 32380 14170
rect 32404 14118 32434 14170
rect 32434 14118 32446 14170
rect 32446 14118 32460 14170
rect 32484 14118 32498 14170
rect 32498 14118 32510 14170
rect 32510 14118 32540 14170
rect 32564 14118 32574 14170
rect 32574 14118 32620 14170
rect 32324 14116 32380 14118
rect 32404 14116 32460 14118
rect 32484 14116 32540 14118
rect 32564 14116 32620 14118
rect 4877 13626 4933 13628
rect 4957 13626 5013 13628
rect 5037 13626 5093 13628
rect 5117 13626 5173 13628
rect 4877 13574 4923 13626
rect 4923 13574 4933 13626
rect 4957 13574 4987 13626
rect 4987 13574 4999 13626
rect 4999 13574 5013 13626
rect 5037 13574 5051 13626
rect 5051 13574 5063 13626
rect 5063 13574 5093 13626
rect 5117 13574 5127 13626
rect 5127 13574 5173 13626
rect 4877 13572 4933 13574
rect 4957 13572 5013 13574
rect 5037 13572 5093 13574
rect 5117 13572 5173 13574
rect 12719 13626 12775 13628
rect 12799 13626 12855 13628
rect 12879 13626 12935 13628
rect 12959 13626 13015 13628
rect 12719 13574 12765 13626
rect 12765 13574 12775 13626
rect 12799 13574 12829 13626
rect 12829 13574 12841 13626
rect 12841 13574 12855 13626
rect 12879 13574 12893 13626
rect 12893 13574 12905 13626
rect 12905 13574 12935 13626
rect 12959 13574 12969 13626
rect 12969 13574 13015 13626
rect 12719 13572 12775 13574
rect 12799 13572 12855 13574
rect 12879 13572 12935 13574
rect 12959 13572 13015 13574
rect 20561 13626 20617 13628
rect 20641 13626 20697 13628
rect 20721 13626 20777 13628
rect 20801 13626 20857 13628
rect 20561 13574 20607 13626
rect 20607 13574 20617 13626
rect 20641 13574 20671 13626
rect 20671 13574 20683 13626
rect 20683 13574 20697 13626
rect 20721 13574 20735 13626
rect 20735 13574 20747 13626
rect 20747 13574 20777 13626
rect 20801 13574 20811 13626
rect 20811 13574 20857 13626
rect 20561 13572 20617 13574
rect 20641 13572 20697 13574
rect 20721 13572 20777 13574
rect 20801 13572 20857 13574
rect 28403 13626 28459 13628
rect 28483 13626 28539 13628
rect 28563 13626 28619 13628
rect 28643 13626 28699 13628
rect 28403 13574 28449 13626
rect 28449 13574 28459 13626
rect 28483 13574 28513 13626
rect 28513 13574 28525 13626
rect 28525 13574 28539 13626
rect 28563 13574 28577 13626
rect 28577 13574 28589 13626
rect 28589 13574 28619 13626
rect 28643 13574 28653 13626
rect 28653 13574 28699 13626
rect 28403 13572 28459 13574
rect 28483 13572 28539 13574
rect 28563 13572 28619 13574
rect 28643 13572 28699 13574
rect 8798 13082 8854 13084
rect 8878 13082 8934 13084
rect 8958 13082 9014 13084
rect 9038 13082 9094 13084
rect 8798 13030 8844 13082
rect 8844 13030 8854 13082
rect 8878 13030 8908 13082
rect 8908 13030 8920 13082
rect 8920 13030 8934 13082
rect 8958 13030 8972 13082
rect 8972 13030 8984 13082
rect 8984 13030 9014 13082
rect 9038 13030 9048 13082
rect 9048 13030 9094 13082
rect 8798 13028 8854 13030
rect 8878 13028 8934 13030
rect 8958 13028 9014 13030
rect 9038 13028 9094 13030
rect 16640 13082 16696 13084
rect 16720 13082 16776 13084
rect 16800 13082 16856 13084
rect 16880 13082 16936 13084
rect 16640 13030 16686 13082
rect 16686 13030 16696 13082
rect 16720 13030 16750 13082
rect 16750 13030 16762 13082
rect 16762 13030 16776 13082
rect 16800 13030 16814 13082
rect 16814 13030 16826 13082
rect 16826 13030 16856 13082
rect 16880 13030 16890 13082
rect 16890 13030 16936 13082
rect 16640 13028 16696 13030
rect 16720 13028 16776 13030
rect 16800 13028 16856 13030
rect 16880 13028 16936 13030
rect 24482 13082 24538 13084
rect 24562 13082 24618 13084
rect 24642 13082 24698 13084
rect 24722 13082 24778 13084
rect 24482 13030 24528 13082
rect 24528 13030 24538 13082
rect 24562 13030 24592 13082
rect 24592 13030 24604 13082
rect 24604 13030 24618 13082
rect 24642 13030 24656 13082
rect 24656 13030 24668 13082
rect 24668 13030 24698 13082
rect 24722 13030 24732 13082
rect 24732 13030 24778 13082
rect 24482 13028 24538 13030
rect 24562 13028 24618 13030
rect 24642 13028 24698 13030
rect 24722 13028 24778 13030
rect 32324 13082 32380 13084
rect 32404 13082 32460 13084
rect 32484 13082 32540 13084
rect 32564 13082 32620 13084
rect 32324 13030 32370 13082
rect 32370 13030 32380 13082
rect 32404 13030 32434 13082
rect 32434 13030 32446 13082
rect 32446 13030 32460 13082
rect 32484 13030 32498 13082
rect 32498 13030 32510 13082
rect 32510 13030 32540 13082
rect 32564 13030 32574 13082
rect 32574 13030 32620 13082
rect 32324 13028 32380 13030
rect 32404 13028 32460 13030
rect 32484 13028 32540 13030
rect 32564 13028 32620 13030
rect 4877 12538 4933 12540
rect 4957 12538 5013 12540
rect 5037 12538 5093 12540
rect 5117 12538 5173 12540
rect 4877 12486 4923 12538
rect 4923 12486 4933 12538
rect 4957 12486 4987 12538
rect 4987 12486 4999 12538
rect 4999 12486 5013 12538
rect 5037 12486 5051 12538
rect 5051 12486 5063 12538
rect 5063 12486 5093 12538
rect 5117 12486 5127 12538
rect 5127 12486 5173 12538
rect 4877 12484 4933 12486
rect 4957 12484 5013 12486
rect 5037 12484 5093 12486
rect 5117 12484 5173 12486
rect 12719 12538 12775 12540
rect 12799 12538 12855 12540
rect 12879 12538 12935 12540
rect 12959 12538 13015 12540
rect 12719 12486 12765 12538
rect 12765 12486 12775 12538
rect 12799 12486 12829 12538
rect 12829 12486 12841 12538
rect 12841 12486 12855 12538
rect 12879 12486 12893 12538
rect 12893 12486 12905 12538
rect 12905 12486 12935 12538
rect 12959 12486 12969 12538
rect 12969 12486 13015 12538
rect 12719 12484 12775 12486
rect 12799 12484 12855 12486
rect 12879 12484 12935 12486
rect 12959 12484 13015 12486
rect 20561 12538 20617 12540
rect 20641 12538 20697 12540
rect 20721 12538 20777 12540
rect 20801 12538 20857 12540
rect 20561 12486 20607 12538
rect 20607 12486 20617 12538
rect 20641 12486 20671 12538
rect 20671 12486 20683 12538
rect 20683 12486 20697 12538
rect 20721 12486 20735 12538
rect 20735 12486 20747 12538
rect 20747 12486 20777 12538
rect 20801 12486 20811 12538
rect 20811 12486 20857 12538
rect 20561 12484 20617 12486
rect 20641 12484 20697 12486
rect 20721 12484 20777 12486
rect 20801 12484 20857 12486
rect 28403 12538 28459 12540
rect 28483 12538 28539 12540
rect 28563 12538 28619 12540
rect 28643 12538 28699 12540
rect 28403 12486 28449 12538
rect 28449 12486 28459 12538
rect 28483 12486 28513 12538
rect 28513 12486 28525 12538
rect 28525 12486 28539 12538
rect 28563 12486 28577 12538
rect 28577 12486 28589 12538
rect 28589 12486 28619 12538
rect 28643 12486 28653 12538
rect 28653 12486 28699 12538
rect 28403 12484 28459 12486
rect 28483 12484 28539 12486
rect 28563 12484 28619 12486
rect 28643 12484 28699 12486
rect 8798 11994 8854 11996
rect 8878 11994 8934 11996
rect 8958 11994 9014 11996
rect 9038 11994 9094 11996
rect 8798 11942 8844 11994
rect 8844 11942 8854 11994
rect 8878 11942 8908 11994
rect 8908 11942 8920 11994
rect 8920 11942 8934 11994
rect 8958 11942 8972 11994
rect 8972 11942 8984 11994
rect 8984 11942 9014 11994
rect 9038 11942 9048 11994
rect 9048 11942 9094 11994
rect 8798 11940 8854 11942
rect 8878 11940 8934 11942
rect 8958 11940 9014 11942
rect 9038 11940 9094 11942
rect 16640 11994 16696 11996
rect 16720 11994 16776 11996
rect 16800 11994 16856 11996
rect 16880 11994 16936 11996
rect 16640 11942 16686 11994
rect 16686 11942 16696 11994
rect 16720 11942 16750 11994
rect 16750 11942 16762 11994
rect 16762 11942 16776 11994
rect 16800 11942 16814 11994
rect 16814 11942 16826 11994
rect 16826 11942 16856 11994
rect 16880 11942 16890 11994
rect 16890 11942 16936 11994
rect 16640 11940 16696 11942
rect 16720 11940 16776 11942
rect 16800 11940 16856 11942
rect 16880 11940 16936 11942
rect 24482 11994 24538 11996
rect 24562 11994 24618 11996
rect 24642 11994 24698 11996
rect 24722 11994 24778 11996
rect 24482 11942 24528 11994
rect 24528 11942 24538 11994
rect 24562 11942 24592 11994
rect 24592 11942 24604 11994
rect 24604 11942 24618 11994
rect 24642 11942 24656 11994
rect 24656 11942 24668 11994
rect 24668 11942 24698 11994
rect 24722 11942 24732 11994
rect 24732 11942 24778 11994
rect 24482 11940 24538 11942
rect 24562 11940 24618 11942
rect 24642 11940 24698 11942
rect 24722 11940 24778 11942
rect 32324 11994 32380 11996
rect 32404 11994 32460 11996
rect 32484 11994 32540 11996
rect 32564 11994 32620 11996
rect 32324 11942 32370 11994
rect 32370 11942 32380 11994
rect 32404 11942 32434 11994
rect 32434 11942 32446 11994
rect 32446 11942 32460 11994
rect 32484 11942 32498 11994
rect 32498 11942 32510 11994
rect 32510 11942 32540 11994
rect 32564 11942 32574 11994
rect 32574 11942 32620 11994
rect 32324 11940 32380 11942
rect 32404 11940 32460 11942
rect 32484 11940 32540 11942
rect 32564 11940 32620 11942
rect 4877 11450 4933 11452
rect 4957 11450 5013 11452
rect 5037 11450 5093 11452
rect 5117 11450 5173 11452
rect 4877 11398 4923 11450
rect 4923 11398 4933 11450
rect 4957 11398 4987 11450
rect 4987 11398 4999 11450
rect 4999 11398 5013 11450
rect 5037 11398 5051 11450
rect 5051 11398 5063 11450
rect 5063 11398 5093 11450
rect 5117 11398 5127 11450
rect 5127 11398 5173 11450
rect 4877 11396 4933 11398
rect 4957 11396 5013 11398
rect 5037 11396 5093 11398
rect 5117 11396 5173 11398
rect 12719 11450 12775 11452
rect 12799 11450 12855 11452
rect 12879 11450 12935 11452
rect 12959 11450 13015 11452
rect 12719 11398 12765 11450
rect 12765 11398 12775 11450
rect 12799 11398 12829 11450
rect 12829 11398 12841 11450
rect 12841 11398 12855 11450
rect 12879 11398 12893 11450
rect 12893 11398 12905 11450
rect 12905 11398 12935 11450
rect 12959 11398 12969 11450
rect 12969 11398 13015 11450
rect 12719 11396 12775 11398
rect 12799 11396 12855 11398
rect 12879 11396 12935 11398
rect 12959 11396 13015 11398
rect 20561 11450 20617 11452
rect 20641 11450 20697 11452
rect 20721 11450 20777 11452
rect 20801 11450 20857 11452
rect 20561 11398 20607 11450
rect 20607 11398 20617 11450
rect 20641 11398 20671 11450
rect 20671 11398 20683 11450
rect 20683 11398 20697 11450
rect 20721 11398 20735 11450
rect 20735 11398 20747 11450
rect 20747 11398 20777 11450
rect 20801 11398 20811 11450
rect 20811 11398 20857 11450
rect 20561 11396 20617 11398
rect 20641 11396 20697 11398
rect 20721 11396 20777 11398
rect 20801 11396 20857 11398
rect 28403 11450 28459 11452
rect 28483 11450 28539 11452
rect 28563 11450 28619 11452
rect 28643 11450 28699 11452
rect 28403 11398 28449 11450
rect 28449 11398 28459 11450
rect 28483 11398 28513 11450
rect 28513 11398 28525 11450
rect 28525 11398 28539 11450
rect 28563 11398 28577 11450
rect 28577 11398 28589 11450
rect 28589 11398 28619 11450
rect 28643 11398 28653 11450
rect 28653 11398 28699 11450
rect 28403 11396 28459 11398
rect 28483 11396 28539 11398
rect 28563 11396 28619 11398
rect 28643 11396 28699 11398
rect 8798 10906 8854 10908
rect 8878 10906 8934 10908
rect 8958 10906 9014 10908
rect 9038 10906 9094 10908
rect 8798 10854 8844 10906
rect 8844 10854 8854 10906
rect 8878 10854 8908 10906
rect 8908 10854 8920 10906
rect 8920 10854 8934 10906
rect 8958 10854 8972 10906
rect 8972 10854 8984 10906
rect 8984 10854 9014 10906
rect 9038 10854 9048 10906
rect 9048 10854 9094 10906
rect 8798 10852 8854 10854
rect 8878 10852 8934 10854
rect 8958 10852 9014 10854
rect 9038 10852 9094 10854
rect 16640 10906 16696 10908
rect 16720 10906 16776 10908
rect 16800 10906 16856 10908
rect 16880 10906 16936 10908
rect 16640 10854 16686 10906
rect 16686 10854 16696 10906
rect 16720 10854 16750 10906
rect 16750 10854 16762 10906
rect 16762 10854 16776 10906
rect 16800 10854 16814 10906
rect 16814 10854 16826 10906
rect 16826 10854 16856 10906
rect 16880 10854 16890 10906
rect 16890 10854 16936 10906
rect 16640 10852 16696 10854
rect 16720 10852 16776 10854
rect 16800 10852 16856 10854
rect 16880 10852 16936 10854
rect 24482 10906 24538 10908
rect 24562 10906 24618 10908
rect 24642 10906 24698 10908
rect 24722 10906 24778 10908
rect 24482 10854 24528 10906
rect 24528 10854 24538 10906
rect 24562 10854 24592 10906
rect 24592 10854 24604 10906
rect 24604 10854 24618 10906
rect 24642 10854 24656 10906
rect 24656 10854 24668 10906
rect 24668 10854 24698 10906
rect 24722 10854 24732 10906
rect 24732 10854 24778 10906
rect 24482 10852 24538 10854
rect 24562 10852 24618 10854
rect 24642 10852 24698 10854
rect 24722 10852 24778 10854
rect 32324 10906 32380 10908
rect 32404 10906 32460 10908
rect 32484 10906 32540 10908
rect 32564 10906 32620 10908
rect 32324 10854 32370 10906
rect 32370 10854 32380 10906
rect 32404 10854 32434 10906
rect 32434 10854 32446 10906
rect 32446 10854 32460 10906
rect 32484 10854 32498 10906
rect 32498 10854 32510 10906
rect 32510 10854 32540 10906
rect 32564 10854 32574 10906
rect 32574 10854 32620 10906
rect 32324 10852 32380 10854
rect 32404 10852 32460 10854
rect 32484 10852 32540 10854
rect 32564 10852 32620 10854
rect 4877 10362 4933 10364
rect 4957 10362 5013 10364
rect 5037 10362 5093 10364
rect 5117 10362 5173 10364
rect 4877 10310 4923 10362
rect 4923 10310 4933 10362
rect 4957 10310 4987 10362
rect 4987 10310 4999 10362
rect 4999 10310 5013 10362
rect 5037 10310 5051 10362
rect 5051 10310 5063 10362
rect 5063 10310 5093 10362
rect 5117 10310 5127 10362
rect 5127 10310 5173 10362
rect 4877 10308 4933 10310
rect 4957 10308 5013 10310
rect 5037 10308 5093 10310
rect 5117 10308 5173 10310
rect 12719 10362 12775 10364
rect 12799 10362 12855 10364
rect 12879 10362 12935 10364
rect 12959 10362 13015 10364
rect 12719 10310 12765 10362
rect 12765 10310 12775 10362
rect 12799 10310 12829 10362
rect 12829 10310 12841 10362
rect 12841 10310 12855 10362
rect 12879 10310 12893 10362
rect 12893 10310 12905 10362
rect 12905 10310 12935 10362
rect 12959 10310 12969 10362
rect 12969 10310 13015 10362
rect 12719 10308 12775 10310
rect 12799 10308 12855 10310
rect 12879 10308 12935 10310
rect 12959 10308 13015 10310
rect 20561 10362 20617 10364
rect 20641 10362 20697 10364
rect 20721 10362 20777 10364
rect 20801 10362 20857 10364
rect 20561 10310 20607 10362
rect 20607 10310 20617 10362
rect 20641 10310 20671 10362
rect 20671 10310 20683 10362
rect 20683 10310 20697 10362
rect 20721 10310 20735 10362
rect 20735 10310 20747 10362
rect 20747 10310 20777 10362
rect 20801 10310 20811 10362
rect 20811 10310 20857 10362
rect 20561 10308 20617 10310
rect 20641 10308 20697 10310
rect 20721 10308 20777 10310
rect 20801 10308 20857 10310
rect 28403 10362 28459 10364
rect 28483 10362 28539 10364
rect 28563 10362 28619 10364
rect 28643 10362 28699 10364
rect 28403 10310 28449 10362
rect 28449 10310 28459 10362
rect 28483 10310 28513 10362
rect 28513 10310 28525 10362
rect 28525 10310 28539 10362
rect 28563 10310 28577 10362
rect 28577 10310 28589 10362
rect 28589 10310 28619 10362
rect 28643 10310 28653 10362
rect 28653 10310 28699 10362
rect 28403 10308 28459 10310
rect 28483 10308 28539 10310
rect 28563 10308 28619 10310
rect 28643 10308 28699 10310
rect 8798 9818 8854 9820
rect 8878 9818 8934 9820
rect 8958 9818 9014 9820
rect 9038 9818 9094 9820
rect 8798 9766 8844 9818
rect 8844 9766 8854 9818
rect 8878 9766 8908 9818
rect 8908 9766 8920 9818
rect 8920 9766 8934 9818
rect 8958 9766 8972 9818
rect 8972 9766 8984 9818
rect 8984 9766 9014 9818
rect 9038 9766 9048 9818
rect 9048 9766 9094 9818
rect 8798 9764 8854 9766
rect 8878 9764 8934 9766
rect 8958 9764 9014 9766
rect 9038 9764 9094 9766
rect 16640 9818 16696 9820
rect 16720 9818 16776 9820
rect 16800 9818 16856 9820
rect 16880 9818 16936 9820
rect 16640 9766 16686 9818
rect 16686 9766 16696 9818
rect 16720 9766 16750 9818
rect 16750 9766 16762 9818
rect 16762 9766 16776 9818
rect 16800 9766 16814 9818
rect 16814 9766 16826 9818
rect 16826 9766 16856 9818
rect 16880 9766 16890 9818
rect 16890 9766 16936 9818
rect 16640 9764 16696 9766
rect 16720 9764 16776 9766
rect 16800 9764 16856 9766
rect 16880 9764 16936 9766
rect 24482 9818 24538 9820
rect 24562 9818 24618 9820
rect 24642 9818 24698 9820
rect 24722 9818 24778 9820
rect 24482 9766 24528 9818
rect 24528 9766 24538 9818
rect 24562 9766 24592 9818
rect 24592 9766 24604 9818
rect 24604 9766 24618 9818
rect 24642 9766 24656 9818
rect 24656 9766 24668 9818
rect 24668 9766 24698 9818
rect 24722 9766 24732 9818
rect 24732 9766 24778 9818
rect 24482 9764 24538 9766
rect 24562 9764 24618 9766
rect 24642 9764 24698 9766
rect 24722 9764 24778 9766
rect 32324 9818 32380 9820
rect 32404 9818 32460 9820
rect 32484 9818 32540 9820
rect 32564 9818 32620 9820
rect 32324 9766 32370 9818
rect 32370 9766 32380 9818
rect 32404 9766 32434 9818
rect 32434 9766 32446 9818
rect 32446 9766 32460 9818
rect 32484 9766 32498 9818
rect 32498 9766 32510 9818
rect 32510 9766 32540 9818
rect 32564 9766 32574 9818
rect 32574 9766 32620 9818
rect 32324 9764 32380 9766
rect 32404 9764 32460 9766
rect 32484 9764 32540 9766
rect 32564 9764 32620 9766
rect 4877 9274 4933 9276
rect 4957 9274 5013 9276
rect 5037 9274 5093 9276
rect 5117 9274 5173 9276
rect 4877 9222 4923 9274
rect 4923 9222 4933 9274
rect 4957 9222 4987 9274
rect 4987 9222 4999 9274
rect 4999 9222 5013 9274
rect 5037 9222 5051 9274
rect 5051 9222 5063 9274
rect 5063 9222 5093 9274
rect 5117 9222 5127 9274
rect 5127 9222 5173 9274
rect 4877 9220 4933 9222
rect 4957 9220 5013 9222
rect 5037 9220 5093 9222
rect 5117 9220 5173 9222
rect 12719 9274 12775 9276
rect 12799 9274 12855 9276
rect 12879 9274 12935 9276
rect 12959 9274 13015 9276
rect 12719 9222 12765 9274
rect 12765 9222 12775 9274
rect 12799 9222 12829 9274
rect 12829 9222 12841 9274
rect 12841 9222 12855 9274
rect 12879 9222 12893 9274
rect 12893 9222 12905 9274
rect 12905 9222 12935 9274
rect 12959 9222 12969 9274
rect 12969 9222 13015 9274
rect 12719 9220 12775 9222
rect 12799 9220 12855 9222
rect 12879 9220 12935 9222
rect 12959 9220 13015 9222
rect 20561 9274 20617 9276
rect 20641 9274 20697 9276
rect 20721 9274 20777 9276
rect 20801 9274 20857 9276
rect 20561 9222 20607 9274
rect 20607 9222 20617 9274
rect 20641 9222 20671 9274
rect 20671 9222 20683 9274
rect 20683 9222 20697 9274
rect 20721 9222 20735 9274
rect 20735 9222 20747 9274
rect 20747 9222 20777 9274
rect 20801 9222 20811 9274
rect 20811 9222 20857 9274
rect 20561 9220 20617 9222
rect 20641 9220 20697 9222
rect 20721 9220 20777 9222
rect 20801 9220 20857 9222
rect 28403 9274 28459 9276
rect 28483 9274 28539 9276
rect 28563 9274 28619 9276
rect 28643 9274 28699 9276
rect 28403 9222 28449 9274
rect 28449 9222 28459 9274
rect 28483 9222 28513 9274
rect 28513 9222 28525 9274
rect 28525 9222 28539 9274
rect 28563 9222 28577 9274
rect 28577 9222 28589 9274
rect 28589 9222 28619 9274
rect 28643 9222 28653 9274
rect 28653 9222 28699 9274
rect 28403 9220 28459 9222
rect 28483 9220 28539 9222
rect 28563 9220 28619 9222
rect 28643 9220 28699 9222
rect 8798 8730 8854 8732
rect 8878 8730 8934 8732
rect 8958 8730 9014 8732
rect 9038 8730 9094 8732
rect 8798 8678 8844 8730
rect 8844 8678 8854 8730
rect 8878 8678 8908 8730
rect 8908 8678 8920 8730
rect 8920 8678 8934 8730
rect 8958 8678 8972 8730
rect 8972 8678 8984 8730
rect 8984 8678 9014 8730
rect 9038 8678 9048 8730
rect 9048 8678 9094 8730
rect 8798 8676 8854 8678
rect 8878 8676 8934 8678
rect 8958 8676 9014 8678
rect 9038 8676 9094 8678
rect 16640 8730 16696 8732
rect 16720 8730 16776 8732
rect 16800 8730 16856 8732
rect 16880 8730 16936 8732
rect 16640 8678 16686 8730
rect 16686 8678 16696 8730
rect 16720 8678 16750 8730
rect 16750 8678 16762 8730
rect 16762 8678 16776 8730
rect 16800 8678 16814 8730
rect 16814 8678 16826 8730
rect 16826 8678 16856 8730
rect 16880 8678 16890 8730
rect 16890 8678 16936 8730
rect 16640 8676 16696 8678
rect 16720 8676 16776 8678
rect 16800 8676 16856 8678
rect 16880 8676 16936 8678
rect 24482 8730 24538 8732
rect 24562 8730 24618 8732
rect 24642 8730 24698 8732
rect 24722 8730 24778 8732
rect 24482 8678 24528 8730
rect 24528 8678 24538 8730
rect 24562 8678 24592 8730
rect 24592 8678 24604 8730
rect 24604 8678 24618 8730
rect 24642 8678 24656 8730
rect 24656 8678 24668 8730
rect 24668 8678 24698 8730
rect 24722 8678 24732 8730
rect 24732 8678 24778 8730
rect 24482 8676 24538 8678
rect 24562 8676 24618 8678
rect 24642 8676 24698 8678
rect 24722 8676 24778 8678
rect 32324 8730 32380 8732
rect 32404 8730 32460 8732
rect 32484 8730 32540 8732
rect 32564 8730 32620 8732
rect 32324 8678 32370 8730
rect 32370 8678 32380 8730
rect 32404 8678 32434 8730
rect 32434 8678 32446 8730
rect 32446 8678 32460 8730
rect 32484 8678 32498 8730
rect 32498 8678 32510 8730
rect 32510 8678 32540 8730
rect 32564 8678 32574 8730
rect 32574 8678 32620 8730
rect 32324 8676 32380 8678
rect 32404 8676 32460 8678
rect 32484 8676 32540 8678
rect 32564 8676 32620 8678
rect 4877 8186 4933 8188
rect 4957 8186 5013 8188
rect 5037 8186 5093 8188
rect 5117 8186 5173 8188
rect 4877 8134 4923 8186
rect 4923 8134 4933 8186
rect 4957 8134 4987 8186
rect 4987 8134 4999 8186
rect 4999 8134 5013 8186
rect 5037 8134 5051 8186
rect 5051 8134 5063 8186
rect 5063 8134 5093 8186
rect 5117 8134 5127 8186
rect 5127 8134 5173 8186
rect 4877 8132 4933 8134
rect 4957 8132 5013 8134
rect 5037 8132 5093 8134
rect 5117 8132 5173 8134
rect 12719 8186 12775 8188
rect 12799 8186 12855 8188
rect 12879 8186 12935 8188
rect 12959 8186 13015 8188
rect 12719 8134 12765 8186
rect 12765 8134 12775 8186
rect 12799 8134 12829 8186
rect 12829 8134 12841 8186
rect 12841 8134 12855 8186
rect 12879 8134 12893 8186
rect 12893 8134 12905 8186
rect 12905 8134 12935 8186
rect 12959 8134 12969 8186
rect 12969 8134 13015 8186
rect 12719 8132 12775 8134
rect 12799 8132 12855 8134
rect 12879 8132 12935 8134
rect 12959 8132 13015 8134
rect 20561 8186 20617 8188
rect 20641 8186 20697 8188
rect 20721 8186 20777 8188
rect 20801 8186 20857 8188
rect 20561 8134 20607 8186
rect 20607 8134 20617 8186
rect 20641 8134 20671 8186
rect 20671 8134 20683 8186
rect 20683 8134 20697 8186
rect 20721 8134 20735 8186
rect 20735 8134 20747 8186
rect 20747 8134 20777 8186
rect 20801 8134 20811 8186
rect 20811 8134 20857 8186
rect 20561 8132 20617 8134
rect 20641 8132 20697 8134
rect 20721 8132 20777 8134
rect 20801 8132 20857 8134
rect 28403 8186 28459 8188
rect 28483 8186 28539 8188
rect 28563 8186 28619 8188
rect 28643 8186 28699 8188
rect 28403 8134 28449 8186
rect 28449 8134 28459 8186
rect 28483 8134 28513 8186
rect 28513 8134 28525 8186
rect 28525 8134 28539 8186
rect 28563 8134 28577 8186
rect 28577 8134 28589 8186
rect 28589 8134 28619 8186
rect 28643 8134 28653 8186
rect 28653 8134 28699 8186
rect 28403 8132 28459 8134
rect 28483 8132 28539 8134
rect 28563 8132 28619 8134
rect 28643 8132 28699 8134
rect 8798 7642 8854 7644
rect 8878 7642 8934 7644
rect 8958 7642 9014 7644
rect 9038 7642 9094 7644
rect 8798 7590 8844 7642
rect 8844 7590 8854 7642
rect 8878 7590 8908 7642
rect 8908 7590 8920 7642
rect 8920 7590 8934 7642
rect 8958 7590 8972 7642
rect 8972 7590 8984 7642
rect 8984 7590 9014 7642
rect 9038 7590 9048 7642
rect 9048 7590 9094 7642
rect 8798 7588 8854 7590
rect 8878 7588 8934 7590
rect 8958 7588 9014 7590
rect 9038 7588 9094 7590
rect 16640 7642 16696 7644
rect 16720 7642 16776 7644
rect 16800 7642 16856 7644
rect 16880 7642 16936 7644
rect 16640 7590 16686 7642
rect 16686 7590 16696 7642
rect 16720 7590 16750 7642
rect 16750 7590 16762 7642
rect 16762 7590 16776 7642
rect 16800 7590 16814 7642
rect 16814 7590 16826 7642
rect 16826 7590 16856 7642
rect 16880 7590 16890 7642
rect 16890 7590 16936 7642
rect 16640 7588 16696 7590
rect 16720 7588 16776 7590
rect 16800 7588 16856 7590
rect 16880 7588 16936 7590
rect 24482 7642 24538 7644
rect 24562 7642 24618 7644
rect 24642 7642 24698 7644
rect 24722 7642 24778 7644
rect 24482 7590 24528 7642
rect 24528 7590 24538 7642
rect 24562 7590 24592 7642
rect 24592 7590 24604 7642
rect 24604 7590 24618 7642
rect 24642 7590 24656 7642
rect 24656 7590 24668 7642
rect 24668 7590 24698 7642
rect 24722 7590 24732 7642
rect 24732 7590 24778 7642
rect 24482 7588 24538 7590
rect 24562 7588 24618 7590
rect 24642 7588 24698 7590
rect 24722 7588 24778 7590
rect 32324 7642 32380 7644
rect 32404 7642 32460 7644
rect 32484 7642 32540 7644
rect 32564 7642 32620 7644
rect 32324 7590 32370 7642
rect 32370 7590 32380 7642
rect 32404 7590 32434 7642
rect 32434 7590 32446 7642
rect 32446 7590 32460 7642
rect 32484 7590 32498 7642
rect 32498 7590 32510 7642
rect 32510 7590 32540 7642
rect 32564 7590 32574 7642
rect 32574 7590 32620 7642
rect 32324 7588 32380 7590
rect 32404 7588 32460 7590
rect 32484 7588 32540 7590
rect 32564 7588 32620 7590
rect 4877 7098 4933 7100
rect 4957 7098 5013 7100
rect 5037 7098 5093 7100
rect 5117 7098 5173 7100
rect 4877 7046 4923 7098
rect 4923 7046 4933 7098
rect 4957 7046 4987 7098
rect 4987 7046 4999 7098
rect 4999 7046 5013 7098
rect 5037 7046 5051 7098
rect 5051 7046 5063 7098
rect 5063 7046 5093 7098
rect 5117 7046 5127 7098
rect 5127 7046 5173 7098
rect 4877 7044 4933 7046
rect 4957 7044 5013 7046
rect 5037 7044 5093 7046
rect 5117 7044 5173 7046
rect 12719 7098 12775 7100
rect 12799 7098 12855 7100
rect 12879 7098 12935 7100
rect 12959 7098 13015 7100
rect 12719 7046 12765 7098
rect 12765 7046 12775 7098
rect 12799 7046 12829 7098
rect 12829 7046 12841 7098
rect 12841 7046 12855 7098
rect 12879 7046 12893 7098
rect 12893 7046 12905 7098
rect 12905 7046 12935 7098
rect 12959 7046 12969 7098
rect 12969 7046 13015 7098
rect 12719 7044 12775 7046
rect 12799 7044 12855 7046
rect 12879 7044 12935 7046
rect 12959 7044 13015 7046
rect 20561 7098 20617 7100
rect 20641 7098 20697 7100
rect 20721 7098 20777 7100
rect 20801 7098 20857 7100
rect 20561 7046 20607 7098
rect 20607 7046 20617 7098
rect 20641 7046 20671 7098
rect 20671 7046 20683 7098
rect 20683 7046 20697 7098
rect 20721 7046 20735 7098
rect 20735 7046 20747 7098
rect 20747 7046 20777 7098
rect 20801 7046 20811 7098
rect 20811 7046 20857 7098
rect 20561 7044 20617 7046
rect 20641 7044 20697 7046
rect 20721 7044 20777 7046
rect 20801 7044 20857 7046
rect 28403 7098 28459 7100
rect 28483 7098 28539 7100
rect 28563 7098 28619 7100
rect 28643 7098 28699 7100
rect 28403 7046 28449 7098
rect 28449 7046 28459 7098
rect 28483 7046 28513 7098
rect 28513 7046 28525 7098
rect 28525 7046 28539 7098
rect 28563 7046 28577 7098
rect 28577 7046 28589 7098
rect 28589 7046 28619 7098
rect 28643 7046 28653 7098
rect 28653 7046 28699 7098
rect 28403 7044 28459 7046
rect 28483 7044 28539 7046
rect 28563 7044 28619 7046
rect 28643 7044 28699 7046
rect 8798 6554 8854 6556
rect 8878 6554 8934 6556
rect 8958 6554 9014 6556
rect 9038 6554 9094 6556
rect 8798 6502 8844 6554
rect 8844 6502 8854 6554
rect 8878 6502 8908 6554
rect 8908 6502 8920 6554
rect 8920 6502 8934 6554
rect 8958 6502 8972 6554
rect 8972 6502 8984 6554
rect 8984 6502 9014 6554
rect 9038 6502 9048 6554
rect 9048 6502 9094 6554
rect 8798 6500 8854 6502
rect 8878 6500 8934 6502
rect 8958 6500 9014 6502
rect 9038 6500 9094 6502
rect 16640 6554 16696 6556
rect 16720 6554 16776 6556
rect 16800 6554 16856 6556
rect 16880 6554 16936 6556
rect 16640 6502 16686 6554
rect 16686 6502 16696 6554
rect 16720 6502 16750 6554
rect 16750 6502 16762 6554
rect 16762 6502 16776 6554
rect 16800 6502 16814 6554
rect 16814 6502 16826 6554
rect 16826 6502 16856 6554
rect 16880 6502 16890 6554
rect 16890 6502 16936 6554
rect 16640 6500 16696 6502
rect 16720 6500 16776 6502
rect 16800 6500 16856 6502
rect 16880 6500 16936 6502
rect 24482 6554 24538 6556
rect 24562 6554 24618 6556
rect 24642 6554 24698 6556
rect 24722 6554 24778 6556
rect 24482 6502 24528 6554
rect 24528 6502 24538 6554
rect 24562 6502 24592 6554
rect 24592 6502 24604 6554
rect 24604 6502 24618 6554
rect 24642 6502 24656 6554
rect 24656 6502 24668 6554
rect 24668 6502 24698 6554
rect 24722 6502 24732 6554
rect 24732 6502 24778 6554
rect 24482 6500 24538 6502
rect 24562 6500 24618 6502
rect 24642 6500 24698 6502
rect 24722 6500 24778 6502
rect 32324 6554 32380 6556
rect 32404 6554 32460 6556
rect 32484 6554 32540 6556
rect 32564 6554 32620 6556
rect 32324 6502 32370 6554
rect 32370 6502 32380 6554
rect 32404 6502 32434 6554
rect 32434 6502 32446 6554
rect 32446 6502 32460 6554
rect 32484 6502 32498 6554
rect 32498 6502 32510 6554
rect 32510 6502 32540 6554
rect 32564 6502 32574 6554
rect 32574 6502 32620 6554
rect 32324 6500 32380 6502
rect 32404 6500 32460 6502
rect 32484 6500 32540 6502
rect 32564 6500 32620 6502
rect 4877 6010 4933 6012
rect 4957 6010 5013 6012
rect 5037 6010 5093 6012
rect 5117 6010 5173 6012
rect 4877 5958 4923 6010
rect 4923 5958 4933 6010
rect 4957 5958 4987 6010
rect 4987 5958 4999 6010
rect 4999 5958 5013 6010
rect 5037 5958 5051 6010
rect 5051 5958 5063 6010
rect 5063 5958 5093 6010
rect 5117 5958 5127 6010
rect 5127 5958 5173 6010
rect 4877 5956 4933 5958
rect 4957 5956 5013 5958
rect 5037 5956 5093 5958
rect 5117 5956 5173 5958
rect 12719 6010 12775 6012
rect 12799 6010 12855 6012
rect 12879 6010 12935 6012
rect 12959 6010 13015 6012
rect 12719 5958 12765 6010
rect 12765 5958 12775 6010
rect 12799 5958 12829 6010
rect 12829 5958 12841 6010
rect 12841 5958 12855 6010
rect 12879 5958 12893 6010
rect 12893 5958 12905 6010
rect 12905 5958 12935 6010
rect 12959 5958 12969 6010
rect 12969 5958 13015 6010
rect 12719 5956 12775 5958
rect 12799 5956 12855 5958
rect 12879 5956 12935 5958
rect 12959 5956 13015 5958
rect 20561 6010 20617 6012
rect 20641 6010 20697 6012
rect 20721 6010 20777 6012
rect 20801 6010 20857 6012
rect 20561 5958 20607 6010
rect 20607 5958 20617 6010
rect 20641 5958 20671 6010
rect 20671 5958 20683 6010
rect 20683 5958 20697 6010
rect 20721 5958 20735 6010
rect 20735 5958 20747 6010
rect 20747 5958 20777 6010
rect 20801 5958 20811 6010
rect 20811 5958 20857 6010
rect 20561 5956 20617 5958
rect 20641 5956 20697 5958
rect 20721 5956 20777 5958
rect 20801 5956 20857 5958
rect 28403 6010 28459 6012
rect 28483 6010 28539 6012
rect 28563 6010 28619 6012
rect 28643 6010 28699 6012
rect 28403 5958 28449 6010
rect 28449 5958 28459 6010
rect 28483 5958 28513 6010
rect 28513 5958 28525 6010
rect 28525 5958 28539 6010
rect 28563 5958 28577 6010
rect 28577 5958 28589 6010
rect 28589 5958 28619 6010
rect 28643 5958 28653 6010
rect 28653 5958 28699 6010
rect 28403 5956 28459 5958
rect 28483 5956 28539 5958
rect 28563 5956 28619 5958
rect 28643 5956 28699 5958
rect 8798 5466 8854 5468
rect 8878 5466 8934 5468
rect 8958 5466 9014 5468
rect 9038 5466 9094 5468
rect 8798 5414 8844 5466
rect 8844 5414 8854 5466
rect 8878 5414 8908 5466
rect 8908 5414 8920 5466
rect 8920 5414 8934 5466
rect 8958 5414 8972 5466
rect 8972 5414 8984 5466
rect 8984 5414 9014 5466
rect 9038 5414 9048 5466
rect 9048 5414 9094 5466
rect 8798 5412 8854 5414
rect 8878 5412 8934 5414
rect 8958 5412 9014 5414
rect 9038 5412 9094 5414
rect 16640 5466 16696 5468
rect 16720 5466 16776 5468
rect 16800 5466 16856 5468
rect 16880 5466 16936 5468
rect 16640 5414 16686 5466
rect 16686 5414 16696 5466
rect 16720 5414 16750 5466
rect 16750 5414 16762 5466
rect 16762 5414 16776 5466
rect 16800 5414 16814 5466
rect 16814 5414 16826 5466
rect 16826 5414 16856 5466
rect 16880 5414 16890 5466
rect 16890 5414 16936 5466
rect 16640 5412 16696 5414
rect 16720 5412 16776 5414
rect 16800 5412 16856 5414
rect 16880 5412 16936 5414
rect 24482 5466 24538 5468
rect 24562 5466 24618 5468
rect 24642 5466 24698 5468
rect 24722 5466 24778 5468
rect 24482 5414 24528 5466
rect 24528 5414 24538 5466
rect 24562 5414 24592 5466
rect 24592 5414 24604 5466
rect 24604 5414 24618 5466
rect 24642 5414 24656 5466
rect 24656 5414 24668 5466
rect 24668 5414 24698 5466
rect 24722 5414 24732 5466
rect 24732 5414 24778 5466
rect 24482 5412 24538 5414
rect 24562 5412 24618 5414
rect 24642 5412 24698 5414
rect 24722 5412 24778 5414
rect 32324 5466 32380 5468
rect 32404 5466 32460 5468
rect 32484 5466 32540 5468
rect 32564 5466 32620 5468
rect 32324 5414 32370 5466
rect 32370 5414 32380 5466
rect 32404 5414 32434 5466
rect 32434 5414 32446 5466
rect 32446 5414 32460 5466
rect 32484 5414 32498 5466
rect 32498 5414 32510 5466
rect 32510 5414 32540 5466
rect 32564 5414 32574 5466
rect 32574 5414 32620 5466
rect 32324 5412 32380 5414
rect 32404 5412 32460 5414
rect 32484 5412 32540 5414
rect 32564 5412 32620 5414
rect 4877 4922 4933 4924
rect 4957 4922 5013 4924
rect 5037 4922 5093 4924
rect 5117 4922 5173 4924
rect 4877 4870 4923 4922
rect 4923 4870 4933 4922
rect 4957 4870 4987 4922
rect 4987 4870 4999 4922
rect 4999 4870 5013 4922
rect 5037 4870 5051 4922
rect 5051 4870 5063 4922
rect 5063 4870 5093 4922
rect 5117 4870 5127 4922
rect 5127 4870 5173 4922
rect 4877 4868 4933 4870
rect 4957 4868 5013 4870
rect 5037 4868 5093 4870
rect 5117 4868 5173 4870
rect 12719 4922 12775 4924
rect 12799 4922 12855 4924
rect 12879 4922 12935 4924
rect 12959 4922 13015 4924
rect 12719 4870 12765 4922
rect 12765 4870 12775 4922
rect 12799 4870 12829 4922
rect 12829 4870 12841 4922
rect 12841 4870 12855 4922
rect 12879 4870 12893 4922
rect 12893 4870 12905 4922
rect 12905 4870 12935 4922
rect 12959 4870 12969 4922
rect 12969 4870 13015 4922
rect 12719 4868 12775 4870
rect 12799 4868 12855 4870
rect 12879 4868 12935 4870
rect 12959 4868 13015 4870
rect 20561 4922 20617 4924
rect 20641 4922 20697 4924
rect 20721 4922 20777 4924
rect 20801 4922 20857 4924
rect 20561 4870 20607 4922
rect 20607 4870 20617 4922
rect 20641 4870 20671 4922
rect 20671 4870 20683 4922
rect 20683 4870 20697 4922
rect 20721 4870 20735 4922
rect 20735 4870 20747 4922
rect 20747 4870 20777 4922
rect 20801 4870 20811 4922
rect 20811 4870 20857 4922
rect 20561 4868 20617 4870
rect 20641 4868 20697 4870
rect 20721 4868 20777 4870
rect 20801 4868 20857 4870
rect 28403 4922 28459 4924
rect 28483 4922 28539 4924
rect 28563 4922 28619 4924
rect 28643 4922 28699 4924
rect 28403 4870 28449 4922
rect 28449 4870 28459 4922
rect 28483 4870 28513 4922
rect 28513 4870 28525 4922
rect 28525 4870 28539 4922
rect 28563 4870 28577 4922
rect 28577 4870 28589 4922
rect 28589 4870 28619 4922
rect 28643 4870 28653 4922
rect 28653 4870 28699 4922
rect 28403 4868 28459 4870
rect 28483 4868 28539 4870
rect 28563 4868 28619 4870
rect 28643 4868 28699 4870
rect 8798 4378 8854 4380
rect 8878 4378 8934 4380
rect 8958 4378 9014 4380
rect 9038 4378 9094 4380
rect 8798 4326 8844 4378
rect 8844 4326 8854 4378
rect 8878 4326 8908 4378
rect 8908 4326 8920 4378
rect 8920 4326 8934 4378
rect 8958 4326 8972 4378
rect 8972 4326 8984 4378
rect 8984 4326 9014 4378
rect 9038 4326 9048 4378
rect 9048 4326 9094 4378
rect 8798 4324 8854 4326
rect 8878 4324 8934 4326
rect 8958 4324 9014 4326
rect 9038 4324 9094 4326
rect 16640 4378 16696 4380
rect 16720 4378 16776 4380
rect 16800 4378 16856 4380
rect 16880 4378 16936 4380
rect 16640 4326 16686 4378
rect 16686 4326 16696 4378
rect 16720 4326 16750 4378
rect 16750 4326 16762 4378
rect 16762 4326 16776 4378
rect 16800 4326 16814 4378
rect 16814 4326 16826 4378
rect 16826 4326 16856 4378
rect 16880 4326 16890 4378
rect 16890 4326 16936 4378
rect 16640 4324 16696 4326
rect 16720 4324 16776 4326
rect 16800 4324 16856 4326
rect 16880 4324 16936 4326
rect 24482 4378 24538 4380
rect 24562 4378 24618 4380
rect 24642 4378 24698 4380
rect 24722 4378 24778 4380
rect 24482 4326 24528 4378
rect 24528 4326 24538 4378
rect 24562 4326 24592 4378
rect 24592 4326 24604 4378
rect 24604 4326 24618 4378
rect 24642 4326 24656 4378
rect 24656 4326 24668 4378
rect 24668 4326 24698 4378
rect 24722 4326 24732 4378
rect 24732 4326 24778 4378
rect 24482 4324 24538 4326
rect 24562 4324 24618 4326
rect 24642 4324 24698 4326
rect 24722 4324 24778 4326
rect 32324 4378 32380 4380
rect 32404 4378 32460 4380
rect 32484 4378 32540 4380
rect 32564 4378 32620 4380
rect 32324 4326 32370 4378
rect 32370 4326 32380 4378
rect 32404 4326 32434 4378
rect 32434 4326 32446 4378
rect 32446 4326 32460 4378
rect 32484 4326 32498 4378
rect 32498 4326 32510 4378
rect 32510 4326 32540 4378
rect 32564 4326 32574 4378
rect 32574 4326 32620 4378
rect 32324 4324 32380 4326
rect 32404 4324 32460 4326
rect 32484 4324 32540 4326
rect 32564 4324 32620 4326
rect 4877 3834 4933 3836
rect 4957 3834 5013 3836
rect 5037 3834 5093 3836
rect 5117 3834 5173 3836
rect 4877 3782 4923 3834
rect 4923 3782 4933 3834
rect 4957 3782 4987 3834
rect 4987 3782 4999 3834
rect 4999 3782 5013 3834
rect 5037 3782 5051 3834
rect 5051 3782 5063 3834
rect 5063 3782 5093 3834
rect 5117 3782 5127 3834
rect 5127 3782 5173 3834
rect 4877 3780 4933 3782
rect 4957 3780 5013 3782
rect 5037 3780 5093 3782
rect 5117 3780 5173 3782
rect 12719 3834 12775 3836
rect 12799 3834 12855 3836
rect 12879 3834 12935 3836
rect 12959 3834 13015 3836
rect 12719 3782 12765 3834
rect 12765 3782 12775 3834
rect 12799 3782 12829 3834
rect 12829 3782 12841 3834
rect 12841 3782 12855 3834
rect 12879 3782 12893 3834
rect 12893 3782 12905 3834
rect 12905 3782 12935 3834
rect 12959 3782 12969 3834
rect 12969 3782 13015 3834
rect 12719 3780 12775 3782
rect 12799 3780 12855 3782
rect 12879 3780 12935 3782
rect 12959 3780 13015 3782
rect 20561 3834 20617 3836
rect 20641 3834 20697 3836
rect 20721 3834 20777 3836
rect 20801 3834 20857 3836
rect 20561 3782 20607 3834
rect 20607 3782 20617 3834
rect 20641 3782 20671 3834
rect 20671 3782 20683 3834
rect 20683 3782 20697 3834
rect 20721 3782 20735 3834
rect 20735 3782 20747 3834
rect 20747 3782 20777 3834
rect 20801 3782 20811 3834
rect 20811 3782 20857 3834
rect 20561 3780 20617 3782
rect 20641 3780 20697 3782
rect 20721 3780 20777 3782
rect 20801 3780 20857 3782
rect 28403 3834 28459 3836
rect 28483 3834 28539 3836
rect 28563 3834 28619 3836
rect 28643 3834 28699 3836
rect 28403 3782 28449 3834
rect 28449 3782 28459 3834
rect 28483 3782 28513 3834
rect 28513 3782 28525 3834
rect 28525 3782 28539 3834
rect 28563 3782 28577 3834
rect 28577 3782 28589 3834
rect 28589 3782 28619 3834
rect 28643 3782 28653 3834
rect 28653 3782 28699 3834
rect 28403 3780 28459 3782
rect 28483 3780 28539 3782
rect 28563 3780 28619 3782
rect 28643 3780 28699 3782
rect 8798 3290 8854 3292
rect 8878 3290 8934 3292
rect 8958 3290 9014 3292
rect 9038 3290 9094 3292
rect 8798 3238 8844 3290
rect 8844 3238 8854 3290
rect 8878 3238 8908 3290
rect 8908 3238 8920 3290
rect 8920 3238 8934 3290
rect 8958 3238 8972 3290
rect 8972 3238 8984 3290
rect 8984 3238 9014 3290
rect 9038 3238 9048 3290
rect 9048 3238 9094 3290
rect 8798 3236 8854 3238
rect 8878 3236 8934 3238
rect 8958 3236 9014 3238
rect 9038 3236 9094 3238
rect 16640 3290 16696 3292
rect 16720 3290 16776 3292
rect 16800 3290 16856 3292
rect 16880 3290 16936 3292
rect 16640 3238 16686 3290
rect 16686 3238 16696 3290
rect 16720 3238 16750 3290
rect 16750 3238 16762 3290
rect 16762 3238 16776 3290
rect 16800 3238 16814 3290
rect 16814 3238 16826 3290
rect 16826 3238 16856 3290
rect 16880 3238 16890 3290
rect 16890 3238 16936 3290
rect 16640 3236 16696 3238
rect 16720 3236 16776 3238
rect 16800 3236 16856 3238
rect 16880 3236 16936 3238
rect 24482 3290 24538 3292
rect 24562 3290 24618 3292
rect 24642 3290 24698 3292
rect 24722 3290 24778 3292
rect 24482 3238 24528 3290
rect 24528 3238 24538 3290
rect 24562 3238 24592 3290
rect 24592 3238 24604 3290
rect 24604 3238 24618 3290
rect 24642 3238 24656 3290
rect 24656 3238 24668 3290
rect 24668 3238 24698 3290
rect 24722 3238 24732 3290
rect 24732 3238 24778 3290
rect 24482 3236 24538 3238
rect 24562 3236 24618 3238
rect 24642 3236 24698 3238
rect 24722 3236 24778 3238
rect 32324 3290 32380 3292
rect 32404 3290 32460 3292
rect 32484 3290 32540 3292
rect 32564 3290 32620 3292
rect 32324 3238 32370 3290
rect 32370 3238 32380 3290
rect 32404 3238 32434 3290
rect 32434 3238 32446 3290
rect 32446 3238 32460 3290
rect 32484 3238 32498 3290
rect 32498 3238 32510 3290
rect 32510 3238 32540 3290
rect 32564 3238 32574 3290
rect 32574 3238 32620 3290
rect 32324 3236 32380 3238
rect 32404 3236 32460 3238
rect 32484 3236 32540 3238
rect 32564 3236 32620 3238
rect 4877 2746 4933 2748
rect 4957 2746 5013 2748
rect 5037 2746 5093 2748
rect 5117 2746 5173 2748
rect 4877 2694 4923 2746
rect 4923 2694 4933 2746
rect 4957 2694 4987 2746
rect 4987 2694 4999 2746
rect 4999 2694 5013 2746
rect 5037 2694 5051 2746
rect 5051 2694 5063 2746
rect 5063 2694 5093 2746
rect 5117 2694 5127 2746
rect 5127 2694 5173 2746
rect 4877 2692 4933 2694
rect 4957 2692 5013 2694
rect 5037 2692 5093 2694
rect 5117 2692 5173 2694
rect 12719 2746 12775 2748
rect 12799 2746 12855 2748
rect 12879 2746 12935 2748
rect 12959 2746 13015 2748
rect 12719 2694 12765 2746
rect 12765 2694 12775 2746
rect 12799 2694 12829 2746
rect 12829 2694 12841 2746
rect 12841 2694 12855 2746
rect 12879 2694 12893 2746
rect 12893 2694 12905 2746
rect 12905 2694 12935 2746
rect 12959 2694 12969 2746
rect 12969 2694 13015 2746
rect 12719 2692 12775 2694
rect 12799 2692 12855 2694
rect 12879 2692 12935 2694
rect 12959 2692 13015 2694
rect 20561 2746 20617 2748
rect 20641 2746 20697 2748
rect 20721 2746 20777 2748
rect 20801 2746 20857 2748
rect 20561 2694 20607 2746
rect 20607 2694 20617 2746
rect 20641 2694 20671 2746
rect 20671 2694 20683 2746
rect 20683 2694 20697 2746
rect 20721 2694 20735 2746
rect 20735 2694 20747 2746
rect 20747 2694 20777 2746
rect 20801 2694 20811 2746
rect 20811 2694 20857 2746
rect 20561 2692 20617 2694
rect 20641 2692 20697 2694
rect 20721 2692 20777 2694
rect 20801 2692 20857 2694
rect 28403 2746 28459 2748
rect 28483 2746 28539 2748
rect 28563 2746 28619 2748
rect 28643 2746 28699 2748
rect 28403 2694 28449 2746
rect 28449 2694 28459 2746
rect 28483 2694 28513 2746
rect 28513 2694 28525 2746
rect 28525 2694 28539 2746
rect 28563 2694 28577 2746
rect 28577 2694 28589 2746
rect 28589 2694 28619 2746
rect 28643 2694 28653 2746
rect 28653 2694 28699 2746
rect 28403 2692 28459 2694
rect 28483 2692 28539 2694
rect 28563 2692 28619 2694
rect 28643 2692 28699 2694
rect 8798 2202 8854 2204
rect 8878 2202 8934 2204
rect 8958 2202 9014 2204
rect 9038 2202 9094 2204
rect 8798 2150 8844 2202
rect 8844 2150 8854 2202
rect 8878 2150 8908 2202
rect 8908 2150 8920 2202
rect 8920 2150 8934 2202
rect 8958 2150 8972 2202
rect 8972 2150 8984 2202
rect 8984 2150 9014 2202
rect 9038 2150 9048 2202
rect 9048 2150 9094 2202
rect 8798 2148 8854 2150
rect 8878 2148 8934 2150
rect 8958 2148 9014 2150
rect 9038 2148 9094 2150
rect 16640 2202 16696 2204
rect 16720 2202 16776 2204
rect 16800 2202 16856 2204
rect 16880 2202 16936 2204
rect 16640 2150 16686 2202
rect 16686 2150 16696 2202
rect 16720 2150 16750 2202
rect 16750 2150 16762 2202
rect 16762 2150 16776 2202
rect 16800 2150 16814 2202
rect 16814 2150 16826 2202
rect 16826 2150 16856 2202
rect 16880 2150 16890 2202
rect 16890 2150 16936 2202
rect 16640 2148 16696 2150
rect 16720 2148 16776 2150
rect 16800 2148 16856 2150
rect 16880 2148 16936 2150
rect 24482 2202 24538 2204
rect 24562 2202 24618 2204
rect 24642 2202 24698 2204
rect 24722 2202 24778 2204
rect 24482 2150 24528 2202
rect 24528 2150 24538 2202
rect 24562 2150 24592 2202
rect 24592 2150 24604 2202
rect 24604 2150 24618 2202
rect 24642 2150 24656 2202
rect 24656 2150 24668 2202
rect 24668 2150 24698 2202
rect 24722 2150 24732 2202
rect 24732 2150 24778 2202
rect 24482 2148 24538 2150
rect 24562 2148 24618 2150
rect 24642 2148 24698 2150
rect 24722 2148 24778 2150
rect 32324 2202 32380 2204
rect 32404 2202 32460 2204
rect 32484 2202 32540 2204
rect 32564 2202 32620 2204
rect 32324 2150 32370 2202
rect 32370 2150 32380 2202
rect 32404 2150 32434 2202
rect 32434 2150 32446 2202
rect 32446 2150 32460 2202
rect 32484 2150 32498 2202
rect 32498 2150 32510 2202
rect 32510 2150 32540 2202
rect 32564 2150 32574 2202
rect 32574 2150 32620 2202
rect 32324 2148 32380 2150
rect 32404 2148 32460 2150
rect 32484 2148 32540 2150
rect 32564 2148 32620 2150
rect 4877 1658 4933 1660
rect 4957 1658 5013 1660
rect 5037 1658 5093 1660
rect 5117 1658 5173 1660
rect 4877 1606 4923 1658
rect 4923 1606 4933 1658
rect 4957 1606 4987 1658
rect 4987 1606 4999 1658
rect 4999 1606 5013 1658
rect 5037 1606 5051 1658
rect 5051 1606 5063 1658
rect 5063 1606 5093 1658
rect 5117 1606 5127 1658
rect 5127 1606 5173 1658
rect 4877 1604 4933 1606
rect 4957 1604 5013 1606
rect 5037 1604 5093 1606
rect 5117 1604 5173 1606
rect 12719 1658 12775 1660
rect 12799 1658 12855 1660
rect 12879 1658 12935 1660
rect 12959 1658 13015 1660
rect 12719 1606 12765 1658
rect 12765 1606 12775 1658
rect 12799 1606 12829 1658
rect 12829 1606 12841 1658
rect 12841 1606 12855 1658
rect 12879 1606 12893 1658
rect 12893 1606 12905 1658
rect 12905 1606 12935 1658
rect 12959 1606 12969 1658
rect 12969 1606 13015 1658
rect 12719 1604 12775 1606
rect 12799 1604 12855 1606
rect 12879 1604 12935 1606
rect 12959 1604 13015 1606
rect 20561 1658 20617 1660
rect 20641 1658 20697 1660
rect 20721 1658 20777 1660
rect 20801 1658 20857 1660
rect 20561 1606 20607 1658
rect 20607 1606 20617 1658
rect 20641 1606 20671 1658
rect 20671 1606 20683 1658
rect 20683 1606 20697 1658
rect 20721 1606 20735 1658
rect 20735 1606 20747 1658
rect 20747 1606 20777 1658
rect 20801 1606 20811 1658
rect 20811 1606 20857 1658
rect 20561 1604 20617 1606
rect 20641 1604 20697 1606
rect 20721 1604 20777 1606
rect 20801 1604 20857 1606
rect 28403 1658 28459 1660
rect 28483 1658 28539 1660
rect 28563 1658 28619 1660
rect 28643 1658 28699 1660
rect 28403 1606 28449 1658
rect 28449 1606 28459 1658
rect 28483 1606 28513 1658
rect 28513 1606 28525 1658
rect 28525 1606 28539 1658
rect 28563 1606 28577 1658
rect 28577 1606 28589 1658
rect 28589 1606 28619 1658
rect 28643 1606 28653 1658
rect 28653 1606 28699 1658
rect 28403 1604 28459 1606
rect 28483 1604 28539 1606
rect 28563 1604 28619 1606
rect 28643 1604 28699 1606
rect 8798 1114 8854 1116
rect 8878 1114 8934 1116
rect 8958 1114 9014 1116
rect 9038 1114 9094 1116
rect 8798 1062 8844 1114
rect 8844 1062 8854 1114
rect 8878 1062 8908 1114
rect 8908 1062 8920 1114
rect 8920 1062 8934 1114
rect 8958 1062 8972 1114
rect 8972 1062 8984 1114
rect 8984 1062 9014 1114
rect 9038 1062 9048 1114
rect 9048 1062 9094 1114
rect 8798 1060 8854 1062
rect 8878 1060 8934 1062
rect 8958 1060 9014 1062
rect 9038 1060 9094 1062
rect 16640 1114 16696 1116
rect 16720 1114 16776 1116
rect 16800 1114 16856 1116
rect 16880 1114 16936 1116
rect 16640 1062 16686 1114
rect 16686 1062 16696 1114
rect 16720 1062 16750 1114
rect 16750 1062 16762 1114
rect 16762 1062 16776 1114
rect 16800 1062 16814 1114
rect 16814 1062 16826 1114
rect 16826 1062 16856 1114
rect 16880 1062 16890 1114
rect 16890 1062 16936 1114
rect 16640 1060 16696 1062
rect 16720 1060 16776 1062
rect 16800 1060 16856 1062
rect 16880 1060 16936 1062
rect 24482 1114 24538 1116
rect 24562 1114 24618 1116
rect 24642 1114 24698 1116
rect 24722 1114 24778 1116
rect 24482 1062 24528 1114
rect 24528 1062 24538 1114
rect 24562 1062 24592 1114
rect 24592 1062 24604 1114
rect 24604 1062 24618 1114
rect 24642 1062 24656 1114
rect 24656 1062 24668 1114
rect 24668 1062 24698 1114
rect 24722 1062 24732 1114
rect 24732 1062 24778 1114
rect 24482 1060 24538 1062
rect 24562 1060 24618 1062
rect 24642 1060 24698 1062
rect 24722 1060 24778 1062
rect 32324 1114 32380 1116
rect 32404 1114 32460 1116
rect 32484 1114 32540 1116
rect 32564 1114 32620 1116
rect 32324 1062 32370 1114
rect 32370 1062 32380 1114
rect 32404 1062 32434 1114
rect 32434 1062 32446 1114
rect 32446 1062 32460 1114
rect 32484 1062 32498 1114
rect 32498 1062 32510 1114
rect 32510 1062 32540 1114
rect 32564 1062 32574 1114
rect 32574 1062 32620 1114
rect 32324 1060 32380 1062
rect 32404 1060 32460 1062
rect 32484 1060 32540 1062
rect 32564 1060 32620 1062
<< metal3 >>
rect 19977 21180 20043 21181
rect 23657 21180 23723 21181
rect 19926 21178 19932 21180
rect 19886 21118 19932 21178
rect 19996 21176 20043 21180
rect 23606 21178 23612 21180
rect 20038 21120 20043 21176
rect 19926 21116 19932 21118
rect 19996 21116 20043 21120
rect 23566 21118 23612 21178
rect 23676 21176 23723 21180
rect 23718 21120 23723 21176
rect 23606 21116 23612 21118
rect 23676 21116 23723 21120
rect 19977 21115 20043 21116
rect 23657 21115 23723 21116
rect 22185 21044 22251 21045
rect 22921 21044 22987 21045
rect 22134 21042 22140 21044
rect 22094 20982 22140 21042
rect 22204 21040 22251 21044
rect 22870 21042 22876 21044
rect 22246 20984 22251 21040
rect 22134 20980 22140 20982
rect 22204 20980 22251 20984
rect 22830 20982 22876 21042
rect 22940 21040 22987 21044
rect 22982 20984 22987 21040
rect 22870 20980 22876 20982
rect 22940 20980 22987 20984
rect 22185 20979 22251 20980
rect 22921 20979 22987 20980
rect 5257 20908 5323 20909
rect 5206 20844 5212 20908
rect 5276 20906 5323 20908
rect 5276 20904 5368 20906
rect 5318 20848 5368 20904
rect 5276 20846 5368 20848
rect 5276 20844 5323 20846
rect 8886 20844 8892 20908
rect 8956 20906 8962 20908
rect 9121 20906 9187 20909
rect 8956 20904 9187 20906
rect 8956 20848 9126 20904
rect 9182 20848 9187 20904
rect 8956 20846 9187 20848
rect 8956 20844 8962 20846
rect 5257 20843 5323 20844
rect 9121 20843 9187 20846
rect 16982 20844 16988 20908
rect 17052 20906 17058 20908
rect 17769 20906 17835 20909
rect 17052 20904 17835 20906
rect 17052 20848 17774 20904
rect 17830 20848 17835 20904
rect 17052 20846 17835 20848
rect 17052 20844 17058 20846
rect 17769 20843 17835 20846
rect 20662 20844 20668 20908
rect 20732 20906 20738 20908
rect 20897 20906 20963 20909
rect 20732 20904 20963 20906
rect 20732 20848 20902 20904
rect 20958 20848 20963 20904
rect 20732 20846 20963 20848
rect 20732 20844 20738 20846
rect 20897 20843 20963 20846
rect 17861 20770 17927 20773
rect 31753 20772 31819 20773
rect 19190 20770 19196 20772
rect 17861 20768 19196 20770
rect 17861 20712 17866 20768
rect 17922 20712 19196 20768
rect 17861 20710 19196 20712
rect 17861 20707 17927 20710
rect 19190 20708 19196 20710
rect 19260 20708 19266 20772
rect 31702 20770 31708 20772
rect 31662 20710 31708 20770
rect 31772 20768 31819 20772
rect 31814 20712 31819 20768
rect 31702 20708 31708 20710
rect 31772 20708 31819 20712
rect 31753 20707 31819 20708
rect 8788 20704 9104 20705
rect 8788 20640 8794 20704
rect 8858 20640 8874 20704
rect 8938 20640 8954 20704
rect 9018 20640 9034 20704
rect 9098 20640 9104 20704
rect 8788 20639 9104 20640
rect 16630 20704 16946 20705
rect 16630 20640 16636 20704
rect 16700 20640 16716 20704
rect 16780 20640 16796 20704
rect 16860 20640 16876 20704
rect 16940 20640 16946 20704
rect 16630 20639 16946 20640
rect 24472 20704 24788 20705
rect 24472 20640 24478 20704
rect 24542 20640 24558 20704
rect 24622 20640 24638 20704
rect 24702 20640 24718 20704
rect 24782 20640 24788 20704
rect 24472 20639 24788 20640
rect 32314 20704 32630 20705
rect 32314 20640 32320 20704
rect 32384 20640 32400 20704
rect 32464 20640 32480 20704
rect 32544 20640 32560 20704
rect 32624 20640 32630 20704
rect 32314 20639 32630 20640
rect 11094 20572 11100 20636
rect 11164 20634 11170 20636
rect 11973 20634 12039 20637
rect 11164 20632 12039 20634
rect 11164 20576 11978 20632
rect 12034 20576 12039 20632
rect 11164 20574 12039 20576
rect 11164 20572 11170 20574
rect 11973 20571 12039 20574
rect 12566 20572 12572 20636
rect 12636 20634 12642 20636
rect 12709 20634 12775 20637
rect 14825 20636 14891 20637
rect 12636 20632 12775 20634
rect 12636 20576 12714 20632
rect 12770 20576 12775 20632
rect 12636 20574 12775 20576
rect 12636 20572 12642 20574
rect 12709 20571 12775 20574
rect 14774 20572 14780 20636
rect 14844 20634 14891 20636
rect 14844 20632 14936 20634
rect 14886 20576 14936 20632
rect 14844 20574 14936 20576
rect 14844 20572 14891 20574
rect 18454 20572 18460 20636
rect 18524 20634 18530 20636
rect 18689 20634 18755 20637
rect 18524 20632 18755 20634
rect 18524 20576 18694 20632
rect 18750 20576 18755 20632
rect 18524 20574 18755 20576
rect 18524 20572 18530 20574
rect 14825 20571 14891 20572
rect 18689 20571 18755 20574
rect 8150 20436 8156 20500
rect 8220 20498 8226 20500
rect 11053 20498 11119 20501
rect 21449 20500 21515 20501
rect 21398 20498 21404 20500
rect 8220 20496 11119 20498
rect 8220 20440 11058 20496
rect 11114 20440 11119 20496
rect 8220 20438 11119 20440
rect 21358 20438 21404 20498
rect 21468 20496 21515 20500
rect 21510 20440 21515 20496
rect 8220 20436 8226 20438
rect 11053 20435 11119 20438
rect 21398 20436 21404 20438
rect 21468 20436 21515 20440
rect 21449 20435 21515 20436
rect 4867 20160 5183 20161
rect 4867 20096 4873 20160
rect 4937 20096 4953 20160
rect 5017 20096 5033 20160
rect 5097 20096 5113 20160
rect 5177 20096 5183 20160
rect 4867 20095 5183 20096
rect 12709 20160 13025 20161
rect 12709 20096 12715 20160
rect 12779 20096 12795 20160
rect 12859 20096 12875 20160
rect 12939 20096 12955 20160
rect 13019 20096 13025 20160
rect 12709 20095 13025 20096
rect 20551 20160 20867 20161
rect 20551 20096 20557 20160
rect 20621 20096 20637 20160
rect 20701 20096 20717 20160
rect 20781 20096 20797 20160
rect 20861 20096 20867 20160
rect 20551 20095 20867 20096
rect 28393 20160 28709 20161
rect 28393 20096 28399 20160
rect 28463 20096 28479 20160
rect 28543 20096 28559 20160
rect 28623 20096 28639 20160
rect 28703 20096 28709 20160
rect 28393 20095 28709 20096
rect 2221 20092 2287 20093
rect 3049 20092 3115 20093
rect 2221 20090 2268 20092
rect 2176 20088 2268 20090
rect 2176 20032 2226 20088
rect 2176 20030 2268 20032
rect 2221 20028 2268 20030
rect 2332 20028 2338 20092
rect 2998 20028 3004 20092
rect 3068 20090 3115 20092
rect 4337 20090 4403 20093
rect 4470 20090 4476 20092
rect 3068 20088 3160 20090
rect 3110 20032 3160 20088
rect 3068 20030 3160 20032
rect 4337 20088 4476 20090
rect 4337 20032 4342 20088
rect 4398 20032 4476 20088
rect 4337 20030 4476 20032
rect 3068 20028 3115 20030
rect 2221 20027 2287 20028
rect 3049 20027 3115 20028
rect 4337 20027 4403 20030
rect 4470 20028 4476 20030
rect 4540 20028 4546 20092
rect 5809 20090 5875 20093
rect 5942 20090 5948 20092
rect 5809 20088 5948 20090
rect 5809 20032 5814 20088
rect 5870 20032 5948 20088
rect 5809 20030 5948 20032
rect 5809 20027 5875 20030
rect 5942 20028 5948 20030
rect 6012 20028 6018 20092
rect 6545 20090 6611 20093
rect 6678 20090 6684 20092
rect 6545 20088 6684 20090
rect 6545 20032 6550 20088
rect 6606 20032 6684 20088
rect 6545 20030 6684 20032
rect 6545 20027 6611 20030
rect 6678 20028 6684 20030
rect 6748 20028 6754 20092
rect 13721 20090 13787 20093
rect 14038 20090 14044 20092
rect 13721 20088 14044 20090
rect 13721 20032 13726 20088
rect 13782 20032 14044 20088
rect 13721 20030 14044 20032
rect 13721 20027 13787 20030
rect 14038 20028 14044 20030
rect 14108 20028 14114 20092
rect 7414 19892 7420 19956
rect 7484 19954 7490 19956
rect 11053 19954 11119 19957
rect 7484 19952 11119 19954
rect 7484 19896 11058 19952
rect 11114 19896 11119 19952
rect 7484 19894 11119 19896
rect 7484 19892 7490 19894
rect 11053 19891 11119 19894
rect 30966 19620 30972 19684
rect 31036 19682 31042 19684
rect 31293 19682 31359 19685
rect 31036 19680 31359 19682
rect 31036 19624 31298 19680
rect 31354 19624 31359 19680
rect 31036 19622 31359 19624
rect 31036 19620 31042 19622
rect 31293 19619 31359 19622
rect 8788 19616 9104 19617
rect 8788 19552 8794 19616
rect 8858 19552 8874 19616
rect 8938 19552 8954 19616
rect 9018 19552 9034 19616
rect 9098 19552 9104 19616
rect 8788 19551 9104 19552
rect 16630 19616 16946 19617
rect 16630 19552 16636 19616
rect 16700 19552 16716 19616
rect 16780 19552 16796 19616
rect 16860 19552 16876 19616
rect 16940 19552 16946 19616
rect 16630 19551 16946 19552
rect 24472 19616 24788 19617
rect 24472 19552 24478 19616
rect 24542 19552 24558 19616
rect 24622 19552 24638 19616
rect 24702 19552 24718 19616
rect 24782 19552 24788 19616
rect 24472 19551 24788 19552
rect 32314 19616 32630 19617
rect 32314 19552 32320 19616
rect 32384 19552 32400 19616
rect 32464 19552 32480 19616
rect 32544 19552 32560 19616
rect 32624 19552 32630 19616
rect 32314 19551 32630 19552
rect 1526 19484 1532 19548
rect 1596 19546 1602 19548
rect 2405 19546 2471 19549
rect 1596 19544 2471 19546
rect 1596 19488 2410 19544
rect 2466 19488 2471 19544
rect 1596 19486 2471 19488
rect 1596 19484 1602 19486
rect 2405 19483 2471 19486
rect 3734 19484 3740 19548
rect 3804 19546 3810 19548
rect 3877 19546 3943 19549
rect 3804 19544 3943 19546
rect 3804 19488 3882 19544
rect 3938 19488 3943 19544
rect 3804 19486 3943 19488
rect 3804 19484 3810 19486
rect 3877 19483 3943 19486
rect 9622 19484 9628 19548
rect 9692 19546 9698 19548
rect 10961 19546 11027 19549
rect 11881 19548 11947 19549
rect 9692 19544 11027 19546
rect 9692 19488 10966 19544
rect 11022 19488 11027 19544
rect 9692 19486 11027 19488
rect 9692 19484 9698 19486
rect 10961 19483 11027 19486
rect 11830 19484 11836 19548
rect 11900 19546 11947 19548
rect 16113 19546 16179 19549
rect 16246 19546 16252 19548
rect 11900 19544 11992 19546
rect 11942 19488 11992 19544
rect 11900 19486 11992 19488
rect 16113 19544 16252 19546
rect 16113 19488 16118 19544
rect 16174 19488 16252 19544
rect 16113 19486 16252 19488
rect 11900 19484 11947 19486
rect 11881 19483 11947 19484
rect 16113 19483 16179 19486
rect 16246 19484 16252 19486
rect 16316 19484 16322 19548
rect 17769 19412 17835 19413
rect 17718 19348 17724 19412
rect 17788 19410 17835 19412
rect 17788 19408 17880 19410
rect 17830 19352 17880 19408
rect 17788 19350 17880 19352
rect 17788 19348 17835 19350
rect 17769 19347 17835 19348
rect 13302 19212 13308 19276
rect 13372 19274 13378 19276
rect 13813 19274 13879 19277
rect 13372 19272 13879 19274
rect 13372 19216 13818 19272
rect 13874 19216 13879 19272
rect 13372 19214 13879 19216
rect 13372 19212 13378 19214
rect 13813 19211 13879 19214
rect 24158 19212 24164 19276
rect 24228 19274 24234 19276
rect 24853 19274 24919 19277
rect 24228 19272 24919 19274
rect 24228 19216 24858 19272
rect 24914 19216 24919 19272
rect 24228 19214 24919 19216
rect 24228 19212 24234 19214
rect 24853 19211 24919 19214
rect 4867 19072 5183 19073
rect 4867 19008 4873 19072
rect 4937 19008 4953 19072
rect 5017 19008 5033 19072
rect 5097 19008 5113 19072
rect 5177 19008 5183 19072
rect 4867 19007 5183 19008
rect 12709 19072 13025 19073
rect 12709 19008 12715 19072
rect 12779 19008 12795 19072
rect 12859 19008 12875 19072
rect 12939 19008 12955 19072
rect 13019 19008 13025 19072
rect 12709 19007 13025 19008
rect 20551 19072 20867 19073
rect 20551 19008 20557 19072
rect 20621 19008 20637 19072
rect 20701 19008 20717 19072
rect 20781 19008 20797 19072
rect 20861 19008 20867 19072
rect 20551 19007 20867 19008
rect 28393 19072 28709 19073
rect 28393 19008 28399 19072
rect 28463 19008 28479 19072
rect 28543 19008 28559 19072
rect 28623 19008 28639 19072
rect 28703 19008 28709 19072
rect 28393 19007 28709 19008
rect 10358 18940 10364 19004
rect 10428 19002 10434 19004
rect 11053 19002 11119 19005
rect 10428 19000 11119 19002
rect 10428 18944 11058 19000
rect 11114 18944 11119 19000
rect 10428 18942 11119 18944
rect 10428 18940 10434 18942
rect 11053 18939 11119 18942
rect 15510 18940 15516 19004
rect 15580 19002 15586 19004
rect 16573 19002 16639 19005
rect 15580 19000 16639 19002
rect 15580 18944 16578 19000
rect 16634 18944 16639 19000
rect 15580 18942 16639 18944
rect 15580 18940 15586 18942
rect 16573 18939 16639 18942
rect 8788 18528 9104 18529
rect 8788 18464 8794 18528
rect 8858 18464 8874 18528
rect 8938 18464 8954 18528
rect 9018 18464 9034 18528
rect 9098 18464 9104 18528
rect 8788 18463 9104 18464
rect 16630 18528 16946 18529
rect 16630 18464 16636 18528
rect 16700 18464 16716 18528
rect 16780 18464 16796 18528
rect 16860 18464 16876 18528
rect 16940 18464 16946 18528
rect 16630 18463 16946 18464
rect 24472 18528 24788 18529
rect 24472 18464 24478 18528
rect 24542 18464 24558 18528
rect 24622 18464 24638 18528
rect 24702 18464 24718 18528
rect 24782 18464 24788 18528
rect 24472 18463 24788 18464
rect 32314 18528 32630 18529
rect 32314 18464 32320 18528
rect 32384 18464 32400 18528
rect 32464 18464 32480 18528
rect 32544 18464 32560 18528
rect 32624 18464 32630 18528
rect 32314 18463 32630 18464
rect 4867 17984 5183 17985
rect 4867 17920 4873 17984
rect 4937 17920 4953 17984
rect 5017 17920 5033 17984
rect 5097 17920 5113 17984
rect 5177 17920 5183 17984
rect 4867 17919 5183 17920
rect 12709 17984 13025 17985
rect 12709 17920 12715 17984
rect 12779 17920 12795 17984
rect 12859 17920 12875 17984
rect 12939 17920 12955 17984
rect 13019 17920 13025 17984
rect 12709 17919 13025 17920
rect 20551 17984 20867 17985
rect 20551 17920 20557 17984
rect 20621 17920 20637 17984
rect 20701 17920 20717 17984
rect 20781 17920 20797 17984
rect 20861 17920 20867 17984
rect 20551 17919 20867 17920
rect 28393 17984 28709 17985
rect 28393 17920 28399 17984
rect 28463 17920 28479 17984
rect 28543 17920 28559 17984
rect 28623 17920 28639 17984
rect 28703 17920 28709 17984
rect 28393 17919 28709 17920
rect 30281 17916 30347 17917
rect 30230 17914 30236 17916
rect 30190 17854 30236 17914
rect 30300 17912 30347 17916
rect 30342 17856 30347 17912
rect 30230 17852 30236 17854
rect 30300 17852 30347 17856
rect 30281 17851 30347 17852
rect 8788 17440 9104 17441
rect 8788 17376 8794 17440
rect 8858 17376 8874 17440
rect 8938 17376 8954 17440
rect 9018 17376 9034 17440
rect 9098 17376 9104 17440
rect 8788 17375 9104 17376
rect 16630 17440 16946 17441
rect 16630 17376 16636 17440
rect 16700 17376 16716 17440
rect 16780 17376 16796 17440
rect 16860 17376 16876 17440
rect 16940 17376 16946 17440
rect 16630 17375 16946 17376
rect 24472 17440 24788 17441
rect 24472 17376 24478 17440
rect 24542 17376 24558 17440
rect 24622 17376 24638 17440
rect 24702 17376 24718 17440
rect 24782 17376 24788 17440
rect 24472 17375 24788 17376
rect 32314 17440 32630 17441
rect 32314 17376 32320 17440
rect 32384 17376 32400 17440
rect 32464 17376 32480 17440
rect 32544 17376 32560 17440
rect 32624 17376 32630 17440
rect 32314 17375 32630 17376
rect 4867 16896 5183 16897
rect 4867 16832 4873 16896
rect 4937 16832 4953 16896
rect 5017 16832 5033 16896
rect 5097 16832 5113 16896
rect 5177 16832 5183 16896
rect 4867 16831 5183 16832
rect 12709 16896 13025 16897
rect 12709 16832 12715 16896
rect 12779 16832 12795 16896
rect 12859 16832 12875 16896
rect 12939 16832 12955 16896
rect 13019 16832 13025 16896
rect 12709 16831 13025 16832
rect 20551 16896 20867 16897
rect 20551 16832 20557 16896
rect 20621 16832 20637 16896
rect 20701 16832 20717 16896
rect 20781 16832 20797 16896
rect 20861 16832 20867 16896
rect 20551 16831 20867 16832
rect 28393 16896 28709 16897
rect 28393 16832 28399 16896
rect 28463 16832 28479 16896
rect 28543 16832 28559 16896
rect 28623 16832 28639 16896
rect 28703 16832 28709 16896
rect 28393 16831 28709 16832
rect 8788 16352 9104 16353
rect 8788 16288 8794 16352
rect 8858 16288 8874 16352
rect 8938 16288 8954 16352
rect 9018 16288 9034 16352
rect 9098 16288 9104 16352
rect 8788 16287 9104 16288
rect 16630 16352 16946 16353
rect 16630 16288 16636 16352
rect 16700 16288 16716 16352
rect 16780 16288 16796 16352
rect 16860 16288 16876 16352
rect 16940 16288 16946 16352
rect 16630 16287 16946 16288
rect 24472 16352 24788 16353
rect 24472 16288 24478 16352
rect 24542 16288 24558 16352
rect 24622 16288 24638 16352
rect 24702 16288 24718 16352
rect 24782 16288 24788 16352
rect 24472 16287 24788 16288
rect 32314 16352 32630 16353
rect 32314 16288 32320 16352
rect 32384 16288 32400 16352
rect 32464 16288 32480 16352
rect 32544 16288 32560 16352
rect 32624 16288 32630 16352
rect 32314 16287 32630 16288
rect 4867 15808 5183 15809
rect 4867 15744 4873 15808
rect 4937 15744 4953 15808
rect 5017 15744 5033 15808
rect 5097 15744 5113 15808
rect 5177 15744 5183 15808
rect 4867 15743 5183 15744
rect 12709 15808 13025 15809
rect 12709 15744 12715 15808
rect 12779 15744 12795 15808
rect 12859 15744 12875 15808
rect 12939 15744 12955 15808
rect 13019 15744 13025 15808
rect 12709 15743 13025 15744
rect 20551 15808 20867 15809
rect 20551 15744 20557 15808
rect 20621 15744 20637 15808
rect 20701 15744 20717 15808
rect 20781 15744 20797 15808
rect 20861 15744 20867 15808
rect 20551 15743 20867 15744
rect 28393 15808 28709 15809
rect 28393 15744 28399 15808
rect 28463 15744 28479 15808
rect 28543 15744 28559 15808
rect 28623 15744 28639 15808
rect 28703 15744 28709 15808
rect 28393 15743 28709 15744
rect 8788 15264 9104 15265
rect 8788 15200 8794 15264
rect 8858 15200 8874 15264
rect 8938 15200 8954 15264
rect 9018 15200 9034 15264
rect 9098 15200 9104 15264
rect 8788 15199 9104 15200
rect 16630 15264 16946 15265
rect 16630 15200 16636 15264
rect 16700 15200 16716 15264
rect 16780 15200 16796 15264
rect 16860 15200 16876 15264
rect 16940 15200 16946 15264
rect 16630 15199 16946 15200
rect 24472 15264 24788 15265
rect 24472 15200 24478 15264
rect 24542 15200 24558 15264
rect 24622 15200 24638 15264
rect 24702 15200 24718 15264
rect 24782 15200 24788 15264
rect 24472 15199 24788 15200
rect 32314 15264 32630 15265
rect 32314 15200 32320 15264
rect 32384 15200 32400 15264
rect 32464 15200 32480 15264
rect 32544 15200 32560 15264
rect 32624 15200 32630 15264
rect 32314 15199 32630 15200
rect 4867 14720 5183 14721
rect 4867 14656 4873 14720
rect 4937 14656 4953 14720
rect 5017 14656 5033 14720
rect 5097 14656 5113 14720
rect 5177 14656 5183 14720
rect 4867 14655 5183 14656
rect 12709 14720 13025 14721
rect 12709 14656 12715 14720
rect 12779 14656 12795 14720
rect 12859 14656 12875 14720
rect 12939 14656 12955 14720
rect 13019 14656 13025 14720
rect 12709 14655 13025 14656
rect 20551 14720 20867 14721
rect 20551 14656 20557 14720
rect 20621 14656 20637 14720
rect 20701 14656 20717 14720
rect 20781 14656 20797 14720
rect 20861 14656 20867 14720
rect 20551 14655 20867 14656
rect 28393 14720 28709 14721
rect 28393 14656 28399 14720
rect 28463 14656 28479 14720
rect 28543 14656 28559 14720
rect 28623 14656 28639 14720
rect 28703 14656 28709 14720
rect 28393 14655 28709 14656
rect 8788 14176 9104 14177
rect 8788 14112 8794 14176
rect 8858 14112 8874 14176
rect 8938 14112 8954 14176
rect 9018 14112 9034 14176
rect 9098 14112 9104 14176
rect 8788 14111 9104 14112
rect 16630 14176 16946 14177
rect 16630 14112 16636 14176
rect 16700 14112 16716 14176
rect 16780 14112 16796 14176
rect 16860 14112 16876 14176
rect 16940 14112 16946 14176
rect 16630 14111 16946 14112
rect 24472 14176 24788 14177
rect 24472 14112 24478 14176
rect 24542 14112 24558 14176
rect 24622 14112 24638 14176
rect 24702 14112 24718 14176
rect 24782 14112 24788 14176
rect 24472 14111 24788 14112
rect 32314 14176 32630 14177
rect 32314 14112 32320 14176
rect 32384 14112 32400 14176
rect 32464 14112 32480 14176
rect 32544 14112 32560 14176
rect 32624 14112 32630 14176
rect 32314 14111 32630 14112
rect 4867 13632 5183 13633
rect 4867 13568 4873 13632
rect 4937 13568 4953 13632
rect 5017 13568 5033 13632
rect 5097 13568 5113 13632
rect 5177 13568 5183 13632
rect 4867 13567 5183 13568
rect 12709 13632 13025 13633
rect 12709 13568 12715 13632
rect 12779 13568 12795 13632
rect 12859 13568 12875 13632
rect 12939 13568 12955 13632
rect 13019 13568 13025 13632
rect 12709 13567 13025 13568
rect 20551 13632 20867 13633
rect 20551 13568 20557 13632
rect 20621 13568 20637 13632
rect 20701 13568 20717 13632
rect 20781 13568 20797 13632
rect 20861 13568 20867 13632
rect 20551 13567 20867 13568
rect 28393 13632 28709 13633
rect 28393 13568 28399 13632
rect 28463 13568 28479 13632
rect 28543 13568 28559 13632
rect 28623 13568 28639 13632
rect 28703 13568 28709 13632
rect 28393 13567 28709 13568
rect 8788 13088 9104 13089
rect 8788 13024 8794 13088
rect 8858 13024 8874 13088
rect 8938 13024 8954 13088
rect 9018 13024 9034 13088
rect 9098 13024 9104 13088
rect 8788 13023 9104 13024
rect 16630 13088 16946 13089
rect 16630 13024 16636 13088
rect 16700 13024 16716 13088
rect 16780 13024 16796 13088
rect 16860 13024 16876 13088
rect 16940 13024 16946 13088
rect 16630 13023 16946 13024
rect 24472 13088 24788 13089
rect 24472 13024 24478 13088
rect 24542 13024 24558 13088
rect 24622 13024 24638 13088
rect 24702 13024 24718 13088
rect 24782 13024 24788 13088
rect 24472 13023 24788 13024
rect 32314 13088 32630 13089
rect 32314 13024 32320 13088
rect 32384 13024 32400 13088
rect 32464 13024 32480 13088
rect 32544 13024 32560 13088
rect 32624 13024 32630 13088
rect 32314 13023 32630 13024
rect 4867 12544 5183 12545
rect 4867 12480 4873 12544
rect 4937 12480 4953 12544
rect 5017 12480 5033 12544
rect 5097 12480 5113 12544
rect 5177 12480 5183 12544
rect 4867 12479 5183 12480
rect 12709 12544 13025 12545
rect 12709 12480 12715 12544
rect 12779 12480 12795 12544
rect 12859 12480 12875 12544
rect 12939 12480 12955 12544
rect 13019 12480 13025 12544
rect 12709 12479 13025 12480
rect 20551 12544 20867 12545
rect 20551 12480 20557 12544
rect 20621 12480 20637 12544
rect 20701 12480 20717 12544
rect 20781 12480 20797 12544
rect 20861 12480 20867 12544
rect 20551 12479 20867 12480
rect 28393 12544 28709 12545
rect 28393 12480 28399 12544
rect 28463 12480 28479 12544
rect 28543 12480 28559 12544
rect 28623 12480 28639 12544
rect 28703 12480 28709 12544
rect 28393 12479 28709 12480
rect 8788 12000 9104 12001
rect 8788 11936 8794 12000
rect 8858 11936 8874 12000
rect 8938 11936 8954 12000
rect 9018 11936 9034 12000
rect 9098 11936 9104 12000
rect 8788 11935 9104 11936
rect 16630 12000 16946 12001
rect 16630 11936 16636 12000
rect 16700 11936 16716 12000
rect 16780 11936 16796 12000
rect 16860 11936 16876 12000
rect 16940 11936 16946 12000
rect 16630 11935 16946 11936
rect 24472 12000 24788 12001
rect 24472 11936 24478 12000
rect 24542 11936 24558 12000
rect 24622 11936 24638 12000
rect 24702 11936 24718 12000
rect 24782 11936 24788 12000
rect 24472 11935 24788 11936
rect 32314 12000 32630 12001
rect 32314 11936 32320 12000
rect 32384 11936 32400 12000
rect 32464 11936 32480 12000
rect 32544 11936 32560 12000
rect 32624 11936 32630 12000
rect 32314 11935 32630 11936
rect 4867 11456 5183 11457
rect 4867 11392 4873 11456
rect 4937 11392 4953 11456
rect 5017 11392 5033 11456
rect 5097 11392 5113 11456
rect 5177 11392 5183 11456
rect 4867 11391 5183 11392
rect 12709 11456 13025 11457
rect 12709 11392 12715 11456
rect 12779 11392 12795 11456
rect 12859 11392 12875 11456
rect 12939 11392 12955 11456
rect 13019 11392 13025 11456
rect 12709 11391 13025 11392
rect 20551 11456 20867 11457
rect 20551 11392 20557 11456
rect 20621 11392 20637 11456
rect 20701 11392 20717 11456
rect 20781 11392 20797 11456
rect 20861 11392 20867 11456
rect 20551 11391 20867 11392
rect 28393 11456 28709 11457
rect 28393 11392 28399 11456
rect 28463 11392 28479 11456
rect 28543 11392 28559 11456
rect 28623 11392 28639 11456
rect 28703 11392 28709 11456
rect 28393 11391 28709 11392
rect 8788 10912 9104 10913
rect 8788 10848 8794 10912
rect 8858 10848 8874 10912
rect 8938 10848 8954 10912
rect 9018 10848 9034 10912
rect 9098 10848 9104 10912
rect 8788 10847 9104 10848
rect 16630 10912 16946 10913
rect 16630 10848 16636 10912
rect 16700 10848 16716 10912
rect 16780 10848 16796 10912
rect 16860 10848 16876 10912
rect 16940 10848 16946 10912
rect 16630 10847 16946 10848
rect 24472 10912 24788 10913
rect 24472 10848 24478 10912
rect 24542 10848 24558 10912
rect 24622 10848 24638 10912
rect 24702 10848 24718 10912
rect 24782 10848 24788 10912
rect 24472 10847 24788 10848
rect 32314 10912 32630 10913
rect 32314 10848 32320 10912
rect 32384 10848 32400 10912
rect 32464 10848 32480 10912
rect 32544 10848 32560 10912
rect 32624 10848 32630 10912
rect 32314 10847 32630 10848
rect 4867 10368 5183 10369
rect 4867 10304 4873 10368
rect 4937 10304 4953 10368
rect 5017 10304 5033 10368
rect 5097 10304 5113 10368
rect 5177 10304 5183 10368
rect 4867 10303 5183 10304
rect 12709 10368 13025 10369
rect 12709 10304 12715 10368
rect 12779 10304 12795 10368
rect 12859 10304 12875 10368
rect 12939 10304 12955 10368
rect 13019 10304 13025 10368
rect 12709 10303 13025 10304
rect 20551 10368 20867 10369
rect 20551 10304 20557 10368
rect 20621 10304 20637 10368
rect 20701 10304 20717 10368
rect 20781 10304 20797 10368
rect 20861 10304 20867 10368
rect 20551 10303 20867 10304
rect 28393 10368 28709 10369
rect 28393 10304 28399 10368
rect 28463 10304 28479 10368
rect 28543 10304 28559 10368
rect 28623 10304 28639 10368
rect 28703 10304 28709 10368
rect 28393 10303 28709 10304
rect 8788 9824 9104 9825
rect 8788 9760 8794 9824
rect 8858 9760 8874 9824
rect 8938 9760 8954 9824
rect 9018 9760 9034 9824
rect 9098 9760 9104 9824
rect 8788 9759 9104 9760
rect 16630 9824 16946 9825
rect 16630 9760 16636 9824
rect 16700 9760 16716 9824
rect 16780 9760 16796 9824
rect 16860 9760 16876 9824
rect 16940 9760 16946 9824
rect 16630 9759 16946 9760
rect 24472 9824 24788 9825
rect 24472 9760 24478 9824
rect 24542 9760 24558 9824
rect 24622 9760 24638 9824
rect 24702 9760 24718 9824
rect 24782 9760 24788 9824
rect 24472 9759 24788 9760
rect 32314 9824 32630 9825
rect 32314 9760 32320 9824
rect 32384 9760 32400 9824
rect 32464 9760 32480 9824
rect 32544 9760 32560 9824
rect 32624 9760 32630 9824
rect 32314 9759 32630 9760
rect 4867 9280 5183 9281
rect 4867 9216 4873 9280
rect 4937 9216 4953 9280
rect 5017 9216 5033 9280
rect 5097 9216 5113 9280
rect 5177 9216 5183 9280
rect 4867 9215 5183 9216
rect 12709 9280 13025 9281
rect 12709 9216 12715 9280
rect 12779 9216 12795 9280
rect 12859 9216 12875 9280
rect 12939 9216 12955 9280
rect 13019 9216 13025 9280
rect 12709 9215 13025 9216
rect 20551 9280 20867 9281
rect 20551 9216 20557 9280
rect 20621 9216 20637 9280
rect 20701 9216 20717 9280
rect 20781 9216 20797 9280
rect 20861 9216 20867 9280
rect 20551 9215 20867 9216
rect 28393 9280 28709 9281
rect 28393 9216 28399 9280
rect 28463 9216 28479 9280
rect 28543 9216 28559 9280
rect 28623 9216 28639 9280
rect 28703 9216 28709 9280
rect 28393 9215 28709 9216
rect 8788 8736 9104 8737
rect 8788 8672 8794 8736
rect 8858 8672 8874 8736
rect 8938 8672 8954 8736
rect 9018 8672 9034 8736
rect 9098 8672 9104 8736
rect 8788 8671 9104 8672
rect 16630 8736 16946 8737
rect 16630 8672 16636 8736
rect 16700 8672 16716 8736
rect 16780 8672 16796 8736
rect 16860 8672 16876 8736
rect 16940 8672 16946 8736
rect 16630 8671 16946 8672
rect 24472 8736 24788 8737
rect 24472 8672 24478 8736
rect 24542 8672 24558 8736
rect 24622 8672 24638 8736
rect 24702 8672 24718 8736
rect 24782 8672 24788 8736
rect 24472 8671 24788 8672
rect 32314 8736 32630 8737
rect 32314 8672 32320 8736
rect 32384 8672 32400 8736
rect 32464 8672 32480 8736
rect 32544 8672 32560 8736
rect 32624 8672 32630 8736
rect 32314 8671 32630 8672
rect 4867 8192 5183 8193
rect 4867 8128 4873 8192
rect 4937 8128 4953 8192
rect 5017 8128 5033 8192
rect 5097 8128 5113 8192
rect 5177 8128 5183 8192
rect 4867 8127 5183 8128
rect 12709 8192 13025 8193
rect 12709 8128 12715 8192
rect 12779 8128 12795 8192
rect 12859 8128 12875 8192
rect 12939 8128 12955 8192
rect 13019 8128 13025 8192
rect 12709 8127 13025 8128
rect 20551 8192 20867 8193
rect 20551 8128 20557 8192
rect 20621 8128 20637 8192
rect 20701 8128 20717 8192
rect 20781 8128 20797 8192
rect 20861 8128 20867 8192
rect 20551 8127 20867 8128
rect 28393 8192 28709 8193
rect 28393 8128 28399 8192
rect 28463 8128 28479 8192
rect 28543 8128 28559 8192
rect 28623 8128 28639 8192
rect 28703 8128 28709 8192
rect 28393 8127 28709 8128
rect 8788 7648 9104 7649
rect 8788 7584 8794 7648
rect 8858 7584 8874 7648
rect 8938 7584 8954 7648
rect 9018 7584 9034 7648
rect 9098 7584 9104 7648
rect 8788 7583 9104 7584
rect 16630 7648 16946 7649
rect 16630 7584 16636 7648
rect 16700 7584 16716 7648
rect 16780 7584 16796 7648
rect 16860 7584 16876 7648
rect 16940 7584 16946 7648
rect 16630 7583 16946 7584
rect 24472 7648 24788 7649
rect 24472 7584 24478 7648
rect 24542 7584 24558 7648
rect 24622 7584 24638 7648
rect 24702 7584 24718 7648
rect 24782 7584 24788 7648
rect 24472 7583 24788 7584
rect 32314 7648 32630 7649
rect 32314 7584 32320 7648
rect 32384 7584 32400 7648
rect 32464 7584 32480 7648
rect 32544 7584 32560 7648
rect 32624 7584 32630 7648
rect 32314 7583 32630 7584
rect 4867 7104 5183 7105
rect 4867 7040 4873 7104
rect 4937 7040 4953 7104
rect 5017 7040 5033 7104
rect 5097 7040 5113 7104
rect 5177 7040 5183 7104
rect 4867 7039 5183 7040
rect 12709 7104 13025 7105
rect 12709 7040 12715 7104
rect 12779 7040 12795 7104
rect 12859 7040 12875 7104
rect 12939 7040 12955 7104
rect 13019 7040 13025 7104
rect 12709 7039 13025 7040
rect 20551 7104 20867 7105
rect 20551 7040 20557 7104
rect 20621 7040 20637 7104
rect 20701 7040 20717 7104
rect 20781 7040 20797 7104
rect 20861 7040 20867 7104
rect 20551 7039 20867 7040
rect 28393 7104 28709 7105
rect 28393 7040 28399 7104
rect 28463 7040 28479 7104
rect 28543 7040 28559 7104
rect 28623 7040 28639 7104
rect 28703 7040 28709 7104
rect 28393 7039 28709 7040
rect 8788 6560 9104 6561
rect 8788 6496 8794 6560
rect 8858 6496 8874 6560
rect 8938 6496 8954 6560
rect 9018 6496 9034 6560
rect 9098 6496 9104 6560
rect 8788 6495 9104 6496
rect 16630 6560 16946 6561
rect 16630 6496 16636 6560
rect 16700 6496 16716 6560
rect 16780 6496 16796 6560
rect 16860 6496 16876 6560
rect 16940 6496 16946 6560
rect 16630 6495 16946 6496
rect 24472 6560 24788 6561
rect 24472 6496 24478 6560
rect 24542 6496 24558 6560
rect 24622 6496 24638 6560
rect 24702 6496 24718 6560
rect 24782 6496 24788 6560
rect 24472 6495 24788 6496
rect 32314 6560 32630 6561
rect 32314 6496 32320 6560
rect 32384 6496 32400 6560
rect 32464 6496 32480 6560
rect 32544 6496 32560 6560
rect 32624 6496 32630 6560
rect 32314 6495 32630 6496
rect 4867 6016 5183 6017
rect 4867 5952 4873 6016
rect 4937 5952 4953 6016
rect 5017 5952 5033 6016
rect 5097 5952 5113 6016
rect 5177 5952 5183 6016
rect 4867 5951 5183 5952
rect 12709 6016 13025 6017
rect 12709 5952 12715 6016
rect 12779 5952 12795 6016
rect 12859 5952 12875 6016
rect 12939 5952 12955 6016
rect 13019 5952 13025 6016
rect 12709 5951 13025 5952
rect 20551 6016 20867 6017
rect 20551 5952 20557 6016
rect 20621 5952 20637 6016
rect 20701 5952 20717 6016
rect 20781 5952 20797 6016
rect 20861 5952 20867 6016
rect 20551 5951 20867 5952
rect 28393 6016 28709 6017
rect 28393 5952 28399 6016
rect 28463 5952 28479 6016
rect 28543 5952 28559 6016
rect 28623 5952 28639 6016
rect 28703 5952 28709 6016
rect 28393 5951 28709 5952
rect 8788 5472 9104 5473
rect 8788 5408 8794 5472
rect 8858 5408 8874 5472
rect 8938 5408 8954 5472
rect 9018 5408 9034 5472
rect 9098 5408 9104 5472
rect 8788 5407 9104 5408
rect 16630 5472 16946 5473
rect 16630 5408 16636 5472
rect 16700 5408 16716 5472
rect 16780 5408 16796 5472
rect 16860 5408 16876 5472
rect 16940 5408 16946 5472
rect 16630 5407 16946 5408
rect 24472 5472 24788 5473
rect 24472 5408 24478 5472
rect 24542 5408 24558 5472
rect 24622 5408 24638 5472
rect 24702 5408 24718 5472
rect 24782 5408 24788 5472
rect 24472 5407 24788 5408
rect 32314 5472 32630 5473
rect 32314 5408 32320 5472
rect 32384 5408 32400 5472
rect 32464 5408 32480 5472
rect 32544 5408 32560 5472
rect 32624 5408 32630 5472
rect 32314 5407 32630 5408
rect 4867 4928 5183 4929
rect 4867 4864 4873 4928
rect 4937 4864 4953 4928
rect 5017 4864 5033 4928
rect 5097 4864 5113 4928
rect 5177 4864 5183 4928
rect 4867 4863 5183 4864
rect 12709 4928 13025 4929
rect 12709 4864 12715 4928
rect 12779 4864 12795 4928
rect 12859 4864 12875 4928
rect 12939 4864 12955 4928
rect 13019 4864 13025 4928
rect 12709 4863 13025 4864
rect 20551 4928 20867 4929
rect 20551 4864 20557 4928
rect 20621 4864 20637 4928
rect 20701 4864 20717 4928
rect 20781 4864 20797 4928
rect 20861 4864 20867 4928
rect 20551 4863 20867 4864
rect 28393 4928 28709 4929
rect 28393 4864 28399 4928
rect 28463 4864 28479 4928
rect 28543 4864 28559 4928
rect 28623 4864 28639 4928
rect 28703 4864 28709 4928
rect 28393 4863 28709 4864
rect 8788 4384 9104 4385
rect 8788 4320 8794 4384
rect 8858 4320 8874 4384
rect 8938 4320 8954 4384
rect 9018 4320 9034 4384
rect 9098 4320 9104 4384
rect 8788 4319 9104 4320
rect 16630 4384 16946 4385
rect 16630 4320 16636 4384
rect 16700 4320 16716 4384
rect 16780 4320 16796 4384
rect 16860 4320 16876 4384
rect 16940 4320 16946 4384
rect 16630 4319 16946 4320
rect 24472 4384 24788 4385
rect 24472 4320 24478 4384
rect 24542 4320 24558 4384
rect 24622 4320 24638 4384
rect 24702 4320 24718 4384
rect 24782 4320 24788 4384
rect 24472 4319 24788 4320
rect 32314 4384 32630 4385
rect 32314 4320 32320 4384
rect 32384 4320 32400 4384
rect 32464 4320 32480 4384
rect 32544 4320 32560 4384
rect 32624 4320 32630 4384
rect 32314 4319 32630 4320
rect 4867 3840 5183 3841
rect 4867 3776 4873 3840
rect 4937 3776 4953 3840
rect 5017 3776 5033 3840
rect 5097 3776 5113 3840
rect 5177 3776 5183 3840
rect 4867 3775 5183 3776
rect 12709 3840 13025 3841
rect 12709 3776 12715 3840
rect 12779 3776 12795 3840
rect 12859 3776 12875 3840
rect 12939 3776 12955 3840
rect 13019 3776 13025 3840
rect 12709 3775 13025 3776
rect 20551 3840 20867 3841
rect 20551 3776 20557 3840
rect 20621 3776 20637 3840
rect 20701 3776 20717 3840
rect 20781 3776 20797 3840
rect 20861 3776 20867 3840
rect 20551 3775 20867 3776
rect 28393 3840 28709 3841
rect 28393 3776 28399 3840
rect 28463 3776 28479 3840
rect 28543 3776 28559 3840
rect 28623 3776 28639 3840
rect 28703 3776 28709 3840
rect 28393 3775 28709 3776
rect 8788 3296 9104 3297
rect 8788 3232 8794 3296
rect 8858 3232 8874 3296
rect 8938 3232 8954 3296
rect 9018 3232 9034 3296
rect 9098 3232 9104 3296
rect 8788 3231 9104 3232
rect 16630 3296 16946 3297
rect 16630 3232 16636 3296
rect 16700 3232 16716 3296
rect 16780 3232 16796 3296
rect 16860 3232 16876 3296
rect 16940 3232 16946 3296
rect 16630 3231 16946 3232
rect 24472 3296 24788 3297
rect 24472 3232 24478 3296
rect 24542 3232 24558 3296
rect 24622 3232 24638 3296
rect 24702 3232 24718 3296
rect 24782 3232 24788 3296
rect 24472 3231 24788 3232
rect 32314 3296 32630 3297
rect 32314 3232 32320 3296
rect 32384 3232 32400 3296
rect 32464 3232 32480 3296
rect 32544 3232 32560 3296
rect 32624 3232 32630 3296
rect 32314 3231 32630 3232
rect 4867 2752 5183 2753
rect 4867 2688 4873 2752
rect 4937 2688 4953 2752
rect 5017 2688 5033 2752
rect 5097 2688 5113 2752
rect 5177 2688 5183 2752
rect 4867 2687 5183 2688
rect 12709 2752 13025 2753
rect 12709 2688 12715 2752
rect 12779 2688 12795 2752
rect 12859 2688 12875 2752
rect 12939 2688 12955 2752
rect 13019 2688 13025 2752
rect 12709 2687 13025 2688
rect 20551 2752 20867 2753
rect 20551 2688 20557 2752
rect 20621 2688 20637 2752
rect 20701 2688 20717 2752
rect 20781 2688 20797 2752
rect 20861 2688 20867 2752
rect 20551 2687 20867 2688
rect 28393 2752 28709 2753
rect 28393 2688 28399 2752
rect 28463 2688 28479 2752
rect 28543 2688 28559 2752
rect 28623 2688 28639 2752
rect 28703 2688 28709 2752
rect 28393 2687 28709 2688
rect 8788 2208 9104 2209
rect 8788 2144 8794 2208
rect 8858 2144 8874 2208
rect 8938 2144 8954 2208
rect 9018 2144 9034 2208
rect 9098 2144 9104 2208
rect 8788 2143 9104 2144
rect 16630 2208 16946 2209
rect 16630 2144 16636 2208
rect 16700 2144 16716 2208
rect 16780 2144 16796 2208
rect 16860 2144 16876 2208
rect 16940 2144 16946 2208
rect 16630 2143 16946 2144
rect 24472 2208 24788 2209
rect 24472 2144 24478 2208
rect 24542 2144 24558 2208
rect 24622 2144 24638 2208
rect 24702 2144 24718 2208
rect 24782 2144 24788 2208
rect 24472 2143 24788 2144
rect 32314 2208 32630 2209
rect 32314 2144 32320 2208
rect 32384 2144 32400 2208
rect 32464 2144 32480 2208
rect 32544 2144 32560 2208
rect 32624 2144 32630 2208
rect 32314 2143 32630 2144
rect 4867 1664 5183 1665
rect 4867 1600 4873 1664
rect 4937 1600 4953 1664
rect 5017 1600 5033 1664
rect 5097 1600 5113 1664
rect 5177 1600 5183 1664
rect 4867 1599 5183 1600
rect 12709 1664 13025 1665
rect 12709 1600 12715 1664
rect 12779 1600 12795 1664
rect 12859 1600 12875 1664
rect 12939 1600 12955 1664
rect 13019 1600 13025 1664
rect 12709 1599 13025 1600
rect 20551 1664 20867 1665
rect 20551 1600 20557 1664
rect 20621 1600 20637 1664
rect 20701 1600 20717 1664
rect 20781 1600 20797 1664
rect 20861 1600 20867 1664
rect 20551 1599 20867 1600
rect 28393 1664 28709 1665
rect 28393 1600 28399 1664
rect 28463 1600 28479 1664
rect 28543 1600 28559 1664
rect 28623 1600 28639 1664
rect 28703 1600 28709 1664
rect 28393 1599 28709 1600
rect 8788 1120 9104 1121
rect 8788 1056 8794 1120
rect 8858 1056 8874 1120
rect 8938 1056 8954 1120
rect 9018 1056 9034 1120
rect 9098 1056 9104 1120
rect 8788 1055 9104 1056
rect 16630 1120 16946 1121
rect 16630 1056 16636 1120
rect 16700 1056 16716 1120
rect 16780 1056 16796 1120
rect 16860 1056 16876 1120
rect 16940 1056 16946 1120
rect 16630 1055 16946 1056
rect 24472 1120 24788 1121
rect 24472 1056 24478 1120
rect 24542 1056 24558 1120
rect 24622 1056 24638 1120
rect 24702 1056 24718 1120
rect 24782 1056 24788 1120
rect 24472 1055 24788 1056
rect 32314 1120 32630 1121
rect 32314 1056 32320 1120
rect 32384 1056 32400 1120
rect 32464 1056 32480 1120
rect 32544 1056 32560 1120
rect 32624 1056 32630 1120
rect 32314 1055 32630 1056
<< via3 >>
rect 19932 21176 19996 21180
rect 19932 21120 19982 21176
rect 19982 21120 19996 21176
rect 19932 21116 19996 21120
rect 23612 21176 23676 21180
rect 23612 21120 23662 21176
rect 23662 21120 23676 21176
rect 23612 21116 23676 21120
rect 22140 21040 22204 21044
rect 22140 20984 22190 21040
rect 22190 20984 22204 21040
rect 22140 20980 22204 20984
rect 22876 21040 22940 21044
rect 22876 20984 22926 21040
rect 22926 20984 22940 21040
rect 22876 20980 22940 20984
rect 5212 20904 5276 20908
rect 5212 20848 5262 20904
rect 5262 20848 5276 20904
rect 5212 20844 5276 20848
rect 8892 20844 8956 20908
rect 16988 20844 17052 20908
rect 20668 20844 20732 20908
rect 19196 20708 19260 20772
rect 31708 20768 31772 20772
rect 31708 20712 31758 20768
rect 31758 20712 31772 20768
rect 31708 20708 31772 20712
rect 8794 20700 8858 20704
rect 8794 20644 8798 20700
rect 8798 20644 8854 20700
rect 8854 20644 8858 20700
rect 8794 20640 8858 20644
rect 8874 20700 8938 20704
rect 8874 20644 8878 20700
rect 8878 20644 8934 20700
rect 8934 20644 8938 20700
rect 8874 20640 8938 20644
rect 8954 20700 9018 20704
rect 8954 20644 8958 20700
rect 8958 20644 9014 20700
rect 9014 20644 9018 20700
rect 8954 20640 9018 20644
rect 9034 20700 9098 20704
rect 9034 20644 9038 20700
rect 9038 20644 9094 20700
rect 9094 20644 9098 20700
rect 9034 20640 9098 20644
rect 16636 20700 16700 20704
rect 16636 20644 16640 20700
rect 16640 20644 16696 20700
rect 16696 20644 16700 20700
rect 16636 20640 16700 20644
rect 16716 20700 16780 20704
rect 16716 20644 16720 20700
rect 16720 20644 16776 20700
rect 16776 20644 16780 20700
rect 16716 20640 16780 20644
rect 16796 20700 16860 20704
rect 16796 20644 16800 20700
rect 16800 20644 16856 20700
rect 16856 20644 16860 20700
rect 16796 20640 16860 20644
rect 16876 20700 16940 20704
rect 16876 20644 16880 20700
rect 16880 20644 16936 20700
rect 16936 20644 16940 20700
rect 16876 20640 16940 20644
rect 24478 20700 24542 20704
rect 24478 20644 24482 20700
rect 24482 20644 24538 20700
rect 24538 20644 24542 20700
rect 24478 20640 24542 20644
rect 24558 20700 24622 20704
rect 24558 20644 24562 20700
rect 24562 20644 24618 20700
rect 24618 20644 24622 20700
rect 24558 20640 24622 20644
rect 24638 20700 24702 20704
rect 24638 20644 24642 20700
rect 24642 20644 24698 20700
rect 24698 20644 24702 20700
rect 24638 20640 24702 20644
rect 24718 20700 24782 20704
rect 24718 20644 24722 20700
rect 24722 20644 24778 20700
rect 24778 20644 24782 20700
rect 24718 20640 24782 20644
rect 32320 20700 32384 20704
rect 32320 20644 32324 20700
rect 32324 20644 32380 20700
rect 32380 20644 32384 20700
rect 32320 20640 32384 20644
rect 32400 20700 32464 20704
rect 32400 20644 32404 20700
rect 32404 20644 32460 20700
rect 32460 20644 32464 20700
rect 32400 20640 32464 20644
rect 32480 20700 32544 20704
rect 32480 20644 32484 20700
rect 32484 20644 32540 20700
rect 32540 20644 32544 20700
rect 32480 20640 32544 20644
rect 32560 20700 32624 20704
rect 32560 20644 32564 20700
rect 32564 20644 32620 20700
rect 32620 20644 32624 20700
rect 32560 20640 32624 20644
rect 11100 20572 11164 20636
rect 12572 20572 12636 20636
rect 14780 20632 14844 20636
rect 14780 20576 14830 20632
rect 14830 20576 14844 20632
rect 14780 20572 14844 20576
rect 18460 20572 18524 20636
rect 8156 20436 8220 20500
rect 21404 20496 21468 20500
rect 21404 20440 21454 20496
rect 21454 20440 21468 20496
rect 21404 20436 21468 20440
rect 4873 20156 4937 20160
rect 4873 20100 4877 20156
rect 4877 20100 4933 20156
rect 4933 20100 4937 20156
rect 4873 20096 4937 20100
rect 4953 20156 5017 20160
rect 4953 20100 4957 20156
rect 4957 20100 5013 20156
rect 5013 20100 5017 20156
rect 4953 20096 5017 20100
rect 5033 20156 5097 20160
rect 5033 20100 5037 20156
rect 5037 20100 5093 20156
rect 5093 20100 5097 20156
rect 5033 20096 5097 20100
rect 5113 20156 5177 20160
rect 5113 20100 5117 20156
rect 5117 20100 5173 20156
rect 5173 20100 5177 20156
rect 5113 20096 5177 20100
rect 12715 20156 12779 20160
rect 12715 20100 12719 20156
rect 12719 20100 12775 20156
rect 12775 20100 12779 20156
rect 12715 20096 12779 20100
rect 12795 20156 12859 20160
rect 12795 20100 12799 20156
rect 12799 20100 12855 20156
rect 12855 20100 12859 20156
rect 12795 20096 12859 20100
rect 12875 20156 12939 20160
rect 12875 20100 12879 20156
rect 12879 20100 12935 20156
rect 12935 20100 12939 20156
rect 12875 20096 12939 20100
rect 12955 20156 13019 20160
rect 12955 20100 12959 20156
rect 12959 20100 13015 20156
rect 13015 20100 13019 20156
rect 12955 20096 13019 20100
rect 20557 20156 20621 20160
rect 20557 20100 20561 20156
rect 20561 20100 20617 20156
rect 20617 20100 20621 20156
rect 20557 20096 20621 20100
rect 20637 20156 20701 20160
rect 20637 20100 20641 20156
rect 20641 20100 20697 20156
rect 20697 20100 20701 20156
rect 20637 20096 20701 20100
rect 20717 20156 20781 20160
rect 20717 20100 20721 20156
rect 20721 20100 20777 20156
rect 20777 20100 20781 20156
rect 20717 20096 20781 20100
rect 20797 20156 20861 20160
rect 20797 20100 20801 20156
rect 20801 20100 20857 20156
rect 20857 20100 20861 20156
rect 20797 20096 20861 20100
rect 28399 20156 28463 20160
rect 28399 20100 28403 20156
rect 28403 20100 28459 20156
rect 28459 20100 28463 20156
rect 28399 20096 28463 20100
rect 28479 20156 28543 20160
rect 28479 20100 28483 20156
rect 28483 20100 28539 20156
rect 28539 20100 28543 20156
rect 28479 20096 28543 20100
rect 28559 20156 28623 20160
rect 28559 20100 28563 20156
rect 28563 20100 28619 20156
rect 28619 20100 28623 20156
rect 28559 20096 28623 20100
rect 28639 20156 28703 20160
rect 28639 20100 28643 20156
rect 28643 20100 28699 20156
rect 28699 20100 28703 20156
rect 28639 20096 28703 20100
rect 2268 20088 2332 20092
rect 2268 20032 2282 20088
rect 2282 20032 2332 20088
rect 2268 20028 2332 20032
rect 3004 20088 3068 20092
rect 3004 20032 3054 20088
rect 3054 20032 3068 20088
rect 3004 20028 3068 20032
rect 4476 20028 4540 20092
rect 5948 20028 6012 20092
rect 6684 20028 6748 20092
rect 14044 20028 14108 20092
rect 7420 19892 7484 19956
rect 30972 19620 31036 19684
rect 8794 19612 8858 19616
rect 8794 19556 8798 19612
rect 8798 19556 8854 19612
rect 8854 19556 8858 19612
rect 8794 19552 8858 19556
rect 8874 19612 8938 19616
rect 8874 19556 8878 19612
rect 8878 19556 8934 19612
rect 8934 19556 8938 19612
rect 8874 19552 8938 19556
rect 8954 19612 9018 19616
rect 8954 19556 8958 19612
rect 8958 19556 9014 19612
rect 9014 19556 9018 19612
rect 8954 19552 9018 19556
rect 9034 19612 9098 19616
rect 9034 19556 9038 19612
rect 9038 19556 9094 19612
rect 9094 19556 9098 19612
rect 9034 19552 9098 19556
rect 16636 19612 16700 19616
rect 16636 19556 16640 19612
rect 16640 19556 16696 19612
rect 16696 19556 16700 19612
rect 16636 19552 16700 19556
rect 16716 19612 16780 19616
rect 16716 19556 16720 19612
rect 16720 19556 16776 19612
rect 16776 19556 16780 19612
rect 16716 19552 16780 19556
rect 16796 19612 16860 19616
rect 16796 19556 16800 19612
rect 16800 19556 16856 19612
rect 16856 19556 16860 19612
rect 16796 19552 16860 19556
rect 16876 19612 16940 19616
rect 16876 19556 16880 19612
rect 16880 19556 16936 19612
rect 16936 19556 16940 19612
rect 16876 19552 16940 19556
rect 24478 19612 24542 19616
rect 24478 19556 24482 19612
rect 24482 19556 24538 19612
rect 24538 19556 24542 19612
rect 24478 19552 24542 19556
rect 24558 19612 24622 19616
rect 24558 19556 24562 19612
rect 24562 19556 24618 19612
rect 24618 19556 24622 19612
rect 24558 19552 24622 19556
rect 24638 19612 24702 19616
rect 24638 19556 24642 19612
rect 24642 19556 24698 19612
rect 24698 19556 24702 19612
rect 24638 19552 24702 19556
rect 24718 19612 24782 19616
rect 24718 19556 24722 19612
rect 24722 19556 24778 19612
rect 24778 19556 24782 19612
rect 24718 19552 24782 19556
rect 32320 19612 32384 19616
rect 32320 19556 32324 19612
rect 32324 19556 32380 19612
rect 32380 19556 32384 19612
rect 32320 19552 32384 19556
rect 32400 19612 32464 19616
rect 32400 19556 32404 19612
rect 32404 19556 32460 19612
rect 32460 19556 32464 19612
rect 32400 19552 32464 19556
rect 32480 19612 32544 19616
rect 32480 19556 32484 19612
rect 32484 19556 32540 19612
rect 32540 19556 32544 19612
rect 32480 19552 32544 19556
rect 32560 19612 32624 19616
rect 32560 19556 32564 19612
rect 32564 19556 32620 19612
rect 32620 19556 32624 19612
rect 32560 19552 32624 19556
rect 1532 19484 1596 19548
rect 3740 19484 3804 19548
rect 9628 19484 9692 19548
rect 11836 19544 11900 19548
rect 11836 19488 11886 19544
rect 11886 19488 11900 19544
rect 11836 19484 11900 19488
rect 16252 19484 16316 19548
rect 17724 19408 17788 19412
rect 17724 19352 17774 19408
rect 17774 19352 17788 19408
rect 17724 19348 17788 19352
rect 13308 19212 13372 19276
rect 24164 19212 24228 19276
rect 4873 19068 4937 19072
rect 4873 19012 4877 19068
rect 4877 19012 4933 19068
rect 4933 19012 4937 19068
rect 4873 19008 4937 19012
rect 4953 19068 5017 19072
rect 4953 19012 4957 19068
rect 4957 19012 5013 19068
rect 5013 19012 5017 19068
rect 4953 19008 5017 19012
rect 5033 19068 5097 19072
rect 5033 19012 5037 19068
rect 5037 19012 5093 19068
rect 5093 19012 5097 19068
rect 5033 19008 5097 19012
rect 5113 19068 5177 19072
rect 5113 19012 5117 19068
rect 5117 19012 5173 19068
rect 5173 19012 5177 19068
rect 5113 19008 5177 19012
rect 12715 19068 12779 19072
rect 12715 19012 12719 19068
rect 12719 19012 12775 19068
rect 12775 19012 12779 19068
rect 12715 19008 12779 19012
rect 12795 19068 12859 19072
rect 12795 19012 12799 19068
rect 12799 19012 12855 19068
rect 12855 19012 12859 19068
rect 12795 19008 12859 19012
rect 12875 19068 12939 19072
rect 12875 19012 12879 19068
rect 12879 19012 12935 19068
rect 12935 19012 12939 19068
rect 12875 19008 12939 19012
rect 12955 19068 13019 19072
rect 12955 19012 12959 19068
rect 12959 19012 13015 19068
rect 13015 19012 13019 19068
rect 12955 19008 13019 19012
rect 20557 19068 20621 19072
rect 20557 19012 20561 19068
rect 20561 19012 20617 19068
rect 20617 19012 20621 19068
rect 20557 19008 20621 19012
rect 20637 19068 20701 19072
rect 20637 19012 20641 19068
rect 20641 19012 20697 19068
rect 20697 19012 20701 19068
rect 20637 19008 20701 19012
rect 20717 19068 20781 19072
rect 20717 19012 20721 19068
rect 20721 19012 20777 19068
rect 20777 19012 20781 19068
rect 20717 19008 20781 19012
rect 20797 19068 20861 19072
rect 20797 19012 20801 19068
rect 20801 19012 20857 19068
rect 20857 19012 20861 19068
rect 20797 19008 20861 19012
rect 28399 19068 28463 19072
rect 28399 19012 28403 19068
rect 28403 19012 28459 19068
rect 28459 19012 28463 19068
rect 28399 19008 28463 19012
rect 28479 19068 28543 19072
rect 28479 19012 28483 19068
rect 28483 19012 28539 19068
rect 28539 19012 28543 19068
rect 28479 19008 28543 19012
rect 28559 19068 28623 19072
rect 28559 19012 28563 19068
rect 28563 19012 28619 19068
rect 28619 19012 28623 19068
rect 28559 19008 28623 19012
rect 28639 19068 28703 19072
rect 28639 19012 28643 19068
rect 28643 19012 28699 19068
rect 28699 19012 28703 19068
rect 28639 19008 28703 19012
rect 10364 18940 10428 19004
rect 15516 18940 15580 19004
rect 8794 18524 8858 18528
rect 8794 18468 8798 18524
rect 8798 18468 8854 18524
rect 8854 18468 8858 18524
rect 8794 18464 8858 18468
rect 8874 18524 8938 18528
rect 8874 18468 8878 18524
rect 8878 18468 8934 18524
rect 8934 18468 8938 18524
rect 8874 18464 8938 18468
rect 8954 18524 9018 18528
rect 8954 18468 8958 18524
rect 8958 18468 9014 18524
rect 9014 18468 9018 18524
rect 8954 18464 9018 18468
rect 9034 18524 9098 18528
rect 9034 18468 9038 18524
rect 9038 18468 9094 18524
rect 9094 18468 9098 18524
rect 9034 18464 9098 18468
rect 16636 18524 16700 18528
rect 16636 18468 16640 18524
rect 16640 18468 16696 18524
rect 16696 18468 16700 18524
rect 16636 18464 16700 18468
rect 16716 18524 16780 18528
rect 16716 18468 16720 18524
rect 16720 18468 16776 18524
rect 16776 18468 16780 18524
rect 16716 18464 16780 18468
rect 16796 18524 16860 18528
rect 16796 18468 16800 18524
rect 16800 18468 16856 18524
rect 16856 18468 16860 18524
rect 16796 18464 16860 18468
rect 16876 18524 16940 18528
rect 16876 18468 16880 18524
rect 16880 18468 16936 18524
rect 16936 18468 16940 18524
rect 16876 18464 16940 18468
rect 24478 18524 24542 18528
rect 24478 18468 24482 18524
rect 24482 18468 24538 18524
rect 24538 18468 24542 18524
rect 24478 18464 24542 18468
rect 24558 18524 24622 18528
rect 24558 18468 24562 18524
rect 24562 18468 24618 18524
rect 24618 18468 24622 18524
rect 24558 18464 24622 18468
rect 24638 18524 24702 18528
rect 24638 18468 24642 18524
rect 24642 18468 24698 18524
rect 24698 18468 24702 18524
rect 24638 18464 24702 18468
rect 24718 18524 24782 18528
rect 24718 18468 24722 18524
rect 24722 18468 24778 18524
rect 24778 18468 24782 18524
rect 24718 18464 24782 18468
rect 32320 18524 32384 18528
rect 32320 18468 32324 18524
rect 32324 18468 32380 18524
rect 32380 18468 32384 18524
rect 32320 18464 32384 18468
rect 32400 18524 32464 18528
rect 32400 18468 32404 18524
rect 32404 18468 32460 18524
rect 32460 18468 32464 18524
rect 32400 18464 32464 18468
rect 32480 18524 32544 18528
rect 32480 18468 32484 18524
rect 32484 18468 32540 18524
rect 32540 18468 32544 18524
rect 32480 18464 32544 18468
rect 32560 18524 32624 18528
rect 32560 18468 32564 18524
rect 32564 18468 32620 18524
rect 32620 18468 32624 18524
rect 32560 18464 32624 18468
rect 4873 17980 4937 17984
rect 4873 17924 4877 17980
rect 4877 17924 4933 17980
rect 4933 17924 4937 17980
rect 4873 17920 4937 17924
rect 4953 17980 5017 17984
rect 4953 17924 4957 17980
rect 4957 17924 5013 17980
rect 5013 17924 5017 17980
rect 4953 17920 5017 17924
rect 5033 17980 5097 17984
rect 5033 17924 5037 17980
rect 5037 17924 5093 17980
rect 5093 17924 5097 17980
rect 5033 17920 5097 17924
rect 5113 17980 5177 17984
rect 5113 17924 5117 17980
rect 5117 17924 5173 17980
rect 5173 17924 5177 17980
rect 5113 17920 5177 17924
rect 12715 17980 12779 17984
rect 12715 17924 12719 17980
rect 12719 17924 12775 17980
rect 12775 17924 12779 17980
rect 12715 17920 12779 17924
rect 12795 17980 12859 17984
rect 12795 17924 12799 17980
rect 12799 17924 12855 17980
rect 12855 17924 12859 17980
rect 12795 17920 12859 17924
rect 12875 17980 12939 17984
rect 12875 17924 12879 17980
rect 12879 17924 12935 17980
rect 12935 17924 12939 17980
rect 12875 17920 12939 17924
rect 12955 17980 13019 17984
rect 12955 17924 12959 17980
rect 12959 17924 13015 17980
rect 13015 17924 13019 17980
rect 12955 17920 13019 17924
rect 20557 17980 20621 17984
rect 20557 17924 20561 17980
rect 20561 17924 20617 17980
rect 20617 17924 20621 17980
rect 20557 17920 20621 17924
rect 20637 17980 20701 17984
rect 20637 17924 20641 17980
rect 20641 17924 20697 17980
rect 20697 17924 20701 17980
rect 20637 17920 20701 17924
rect 20717 17980 20781 17984
rect 20717 17924 20721 17980
rect 20721 17924 20777 17980
rect 20777 17924 20781 17980
rect 20717 17920 20781 17924
rect 20797 17980 20861 17984
rect 20797 17924 20801 17980
rect 20801 17924 20857 17980
rect 20857 17924 20861 17980
rect 20797 17920 20861 17924
rect 28399 17980 28463 17984
rect 28399 17924 28403 17980
rect 28403 17924 28459 17980
rect 28459 17924 28463 17980
rect 28399 17920 28463 17924
rect 28479 17980 28543 17984
rect 28479 17924 28483 17980
rect 28483 17924 28539 17980
rect 28539 17924 28543 17980
rect 28479 17920 28543 17924
rect 28559 17980 28623 17984
rect 28559 17924 28563 17980
rect 28563 17924 28619 17980
rect 28619 17924 28623 17980
rect 28559 17920 28623 17924
rect 28639 17980 28703 17984
rect 28639 17924 28643 17980
rect 28643 17924 28699 17980
rect 28699 17924 28703 17980
rect 28639 17920 28703 17924
rect 30236 17912 30300 17916
rect 30236 17856 30286 17912
rect 30286 17856 30300 17912
rect 30236 17852 30300 17856
rect 8794 17436 8858 17440
rect 8794 17380 8798 17436
rect 8798 17380 8854 17436
rect 8854 17380 8858 17436
rect 8794 17376 8858 17380
rect 8874 17436 8938 17440
rect 8874 17380 8878 17436
rect 8878 17380 8934 17436
rect 8934 17380 8938 17436
rect 8874 17376 8938 17380
rect 8954 17436 9018 17440
rect 8954 17380 8958 17436
rect 8958 17380 9014 17436
rect 9014 17380 9018 17436
rect 8954 17376 9018 17380
rect 9034 17436 9098 17440
rect 9034 17380 9038 17436
rect 9038 17380 9094 17436
rect 9094 17380 9098 17436
rect 9034 17376 9098 17380
rect 16636 17436 16700 17440
rect 16636 17380 16640 17436
rect 16640 17380 16696 17436
rect 16696 17380 16700 17436
rect 16636 17376 16700 17380
rect 16716 17436 16780 17440
rect 16716 17380 16720 17436
rect 16720 17380 16776 17436
rect 16776 17380 16780 17436
rect 16716 17376 16780 17380
rect 16796 17436 16860 17440
rect 16796 17380 16800 17436
rect 16800 17380 16856 17436
rect 16856 17380 16860 17436
rect 16796 17376 16860 17380
rect 16876 17436 16940 17440
rect 16876 17380 16880 17436
rect 16880 17380 16936 17436
rect 16936 17380 16940 17436
rect 16876 17376 16940 17380
rect 24478 17436 24542 17440
rect 24478 17380 24482 17436
rect 24482 17380 24538 17436
rect 24538 17380 24542 17436
rect 24478 17376 24542 17380
rect 24558 17436 24622 17440
rect 24558 17380 24562 17436
rect 24562 17380 24618 17436
rect 24618 17380 24622 17436
rect 24558 17376 24622 17380
rect 24638 17436 24702 17440
rect 24638 17380 24642 17436
rect 24642 17380 24698 17436
rect 24698 17380 24702 17436
rect 24638 17376 24702 17380
rect 24718 17436 24782 17440
rect 24718 17380 24722 17436
rect 24722 17380 24778 17436
rect 24778 17380 24782 17436
rect 24718 17376 24782 17380
rect 32320 17436 32384 17440
rect 32320 17380 32324 17436
rect 32324 17380 32380 17436
rect 32380 17380 32384 17436
rect 32320 17376 32384 17380
rect 32400 17436 32464 17440
rect 32400 17380 32404 17436
rect 32404 17380 32460 17436
rect 32460 17380 32464 17436
rect 32400 17376 32464 17380
rect 32480 17436 32544 17440
rect 32480 17380 32484 17436
rect 32484 17380 32540 17436
rect 32540 17380 32544 17436
rect 32480 17376 32544 17380
rect 32560 17436 32624 17440
rect 32560 17380 32564 17436
rect 32564 17380 32620 17436
rect 32620 17380 32624 17436
rect 32560 17376 32624 17380
rect 4873 16892 4937 16896
rect 4873 16836 4877 16892
rect 4877 16836 4933 16892
rect 4933 16836 4937 16892
rect 4873 16832 4937 16836
rect 4953 16892 5017 16896
rect 4953 16836 4957 16892
rect 4957 16836 5013 16892
rect 5013 16836 5017 16892
rect 4953 16832 5017 16836
rect 5033 16892 5097 16896
rect 5033 16836 5037 16892
rect 5037 16836 5093 16892
rect 5093 16836 5097 16892
rect 5033 16832 5097 16836
rect 5113 16892 5177 16896
rect 5113 16836 5117 16892
rect 5117 16836 5173 16892
rect 5173 16836 5177 16892
rect 5113 16832 5177 16836
rect 12715 16892 12779 16896
rect 12715 16836 12719 16892
rect 12719 16836 12775 16892
rect 12775 16836 12779 16892
rect 12715 16832 12779 16836
rect 12795 16892 12859 16896
rect 12795 16836 12799 16892
rect 12799 16836 12855 16892
rect 12855 16836 12859 16892
rect 12795 16832 12859 16836
rect 12875 16892 12939 16896
rect 12875 16836 12879 16892
rect 12879 16836 12935 16892
rect 12935 16836 12939 16892
rect 12875 16832 12939 16836
rect 12955 16892 13019 16896
rect 12955 16836 12959 16892
rect 12959 16836 13015 16892
rect 13015 16836 13019 16892
rect 12955 16832 13019 16836
rect 20557 16892 20621 16896
rect 20557 16836 20561 16892
rect 20561 16836 20617 16892
rect 20617 16836 20621 16892
rect 20557 16832 20621 16836
rect 20637 16892 20701 16896
rect 20637 16836 20641 16892
rect 20641 16836 20697 16892
rect 20697 16836 20701 16892
rect 20637 16832 20701 16836
rect 20717 16892 20781 16896
rect 20717 16836 20721 16892
rect 20721 16836 20777 16892
rect 20777 16836 20781 16892
rect 20717 16832 20781 16836
rect 20797 16892 20861 16896
rect 20797 16836 20801 16892
rect 20801 16836 20857 16892
rect 20857 16836 20861 16892
rect 20797 16832 20861 16836
rect 28399 16892 28463 16896
rect 28399 16836 28403 16892
rect 28403 16836 28459 16892
rect 28459 16836 28463 16892
rect 28399 16832 28463 16836
rect 28479 16892 28543 16896
rect 28479 16836 28483 16892
rect 28483 16836 28539 16892
rect 28539 16836 28543 16892
rect 28479 16832 28543 16836
rect 28559 16892 28623 16896
rect 28559 16836 28563 16892
rect 28563 16836 28619 16892
rect 28619 16836 28623 16892
rect 28559 16832 28623 16836
rect 28639 16892 28703 16896
rect 28639 16836 28643 16892
rect 28643 16836 28699 16892
rect 28699 16836 28703 16892
rect 28639 16832 28703 16836
rect 8794 16348 8858 16352
rect 8794 16292 8798 16348
rect 8798 16292 8854 16348
rect 8854 16292 8858 16348
rect 8794 16288 8858 16292
rect 8874 16348 8938 16352
rect 8874 16292 8878 16348
rect 8878 16292 8934 16348
rect 8934 16292 8938 16348
rect 8874 16288 8938 16292
rect 8954 16348 9018 16352
rect 8954 16292 8958 16348
rect 8958 16292 9014 16348
rect 9014 16292 9018 16348
rect 8954 16288 9018 16292
rect 9034 16348 9098 16352
rect 9034 16292 9038 16348
rect 9038 16292 9094 16348
rect 9094 16292 9098 16348
rect 9034 16288 9098 16292
rect 16636 16348 16700 16352
rect 16636 16292 16640 16348
rect 16640 16292 16696 16348
rect 16696 16292 16700 16348
rect 16636 16288 16700 16292
rect 16716 16348 16780 16352
rect 16716 16292 16720 16348
rect 16720 16292 16776 16348
rect 16776 16292 16780 16348
rect 16716 16288 16780 16292
rect 16796 16348 16860 16352
rect 16796 16292 16800 16348
rect 16800 16292 16856 16348
rect 16856 16292 16860 16348
rect 16796 16288 16860 16292
rect 16876 16348 16940 16352
rect 16876 16292 16880 16348
rect 16880 16292 16936 16348
rect 16936 16292 16940 16348
rect 16876 16288 16940 16292
rect 24478 16348 24542 16352
rect 24478 16292 24482 16348
rect 24482 16292 24538 16348
rect 24538 16292 24542 16348
rect 24478 16288 24542 16292
rect 24558 16348 24622 16352
rect 24558 16292 24562 16348
rect 24562 16292 24618 16348
rect 24618 16292 24622 16348
rect 24558 16288 24622 16292
rect 24638 16348 24702 16352
rect 24638 16292 24642 16348
rect 24642 16292 24698 16348
rect 24698 16292 24702 16348
rect 24638 16288 24702 16292
rect 24718 16348 24782 16352
rect 24718 16292 24722 16348
rect 24722 16292 24778 16348
rect 24778 16292 24782 16348
rect 24718 16288 24782 16292
rect 32320 16348 32384 16352
rect 32320 16292 32324 16348
rect 32324 16292 32380 16348
rect 32380 16292 32384 16348
rect 32320 16288 32384 16292
rect 32400 16348 32464 16352
rect 32400 16292 32404 16348
rect 32404 16292 32460 16348
rect 32460 16292 32464 16348
rect 32400 16288 32464 16292
rect 32480 16348 32544 16352
rect 32480 16292 32484 16348
rect 32484 16292 32540 16348
rect 32540 16292 32544 16348
rect 32480 16288 32544 16292
rect 32560 16348 32624 16352
rect 32560 16292 32564 16348
rect 32564 16292 32620 16348
rect 32620 16292 32624 16348
rect 32560 16288 32624 16292
rect 4873 15804 4937 15808
rect 4873 15748 4877 15804
rect 4877 15748 4933 15804
rect 4933 15748 4937 15804
rect 4873 15744 4937 15748
rect 4953 15804 5017 15808
rect 4953 15748 4957 15804
rect 4957 15748 5013 15804
rect 5013 15748 5017 15804
rect 4953 15744 5017 15748
rect 5033 15804 5097 15808
rect 5033 15748 5037 15804
rect 5037 15748 5093 15804
rect 5093 15748 5097 15804
rect 5033 15744 5097 15748
rect 5113 15804 5177 15808
rect 5113 15748 5117 15804
rect 5117 15748 5173 15804
rect 5173 15748 5177 15804
rect 5113 15744 5177 15748
rect 12715 15804 12779 15808
rect 12715 15748 12719 15804
rect 12719 15748 12775 15804
rect 12775 15748 12779 15804
rect 12715 15744 12779 15748
rect 12795 15804 12859 15808
rect 12795 15748 12799 15804
rect 12799 15748 12855 15804
rect 12855 15748 12859 15804
rect 12795 15744 12859 15748
rect 12875 15804 12939 15808
rect 12875 15748 12879 15804
rect 12879 15748 12935 15804
rect 12935 15748 12939 15804
rect 12875 15744 12939 15748
rect 12955 15804 13019 15808
rect 12955 15748 12959 15804
rect 12959 15748 13015 15804
rect 13015 15748 13019 15804
rect 12955 15744 13019 15748
rect 20557 15804 20621 15808
rect 20557 15748 20561 15804
rect 20561 15748 20617 15804
rect 20617 15748 20621 15804
rect 20557 15744 20621 15748
rect 20637 15804 20701 15808
rect 20637 15748 20641 15804
rect 20641 15748 20697 15804
rect 20697 15748 20701 15804
rect 20637 15744 20701 15748
rect 20717 15804 20781 15808
rect 20717 15748 20721 15804
rect 20721 15748 20777 15804
rect 20777 15748 20781 15804
rect 20717 15744 20781 15748
rect 20797 15804 20861 15808
rect 20797 15748 20801 15804
rect 20801 15748 20857 15804
rect 20857 15748 20861 15804
rect 20797 15744 20861 15748
rect 28399 15804 28463 15808
rect 28399 15748 28403 15804
rect 28403 15748 28459 15804
rect 28459 15748 28463 15804
rect 28399 15744 28463 15748
rect 28479 15804 28543 15808
rect 28479 15748 28483 15804
rect 28483 15748 28539 15804
rect 28539 15748 28543 15804
rect 28479 15744 28543 15748
rect 28559 15804 28623 15808
rect 28559 15748 28563 15804
rect 28563 15748 28619 15804
rect 28619 15748 28623 15804
rect 28559 15744 28623 15748
rect 28639 15804 28703 15808
rect 28639 15748 28643 15804
rect 28643 15748 28699 15804
rect 28699 15748 28703 15804
rect 28639 15744 28703 15748
rect 8794 15260 8858 15264
rect 8794 15204 8798 15260
rect 8798 15204 8854 15260
rect 8854 15204 8858 15260
rect 8794 15200 8858 15204
rect 8874 15260 8938 15264
rect 8874 15204 8878 15260
rect 8878 15204 8934 15260
rect 8934 15204 8938 15260
rect 8874 15200 8938 15204
rect 8954 15260 9018 15264
rect 8954 15204 8958 15260
rect 8958 15204 9014 15260
rect 9014 15204 9018 15260
rect 8954 15200 9018 15204
rect 9034 15260 9098 15264
rect 9034 15204 9038 15260
rect 9038 15204 9094 15260
rect 9094 15204 9098 15260
rect 9034 15200 9098 15204
rect 16636 15260 16700 15264
rect 16636 15204 16640 15260
rect 16640 15204 16696 15260
rect 16696 15204 16700 15260
rect 16636 15200 16700 15204
rect 16716 15260 16780 15264
rect 16716 15204 16720 15260
rect 16720 15204 16776 15260
rect 16776 15204 16780 15260
rect 16716 15200 16780 15204
rect 16796 15260 16860 15264
rect 16796 15204 16800 15260
rect 16800 15204 16856 15260
rect 16856 15204 16860 15260
rect 16796 15200 16860 15204
rect 16876 15260 16940 15264
rect 16876 15204 16880 15260
rect 16880 15204 16936 15260
rect 16936 15204 16940 15260
rect 16876 15200 16940 15204
rect 24478 15260 24542 15264
rect 24478 15204 24482 15260
rect 24482 15204 24538 15260
rect 24538 15204 24542 15260
rect 24478 15200 24542 15204
rect 24558 15260 24622 15264
rect 24558 15204 24562 15260
rect 24562 15204 24618 15260
rect 24618 15204 24622 15260
rect 24558 15200 24622 15204
rect 24638 15260 24702 15264
rect 24638 15204 24642 15260
rect 24642 15204 24698 15260
rect 24698 15204 24702 15260
rect 24638 15200 24702 15204
rect 24718 15260 24782 15264
rect 24718 15204 24722 15260
rect 24722 15204 24778 15260
rect 24778 15204 24782 15260
rect 24718 15200 24782 15204
rect 32320 15260 32384 15264
rect 32320 15204 32324 15260
rect 32324 15204 32380 15260
rect 32380 15204 32384 15260
rect 32320 15200 32384 15204
rect 32400 15260 32464 15264
rect 32400 15204 32404 15260
rect 32404 15204 32460 15260
rect 32460 15204 32464 15260
rect 32400 15200 32464 15204
rect 32480 15260 32544 15264
rect 32480 15204 32484 15260
rect 32484 15204 32540 15260
rect 32540 15204 32544 15260
rect 32480 15200 32544 15204
rect 32560 15260 32624 15264
rect 32560 15204 32564 15260
rect 32564 15204 32620 15260
rect 32620 15204 32624 15260
rect 32560 15200 32624 15204
rect 4873 14716 4937 14720
rect 4873 14660 4877 14716
rect 4877 14660 4933 14716
rect 4933 14660 4937 14716
rect 4873 14656 4937 14660
rect 4953 14716 5017 14720
rect 4953 14660 4957 14716
rect 4957 14660 5013 14716
rect 5013 14660 5017 14716
rect 4953 14656 5017 14660
rect 5033 14716 5097 14720
rect 5033 14660 5037 14716
rect 5037 14660 5093 14716
rect 5093 14660 5097 14716
rect 5033 14656 5097 14660
rect 5113 14716 5177 14720
rect 5113 14660 5117 14716
rect 5117 14660 5173 14716
rect 5173 14660 5177 14716
rect 5113 14656 5177 14660
rect 12715 14716 12779 14720
rect 12715 14660 12719 14716
rect 12719 14660 12775 14716
rect 12775 14660 12779 14716
rect 12715 14656 12779 14660
rect 12795 14716 12859 14720
rect 12795 14660 12799 14716
rect 12799 14660 12855 14716
rect 12855 14660 12859 14716
rect 12795 14656 12859 14660
rect 12875 14716 12939 14720
rect 12875 14660 12879 14716
rect 12879 14660 12935 14716
rect 12935 14660 12939 14716
rect 12875 14656 12939 14660
rect 12955 14716 13019 14720
rect 12955 14660 12959 14716
rect 12959 14660 13015 14716
rect 13015 14660 13019 14716
rect 12955 14656 13019 14660
rect 20557 14716 20621 14720
rect 20557 14660 20561 14716
rect 20561 14660 20617 14716
rect 20617 14660 20621 14716
rect 20557 14656 20621 14660
rect 20637 14716 20701 14720
rect 20637 14660 20641 14716
rect 20641 14660 20697 14716
rect 20697 14660 20701 14716
rect 20637 14656 20701 14660
rect 20717 14716 20781 14720
rect 20717 14660 20721 14716
rect 20721 14660 20777 14716
rect 20777 14660 20781 14716
rect 20717 14656 20781 14660
rect 20797 14716 20861 14720
rect 20797 14660 20801 14716
rect 20801 14660 20857 14716
rect 20857 14660 20861 14716
rect 20797 14656 20861 14660
rect 28399 14716 28463 14720
rect 28399 14660 28403 14716
rect 28403 14660 28459 14716
rect 28459 14660 28463 14716
rect 28399 14656 28463 14660
rect 28479 14716 28543 14720
rect 28479 14660 28483 14716
rect 28483 14660 28539 14716
rect 28539 14660 28543 14716
rect 28479 14656 28543 14660
rect 28559 14716 28623 14720
rect 28559 14660 28563 14716
rect 28563 14660 28619 14716
rect 28619 14660 28623 14716
rect 28559 14656 28623 14660
rect 28639 14716 28703 14720
rect 28639 14660 28643 14716
rect 28643 14660 28699 14716
rect 28699 14660 28703 14716
rect 28639 14656 28703 14660
rect 8794 14172 8858 14176
rect 8794 14116 8798 14172
rect 8798 14116 8854 14172
rect 8854 14116 8858 14172
rect 8794 14112 8858 14116
rect 8874 14172 8938 14176
rect 8874 14116 8878 14172
rect 8878 14116 8934 14172
rect 8934 14116 8938 14172
rect 8874 14112 8938 14116
rect 8954 14172 9018 14176
rect 8954 14116 8958 14172
rect 8958 14116 9014 14172
rect 9014 14116 9018 14172
rect 8954 14112 9018 14116
rect 9034 14172 9098 14176
rect 9034 14116 9038 14172
rect 9038 14116 9094 14172
rect 9094 14116 9098 14172
rect 9034 14112 9098 14116
rect 16636 14172 16700 14176
rect 16636 14116 16640 14172
rect 16640 14116 16696 14172
rect 16696 14116 16700 14172
rect 16636 14112 16700 14116
rect 16716 14172 16780 14176
rect 16716 14116 16720 14172
rect 16720 14116 16776 14172
rect 16776 14116 16780 14172
rect 16716 14112 16780 14116
rect 16796 14172 16860 14176
rect 16796 14116 16800 14172
rect 16800 14116 16856 14172
rect 16856 14116 16860 14172
rect 16796 14112 16860 14116
rect 16876 14172 16940 14176
rect 16876 14116 16880 14172
rect 16880 14116 16936 14172
rect 16936 14116 16940 14172
rect 16876 14112 16940 14116
rect 24478 14172 24542 14176
rect 24478 14116 24482 14172
rect 24482 14116 24538 14172
rect 24538 14116 24542 14172
rect 24478 14112 24542 14116
rect 24558 14172 24622 14176
rect 24558 14116 24562 14172
rect 24562 14116 24618 14172
rect 24618 14116 24622 14172
rect 24558 14112 24622 14116
rect 24638 14172 24702 14176
rect 24638 14116 24642 14172
rect 24642 14116 24698 14172
rect 24698 14116 24702 14172
rect 24638 14112 24702 14116
rect 24718 14172 24782 14176
rect 24718 14116 24722 14172
rect 24722 14116 24778 14172
rect 24778 14116 24782 14172
rect 24718 14112 24782 14116
rect 32320 14172 32384 14176
rect 32320 14116 32324 14172
rect 32324 14116 32380 14172
rect 32380 14116 32384 14172
rect 32320 14112 32384 14116
rect 32400 14172 32464 14176
rect 32400 14116 32404 14172
rect 32404 14116 32460 14172
rect 32460 14116 32464 14172
rect 32400 14112 32464 14116
rect 32480 14172 32544 14176
rect 32480 14116 32484 14172
rect 32484 14116 32540 14172
rect 32540 14116 32544 14172
rect 32480 14112 32544 14116
rect 32560 14172 32624 14176
rect 32560 14116 32564 14172
rect 32564 14116 32620 14172
rect 32620 14116 32624 14172
rect 32560 14112 32624 14116
rect 4873 13628 4937 13632
rect 4873 13572 4877 13628
rect 4877 13572 4933 13628
rect 4933 13572 4937 13628
rect 4873 13568 4937 13572
rect 4953 13628 5017 13632
rect 4953 13572 4957 13628
rect 4957 13572 5013 13628
rect 5013 13572 5017 13628
rect 4953 13568 5017 13572
rect 5033 13628 5097 13632
rect 5033 13572 5037 13628
rect 5037 13572 5093 13628
rect 5093 13572 5097 13628
rect 5033 13568 5097 13572
rect 5113 13628 5177 13632
rect 5113 13572 5117 13628
rect 5117 13572 5173 13628
rect 5173 13572 5177 13628
rect 5113 13568 5177 13572
rect 12715 13628 12779 13632
rect 12715 13572 12719 13628
rect 12719 13572 12775 13628
rect 12775 13572 12779 13628
rect 12715 13568 12779 13572
rect 12795 13628 12859 13632
rect 12795 13572 12799 13628
rect 12799 13572 12855 13628
rect 12855 13572 12859 13628
rect 12795 13568 12859 13572
rect 12875 13628 12939 13632
rect 12875 13572 12879 13628
rect 12879 13572 12935 13628
rect 12935 13572 12939 13628
rect 12875 13568 12939 13572
rect 12955 13628 13019 13632
rect 12955 13572 12959 13628
rect 12959 13572 13015 13628
rect 13015 13572 13019 13628
rect 12955 13568 13019 13572
rect 20557 13628 20621 13632
rect 20557 13572 20561 13628
rect 20561 13572 20617 13628
rect 20617 13572 20621 13628
rect 20557 13568 20621 13572
rect 20637 13628 20701 13632
rect 20637 13572 20641 13628
rect 20641 13572 20697 13628
rect 20697 13572 20701 13628
rect 20637 13568 20701 13572
rect 20717 13628 20781 13632
rect 20717 13572 20721 13628
rect 20721 13572 20777 13628
rect 20777 13572 20781 13628
rect 20717 13568 20781 13572
rect 20797 13628 20861 13632
rect 20797 13572 20801 13628
rect 20801 13572 20857 13628
rect 20857 13572 20861 13628
rect 20797 13568 20861 13572
rect 28399 13628 28463 13632
rect 28399 13572 28403 13628
rect 28403 13572 28459 13628
rect 28459 13572 28463 13628
rect 28399 13568 28463 13572
rect 28479 13628 28543 13632
rect 28479 13572 28483 13628
rect 28483 13572 28539 13628
rect 28539 13572 28543 13628
rect 28479 13568 28543 13572
rect 28559 13628 28623 13632
rect 28559 13572 28563 13628
rect 28563 13572 28619 13628
rect 28619 13572 28623 13628
rect 28559 13568 28623 13572
rect 28639 13628 28703 13632
rect 28639 13572 28643 13628
rect 28643 13572 28699 13628
rect 28699 13572 28703 13628
rect 28639 13568 28703 13572
rect 8794 13084 8858 13088
rect 8794 13028 8798 13084
rect 8798 13028 8854 13084
rect 8854 13028 8858 13084
rect 8794 13024 8858 13028
rect 8874 13084 8938 13088
rect 8874 13028 8878 13084
rect 8878 13028 8934 13084
rect 8934 13028 8938 13084
rect 8874 13024 8938 13028
rect 8954 13084 9018 13088
rect 8954 13028 8958 13084
rect 8958 13028 9014 13084
rect 9014 13028 9018 13084
rect 8954 13024 9018 13028
rect 9034 13084 9098 13088
rect 9034 13028 9038 13084
rect 9038 13028 9094 13084
rect 9094 13028 9098 13084
rect 9034 13024 9098 13028
rect 16636 13084 16700 13088
rect 16636 13028 16640 13084
rect 16640 13028 16696 13084
rect 16696 13028 16700 13084
rect 16636 13024 16700 13028
rect 16716 13084 16780 13088
rect 16716 13028 16720 13084
rect 16720 13028 16776 13084
rect 16776 13028 16780 13084
rect 16716 13024 16780 13028
rect 16796 13084 16860 13088
rect 16796 13028 16800 13084
rect 16800 13028 16856 13084
rect 16856 13028 16860 13084
rect 16796 13024 16860 13028
rect 16876 13084 16940 13088
rect 16876 13028 16880 13084
rect 16880 13028 16936 13084
rect 16936 13028 16940 13084
rect 16876 13024 16940 13028
rect 24478 13084 24542 13088
rect 24478 13028 24482 13084
rect 24482 13028 24538 13084
rect 24538 13028 24542 13084
rect 24478 13024 24542 13028
rect 24558 13084 24622 13088
rect 24558 13028 24562 13084
rect 24562 13028 24618 13084
rect 24618 13028 24622 13084
rect 24558 13024 24622 13028
rect 24638 13084 24702 13088
rect 24638 13028 24642 13084
rect 24642 13028 24698 13084
rect 24698 13028 24702 13084
rect 24638 13024 24702 13028
rect 24718 13084 24782 13088
rect 24718 13028 24722 13084
rect 24722 13028 24778 13084
rect 24778 13028 24782 13084
rect 24718 13024 24782 13028
rect 32320 13084 32384 13088
rect 32320 13028 32324 13084
rect 32324 13028 32380 13084
rect 32380 13028 32384 13084
rect 32320 13024 32384 13028
rect 32400 13084 32464 13088
rect 32400 13028 32404 13084
rect 32404 13028 32460 13084
rect 32460 13028 32464 13084
rect 32400 13024 32464 13028
rect 32480 13084 32544 13088
rect 32480 13028 32484 13084
rect 32484 13028 32540 13084
rect 32540 13028 32544 13084
rect 32480 13024 32544 13028
rect 32560 13084 32624 13088
rect 32560 13028 32564 13084
rect 32564 13028 32620 13084
rect 32620 13028 32624 13084
rect 32560 13024 32624 13028
rect 4873 12540 4937 12544
rect 4873 12484 4877 12540
rect 4877 12484 4933 12540
rect 4933 12484 4937 12540
rect 4873 12480 4937 12484
rect 4953 12540 5017 12544
rect 4953 12484 4957 12540
rect 4957 12484 5013 12540
rect 5013 12484 5017 12540
rect 4953 12480 5017 12484
rect 5033 12540 5097 12544
rect 5033 12484 5037 12540
rect 5037 12484 5093 12540
rect 5093 12484 5097 12540
rect 5033 12480 5097 12484
rect 5113 12540 5177 12544
rect 5113 12484 5117 12540
rect 5117 12484 5173 12540
rect 5173 12484 5177 12540
rect 5113 12480 5177 12484
rect 12715 12540 12779 12544
rect 12715 12484 12719 12540
rect 12719 12484 12775 12540
rect 12775 12484 12779 12540
rect 12715 12480 12779 12484
rect 12795 12540 12859 12544
rect 12795 12484 12799 12540
rect 12799 12484 12855 12540
rect 12855 12484 12859 12540
rect 12795 12480 12859 12484
rect 12875 12540 12939 12544
rect 12875 12484 12879 12540
rect 12879 12484 12935 12540
rect 12935 12484 12939 12540
rect 12875 12480 12939 12484
rect 12955 12540 13019 12544
rect 12955 12484 12959 12540
rect 12959 12484 13015 12540
rect 13015 12484 13019 12540
rect 12955 12480 13019 12484
rect 20557 12540 20621 12544
rect 20557 12484 20561 12540
rect 20561 12484 20617 12540
rect 20617 12484 20621 12540
rect 20557 12480 20621 12484
rect 20637 12540 20701 12544
rect 20637 12484 20641 12540
rect 20641 12484 20697 12540
rect 20697 12484 20701 12540
rect 20637 12480 20701 12484
rect 20717 12540 20781 12544
rect 20717 12484 20721 12540
rect 20721 12484 20777 12540
rect 20777 12484 20781 12540
rect 20717 12480 20781 12484
rect 20797 12540 20861 12544
rect 20797 12484 20801 12540
rect 20801 12484 20857 12540
rect 20857 12484 20861 12540
rect 20797 12480 20861 12484
rect 28399 12540 28463 12544
rect 28399 12484 28403 12540
rect 28403 12484 28459 12540
rect 28459 12484 28463 12540
rect 28399 12480 28463 12484
rect 28479 12540 28543 12544
rect 28479 12484 28483 12540
rect 28483 12484 28539 12540
rect 28539 12484 28543 12540
rect 28479 12480 28543 12484
rect 28559 12540 28623 12544
rect 28559 12484 28563 12540
rect 28563 12484 28619 12540
rect 28619 12484 28623 12540
rect 28559 12480 28623 12484
rect 28639 12540 28703 12544
rect 28639 12484 28643 12540
rect 28643 12484 28699 12540
rect 28699 12484 28703 12540
rect 28639 12480 28703 12484
rect 8794 11996 8858 12000
rect 8794 11940 8798 11996
rect 8798 11940 8854 11996
rect 8854 11940 8858 11996
rect 8794 11936 8858 11940
rect 8874 11996 8938 12000
rect 8874 11940 8878 11996
rect 8878 11940 8934 11996
rect 8934 11940 8938 11996
rect 8874 11936 8938 11940
rect 8954 11996 9018 12000
rect 8954 11940 8958 11996
rect 8958 11940 9014 11996
rect 9014 11940 9018 11996
rect 8954 11936 9018 11940
rect 9034 11996 9098 12000
rect 9034 11940 9038 11996
rect 9038 11940 9094 11996
rect 9094 11940 9098 11996
rect 9034 11936 9098 11940
rect 16636 11996 16700 12000
rect 16636 11940 16640 11996
rect 16640 11940 16696 11996
rect 16696 11940 16700 11996
rect 16636 11936 16700 11940
rect 16716 11996 16780 12000
rect 16716 11940 16720 11996
rect 16720 11940 16776 11996
rect 16776 11940 16780 11996
rect 16716 11936 16780 11940
rect 16796 11996 16860 12000
rect 16796 11940 16800 11996
rect 16800 11940 16856 11996
rect 16856 11940 16860 11996
rect 16796 11936 16860 11940
rect 16876 11996 16940 12000
rect 16876 11940 16880 11996
rect 16880 11940 16936 11996
rect 16936 11940 16940 11996
rect 16876 11936 16940 11940
rect 24478 11996 24542 12000
rect 24478 11940 24482 11996
rect 24482 11940 24538 11996
rect 24538 11940 24542 11996
rect 24478 11936 24542 11940
rect 24558 11996 24622 12000
rect 24558 11940 24562 11996
rect 24562 11940 24618 11996
rect 24618 11940 24622 11996
rect 24558 11936 24622 11940
rect 24638 11996 24702 12000
rect 24638 11940 24642 11996
rect 24642 11940 24698 11996
rect 24698 11940 24702 11996
rect 24638 11936 24702 11940
rect 24718 11996 24782 12000
rect 24718 11940 24722 11996
rect 24722 11940 24778 11996
rect 24778 11940 24782 11996
rect 24718 11936 24782 11940
rect 32320 11996 32384 12000
rect 32320 11940 32324 11996
rect 32324 11940 32380 11996
rect 32380 11940 32384 11996
rect 32320 11936 32384 11940
rect 32400 11996 32464 12000
rect 32400 11940 32404 11996
rect 32404 11940 32460 11996
rect 32460 11940 32464 11996
rect 32400 11936 32464 11940
rect 32480 11996 32544 12000
rect 32480 11940 32484 11996
rect 32484 11940 32540 11996
rect 32540 11940 32544 11996
rect 32480 11936 32544 11940
rect 32560 11996 32624 12000
rect 32560 11940 32564 11996
rect 32564 11940 32620 11996
rect 32620 11940 32624 11996
rect 32560 11936 32624 11940
rect 4873 11452 4937 11456
rect 4873 11396 4877 11452
rect 4877 11396 4933 11452
rect 4933 11396 4937 11452
rect 4873 11392 4937 11396
rect 4953 11452 5017 11456
rect 4953 11396 4957 11452
rect 4957 11396 5013 11452
rect 5013 11396 5017 11452
rect 4953 11392 5017 11396
rect 5033 11452 5097 11456
rect 5033 11396 5037 11452
rect 5037 11396 5093 11452
rect 5093 11396 5097 11452
rect 5033 11392 5097 11396
rect 5113 11452 5177 11456
rect 5113 11396 5117 11452
rect 5117 11396 5173 11452
rect 5173 11396 5177 11452
rect 5113 11392 5177 11396
rect 12715 11452 12779 11456
rect 12715 11396 12719 11452
rect 12719 11396 12775 11452
rect 12775 11396 12779 11452
rect 12715 11392 12779 11396
rect 12795 11452 12859 11456
rect 12795 11396 12799 11452
rect 12799 11396 12855 11452
rect 12855 11396 12859 11452
rect 12795 11392 12859 11396
rect 12875 11452 12939 11456
rect 12875 11396 12879 11452
rect 12879 11396 12935 11452
rect 12935 11396 12939 11452
rect 12875 11392 12939 11396
rect 12955 11452 13019 11456
rect 12955 11396 12959 11452
rect 12959 11396 13015 11452
rect 13015 11396 13019 11452
rect 12955 11392 13019 11396
rect 20557 11452 20621 11456
rect 20557 11396 20561 11452
rect 20561 11396 20617 11452
rect 20617 11396 20621 11452
rect 20557 11392 20621 11396
rect 20637 11452 20701 11456
rect 20637 11396 20641 11452
rect 20641 11396 20697 11452
rect 20697 11396 20701 11452
rect 20637 11392 20701 11396
rect 20717 11452 20781 11456
rect 20717 11396 20721 11452
rect 20721 11396 20777 11452
rect 20777 11396 20781 11452
rect 20717 11392 20781 11396
rect 20797 11452 20861 11456
rect 20797 11396 20801 11452
rect 20801 11396 20857 11452
rect 20857 11396 20861 11452
rect 20797 11392 20861 11396
rect 28399 11452 28463 11456
rect 28399 11396 28403 11452
rect 28403 11396 28459 11452
rect 28459 11396 28463 11452
rect 28399 11392 28463 11396
rect 28479 11452 28543 11456
rect 28479 11396 28483 11452
rect 28483 11396 28539 11452
rect 28539 11396 28543 11452
rect 28479 11392 28543 11396
rect 28559 11452 28623 11456
rect 28559 11396 28563 11452
rect 28563 11396 28619 11452
rect 28619 11396 28623 11452
rect 28559 11392 28623 11396
rect 28639 11452 28703 11456
rect 28639 11396 28643 11452
rect 28643 11396 28699 11452
rect 28699 11396 28703 11452
rect 28639 11392 28703 11396
rect 8794 10908 8858 10912
rect 8794 10852 8798 10908
rect 8798 10852 8854 10908
rect 8854 10852 8858 10908
rect 8794 10848 8858 10852
rect 8874 10908 8938 10912
rect 8874 10852 8878 10908
rect 8878 10852 8934 10908
rect 8934 10852 8938 10908
rect 8874 10848 8938 10852
rect 8954 10908 9018 10912
rect 8954 10852 8958 10908
rect 8958 10852 9014 10908
rect 9014 10852 9018 10908
rect 8954 10848 9018 10852
rect 9034 10908 9098 10912
rect 9034 10852 9038 10908
rect 9038 10852 9094 10908
rect 9094 10852 9098 10908
rect 9034 10848 9098 10852
rect 16636 10908 16700 10912
rect 16636 10852 16640 10908
rect 16640 10852 16696 10908
rect 16696 10852 16700 10908
rect 16636 10848 16700 10852
rect 16716 10908 16780 10912
rect 16716 10852 16720 10908
rect 16720 10852 16776 10908
rect 16776 10852 16780 10908
rect 16716 10848 16780 10852
rect 16796 10908 16860 10912
rect 16796 10852 16800 10908
rect 16800 10852 16856 10908
rect 16856 10852 16860 10908
rect 16796 10848 16860 10852
rect 16876 10908 16940 10912
rect 16876 10852 16880 10908
rect 16880 10852 16936 10908
rect 16936 10852 16940 10908
rect 16876 10848 16940 10852
rect 24478 10908 24542 10912
rect 24478 10852 24482 10908
rect 24482 10852 24538 10908
rect 24538 10852 24542 10908
rect 24478 10848 24542 10852
rect 24558 10908 24622 10912
rect 24558 10852 24562 10908
rect 24562 10852 24618 10908
rect 24618 10852 24622 10908
rect 24558 10848 24622 10852
rect 24638 10908 24702 10912
rect 24638 10852 24642 10908
rect 24642 10852 24698 10908
rect 24698 10852 24702 10908
rect 24638 10848 24702 10852
rect 24718 10908 24782 10912
rect 24718 10852 24722 10908
rect 24722 10852 24778 10908
rect 24778 10852 24782 10908
rect 24718 10848 24782 10852
rect 32320 10908 32384 10912
rect 32320 10852 32324 10908
rect 32324 10852 32380 10908
rect 32380 10852 32384 10908
rect 32320 10848 32384 10852
rect 32400 10908 32464 10912
rect 32400 10852 32404 10908
rect 32404 10852 32460 10908
rect 32460 10852 32464 10908
rect 32400 10848 32464 10852
rect 32480 10908 32544 10912
rect 32480 10852 32484 10908
rect 32484 10852 32540 10908
rect 32540 10852 32544 10908
rect 32480 10848 32544 10852
rect 32560 10908 32624 10912
rect 32560 10852 32564 10908
rect 32564 10852 32620 10908
rect 32620 10852 32624 10908
rect 32560 10848 32624 10852
rect 4873 10364 4937 10368
rect 4873 10308 4877 10364
rect 4877 10308 4933 10364
rect 4933 10308 4937 10364
rect 4873 10304 4937 10308
rect 4953 10364 5017 10368
rect 4953 10308 4957 10364
rect 4957 10308 5013 10364
rect 5013 10308 5017 10364
rect 4953 10304 5017 10308
rect 5033 10364 5097 10368
rect 5033 10308 5037 10364
rect 5037 10308 5093 10364
rect 5093 10308 5097 10364
rect 5033 10304 5097 10308
rect 5113 10364 5177 10368
rect 5113 10308 5117 10364
rect 5117 10308 5173 10364
rect 5173 10308 5177 10364
rect 5113 10304 5177 10308
rect 12715 10364 12779 10368
rect 12715 10308 12719 10364
rect 12719 10308 12775 10364
rect 12775 10308 12779 10364
rect 12715 10304 12779 10308
rect 12795 10364 12859 10368
rect 12795 10308 12799 10364
rect 12799 10308 12855 10364
rect 12855 10308 12859 10364
rect 12795 10304 12859 10308
rect 12875 10364 12939 10368
rect 12875 10308 12879 10364
rect 12879 10308 12935 10364
rect 12935 10308 12939 10364
rect 12875 10304 12939 10308
rect 12955 10364 13019 10368
rect 12955 10308 12959 10364
rect 12959 10308 13015 10364
rect 13015 10308 13019 10364
rect 12955 10304 13019 10308
rect 20557 10364 20621 10368
rect 20557 10308 20561 10364
rect 20561 10308 20617 10364
rect 20617 10308 20621 10364
rect 20557 10304 20621 10308
rect 20637 10364 20701 10368
rect 20637 10308 20641 10364
rect 20641 10308 20697 10364
rect 20697 10308 20701 10364
rect 20637 10304 20701 10308
rect 20717 10364 20781 10368
rect 20717 10308 20721 10364
rect 20721 10308 20777 10364
rect 20777 10308 20781 10364
rect 20717 10304 20781 10308
rect 20797 10364 20861 10368
rect 20797 10308 20801 10364
rect 20801 10308 20857 10364
rect 20857 10308 20861 10364
rect 20797 10304 20861 10308
rect 28399 10364 28463 10368
rect 28399 10308 28403 10364
rect 28403 10308 28459 10364
rect 28459 10308 28463 10364
rect 28399 10304 28463 10308
rect 28479 10364 28543 10368
rect 28479 10308 28483 10364
rect 28483 10308 28539 10364
rect 28539 10308 28543 10364
rect 28479 10304 28543 10308
rect 28559 10364 28623 10368
rect 28559 10308 28563 10364
rect 28563 10308 28619 10364
rect 28619 10308 28623 10364
rect 28559 10304 28623 10308
rect 28639 10364 28703 10368
rect 28639 10308 28643 10364
rect 28643 10308 28699 10364
rect 28699 10308 28703 10364
rect 28639 10304 28703 10308
rect 8794 9820 8858 9824
rect 8794 9764 8798 9820
rect 8798 9764 8854 9820
rect 8854 9764 8858 9820
rect 8794 9760 8858 9764
rect 8874 9820 8938 9824
rect 8874 9764 8878 9820
rect 8878 9764 8934 9820
rect 8934 9764 8938 9820
rect 8874 9760 8938 9764
rect 8954 9820 9018 9824
rect 8954 9764 8958 9820
rect 8958 9764 9014 9820
rect 9014 9764 9018 9820
rect 8954 9760 9018 9764
rect 9034 9820 9098 9824
rect 9034 9764 9038 9820
rect 9038 9764 9094 9820
rect 9094 9764 9098 9820
rect 9034 9760 9098 9764
rect 16636 9820 16700 9824
rect 16636 9764 16640 9820
rect 16640 9764 16696 9820
rect 16696 9764 16700 9820
rect 16636 9760 16700 9764
rect 16716 9820 16780 9824
rect 16716 9764 16720 9820
rect 16720 9764 16776 9820
rect 16776 9764 16780 9820
rect 16716 9760 16780 9764
rect 16796 9820 16860 9824
rect 16796 9764 16800 9820
rect 16800 9764 16856 9820
rect 16856 9764 16860 9820
rect 16796 9760 16860 9764
rect 16876 9820 16940 9824
rect 16876 9764 16880 9820
rect 16880 9764 16936 9820
rect 16936 9764 16940 9820
rect 16876 9760 16940 9764
rect 24478 9820 24542 9824
rect 24478 9764 24482 9820
rect 24482 9764 24538 9820
rect 24538 9764 24542 9820
rect 24478 9760 24542 9764
rect 24558 9820 24622 9824
rect 24558 9764 24562 9820
rect 24562 9764 24618 9820
rect 24618 9764 24622 9820
rect 24558 9760 24622 9764
rect 24638 9820 24702 9824
rect 24638 9764 24642 9820
rect 24642 9764 24698 9820
rect 24698 9764 24702 9820
rect 24638 9760 24702 9764
rect 24718 9820 24782 9824
rect 24718 9764 24722 9820
rect 24722 9764 24778 9820
rect 24778 9764 24782 9820
rect 24718 9760 24782 9764
rect 32320 9820 32384 9824
rect 32320 9764 32324 9820
rect 32324 9764 32380 9820
rect 32380 9764 32384 9820
rect 32320 9760 32384 9764
rect 32400 9820 32464 9824
rect 32400 9764 32404 9820
rect 32404 9764 32460 9820
rect 32460 9764 32464 9820
rect 32400 9760 32464 9764
rect 32480 9820 32544 9824
rect 32480 9764 32484 9820
rect 32484 9764 32540 9820
rect 32540 9764 32544 9820
rect 32480 9760 32544 9764
rect 32560 9820 32624 9824
rect 32560 9764 32564 9820
rect 32564 9764 32620 9820
rect 32620 9764 32624 9820
rect 32560 9760 32624 9764
rect 4873 9276 4937 9280
rect 4873 9220 4877 9276
rect 4877 9220 4933 9276
rect 4933 9220 4937 9276
rect 4873 9216 4937 9220
rect 4953 9276 5017 9280
rect 4953 9220 4957 9276
rect 4957 9220 5013 9276
rect 5013 9220 5017 9276
rect 4953 9216 5017 9220
rect 5033 9276 5097 9280
rect 5033 9220 5037 9276
rect 5037 9220 5093 9276
rect 5093 9220 5097 9276
rect 5033 9216 5097 9220
rect 5113 9276 5177 9280
rect 5113 9220 5117 9276
rect 5117 9220 5173 9276
rect 5173 9220 5177 9276
rect 5113 9216 5177 9220
rect 12715 9276 12779 9280
rect 12715 9220 12719 9276
rect 12719 9220 12775 9276
rect 12775 9220 12779 9276
rect 12715 9216 12779 9220
rect 12795 9276 12859 9280
rect 12795 9220 12799 9276
rect 12799 9220 12855 9276
rect 12855 9220 12859 9276
rect 12795 9216 12859 9220
rect 12875 9276 12939 9280
rect 12875 9220 12879 9276
rect 12879 9220 12935 9276
rect 12935 9220 12939 9276
rect 12875 9216 12939 9220
rect 12955 9276 13019 9280
rect 12955 9220 12959 9276
rect 12959 9220 13015 9276
rect 13015 9220 13019 9276
rect 12955 9216 13019 9220
rect 20557 9276 20621 9280
rect 20557 9220 20561 9276
rect 20561 9220 20617 9276
rect 20617 9220 20621 9276
rect 20557 9216 20621 9220
rect 20637 9276 20701 9280
rect 20637 9220 20641 9276
rect 20641 9220 20697 9276
rect 20697 9220 20701 9276
rect 20637 9216 20701 9220
rect 20717 9276 20781 9280
rect 20717 9220 20721 9276
rect 20721 9220 20777 9276
rect 20777 9220 20781 9276
rect 20717 9216 20781 9220
rect 20797 9276 20861 9280
rect 20797 9220 20801 9276
rect 20801 9220 20857 9276
rect 20857 9220 20861 9276
rect 20797 9216 20861 9220
rect 28399 9276 28463 9280
rect 28399 9220 28403 9276
rect 28403 9220 28459 9276
rect 28459 9220 28463 9276
rect 28399 9216 28463 9220
rect 28479 9276 28543 9280
rect 28479 9220 28483 9276
rect 28483 9220 28539 9276
rect 28539 9220 28543 9276
rect 28479 9216 28543 9220
rect 28559 9276 28623 9280
rect 28559 9220 28563 9276
rect 28563 9220 28619 9276
rect 28619 9220 28623 9276
rect 28559 9216 28623 9220
rect 28639 9276 28703 9280
rect 28639 9220 28643 9276
rect 28643 9220 28699 9276
rect 28699 9220 28703 9276
rect 28639 9216 28703 9220
rect 8794 8732 8858 8736
rect 8794 8676 8798 8732
rect 8798 8676 8854 8732
rect 8854 8676 8858 8732
rect 8794 8672 8858 8676
rect 8874 8732 8938 8736
rect 8874 8676 8878 8732
rect 8878 8676 8934 8732
rect 8934 8676 8938 8732
rect 8874 8672 8938 8676
rect 8954 8732 9018 8736
rect 8954 8676 8958 8732
rect 8958 8676 9014 8732
rect 9014 8676 9018 8732
rect 8954 8672 9018 8676
rect 9034 8732 9098 8736
rect 9034 8676 9038 8732
rect 9038 8676 9094 8732
rect 9094 8676 9098 8732
rect 9034 8672 9098 8676
rect 16636 8732 16700 8736
rect 16636 8676 16640 8732
rect 16640 8676 16696 8732
rect 16696 8676 16700 8732
rect 16636 8672 16700 8676
rect 16716 8732 16780 8736
rect 16716 8676 16720 8732
rect 16720 8676 16776 8732
rect 16776 8676 16780 8732
rect 16716 8672 16780 8676
rect 16796 8732 16860 8736
rect 16796 8676 16800 8732
rect 16800 8676 16856 8732
rect 16856 8676 16860 8732
rect 16796 8672 16860 8676
rect 16876 8732 16940 8736
rect 16876 8676 16880 8732
rect 16880 8676 16936 8732
rect 16936 8676 16940 8732
rect 16876 8672 16940 8676
rect 24478 8732 24542 8736
rect 24478 8676 24482 8732
rect 24482 8676 24538 8732
rect 24538 8676 24542 8732
rect 24478 8672 24542 8676
rect 24558 8732 24622 8736
rect 24558 8676 24562 8732
rect 24562 8676 24618 8732
rect 24618 8676 24622 8732
rect 24558 8672 24622 8676
rect 24638 8732 24702 8736
rect 24638 8676 24642 8732
rect 24642 8676 24698 8732
rect 24698 8676 24702 8732
rect 24638 8672 24702 8676
rect 24718 8732 24782 8736
rect 24718 8676 24722 8732
rect 24722 8676 24778 8732
rect 24778 8676 24782 8732
rect 24718 8672 24782 8676
rect 32320 8732 32384 8736
rect 32320 8676 32324 8732
rect 32324 8676 32380 8732
rect 32380 8676 32384 8732
rect 32320 8672 32384 8676
rect 32400 8732 32464 8736
rect 32400 8676 32404 8732
rect 32404 8676 32460 8732
rect 32460 8676 32464 8732
rect 32400 8672 32464 8676
rect 32480 8732 32544 8736
rect 32480 8676 32484 8732
rect 32484 8676 32540 8732
rect 32540 8676 32544 8732
rect 32480 8672 32544 8676
rect 32560 8732 32624 8736
rect 32560 8676 32564 8732
rect 32564 8676 32620 8732
rect 32620 8676 32624 8732
rect 32560 8672 32624 8676
rect 4873 8188 4937 8192
rect 4873 8132 4877 8188
rect 4877 8132 4933 8188
rect 4933 8132 4937 8188
rect 4873 8128 4937 8132
rect 4953 8188 5017 8192
rect 4953 8132 4957 8188
rect 4957 8132 5013 8188
rect 5013 8132 5017 8188
rect 4953 8128 5017 8132
rect 5033 8188 5097 8192
rect 5033 8132 5037 8188
rect 5037 8132 5093 8188
rect 5093 8132 5097 8188
rect 5033 8128 5097 8132
rect 5113 8188 5177 8192
rect 5113 8132 5117 8188
rect 5117 8132 5173 8188
rect 5173 8132 5177 8188
rect 5113 8128 5177 8132
rect 12715 8188 12779 8192
rect 12715 8132 12719 8188
rect 12719 8132 12775 8188
rect 12775 8132 12779 8188
rect 12715 8128 12779 8132
rect 12795 8188 12859 8192
rect 12795 8132 12799 8188
rect 12799 8132 12855 8188
rect 12855 8132 12859 8188
rect 12795 8128 12859 8132
rect 12875 8188 12939 8192
rect 12875 8132 12879 8188
rect 12879 8132 12935 8188
rect 12935 8132 12939 8188
rect 12875 8128 12939 8132
rect 12955 8188 13019 8192
rect 12955 8132 12959 8188
rect 12959 8132 13015 8188
rect 13015 8132 13019 8188
rect 12955 8128 13019 8132
rect 20557 8188 20621 8192
rect 20557 8132 20561 8188
rect 20561 8132 20617 8188
rect 20617 8132 20621 8188
rect 20557 8128 20621 8132
rect 20637 8188 20701 8192
rect 20637 8132 20641 8188
rect 20641 8132 20697 8188
rect 20697 8132 20701 8188
rect 20637 8128 20701 8132
rect 20717 8188 20781 8192
rect 20717 8132 20721 8188
rect 20721 8132 20777 8188
rect 20777 8132 20781 8188
rect 20717 8128 20781 8132
rect 20797 8188 20861 8192
rect 20797 8132 20801 8188
rect 20801 8132 20857 8188
rect 20857 8132 20861 8188
rect 20797 8128 20861 8132
rect 28399 8188 28463 8192
rect 28399 8132 28403 8188
rect 28403 8132 28459 8188
rect 28459 8132 28463 8188
rect 28399 8128 28463 8132
rect 28479 8188 28543 8192
rect 28479 8132 28483 8188
rect 28483 8132 28539 8188
rect 28539 8132 28543 8188
rect 28479 8128 28543 8132
rect 28559 8188 28623 8192
rect 28559 8132 28563 8188
rect 28563 8132 28619 8188
rect 28619 8132 28623 8188
rect 28559 8128 28623 8132
rect 28639 8188 28703 8192
rect 28639 8132 28643 8188
rect 28643 8132 28699 8188
rect 28699 8132 28703 8188
rect 28639 8128 28703 8132
rect 8794 7644 8858 7648
rect 8794 7588 8798 7644
rect 8798 7588 8854 7644
rect 8854 7588 8858 7644
rect 8794 7584 8858 7588
rect 8874 7644 8938 7648
rect 8874 7588 8878 7644
rect 8878 7588 8934 7644
rect 8934 7588 8938 7644
rect 8874 7584 8938 7588
rect 8954 7644 9018 7648
rect 8954 7588 8958 7644
rect 8958 7588 9014 7644
rect 9014 7588 9018 7644
rect 8954 7584 9018 7588
rect 9034 7644 9098 7648
rect 9034 7588 9038 7644
rect 9038 7588 9094 7644
rect 9094 7588 9098 7644
rect 9034 7584 9098 7588
rect 16636 7644 16700 7648
rect 16636 7588 16640 7644
rect 16640 7588 16696 7644
rect 16696 7588 16700 7644
rect 16636 7584 16700 7588
rect 16716 7644 16780 7648
rect 16716 7588 16720 7644
rect 16720 7588 16776 7644
rect 16776 7588 16780 7644
rect 16716 7584 16780 7588
rect 16796 7644 16860 7648
rect 16796 7588 16800 7644
rect 16800 7588 16856 7644
rect 16856 7588 16860 7644
rect 16796 7584 16860 7588
rect 16876 7644 16940 7648
rect 16876 7588 16880 7644
rect 16880 7588 16936 7644
rect 16936 7588 16940 7644
rect 16876 7584 16940 7588
rect 24478 7644 24542 7648
rect 24478 7588 24482 7644
rect 24482 7588 24538 7644
rect 24538 7588 24542 7644
rect 24478 7584 24542 7588
rect 24558 7644 24622 7648
rect 24558 7588 24562 7644
rect 24562 7588 24618 7644
rect 24618 7588 24622 7644
rect 24558 7584 24622 7588
rect 24638 7644 24702 7648
rect 24638 7588 24642 7644
rect 24642 7588 24698 7644
rect 24698 7588 24702 7644
rect 24638 7584 24702 7588
rect 24718 7644 24782 7648
rect 24718 7588 24722 7644
rect 24722 7588 24778 7644
rect 24778 7588 24782 7644
rect 24718 7584 24782 7588
rect 32320 7644 32384 7648
rect 32320 7588 32324 7644
rect 32324 7588 32380 7644
rect 32380 7588 32384 7644
rect 32320 7584 32384 7588
rect 32400 7644 32464 7648
rect 32400 7588 32404 7644
rect 32404 7588 32460 7644
rect 32460 7588 32464 7644
rect 32400 7584 32464 7588
rect 32480 7644 32544 7648
rect 32480 7588 32484 7644
rect 32484 7588 32540 7644
rect 32540 7588 32544 7644
rect 32480 7584 32544 7588
rect 32560 7644 32624 7648
rect 32560 7588 32564 7644
rect 32564 7588 32620 7644
rect 32620 7588 32624 7644
rect 32560 7584 32624 7588
rect 4873 7100 4937 7104
rect 4873 7044 4877 7100
rect 4877 7044 4933 7100
rect 4933 7044 4937 7100
rect 4873 7040 4937 7044
rect 4953 7100 5017 7104
rect 4953 7044 4957 7100
rect 4957 7044 5013 7100
rect 5013 7044 5017 7100
rect 4953 7040 5017 7044
rect 5033 7100 5097 7104
rect 5033 7044 5037 7100
rect 5037 7044 5093 7100
rect 5093 7044 5097 7100
rect 5033 7040 5097 7044
rect 5113 7100 5177 7104
rect 5113 7044 5117 7100
rect 5117 7044 5173 7100
rect 5173 7044 5177 7100
rect 5113 7040 5177 7044
rect 12715 7100 12779 7104
rect 12715 7044 12719 7100
rect 12719 7044 12775 7100
rect 12775 7044 12779 7100
rect 12715 7040 12779 7044
rect 12795 7100 12859 7104
rect 12795 7044 12799 7100
rect 12799 7044 12855 7100
rect 12855 7044 12859 7100
rect 12795 7040 12859 7044
rect 12875 7100 12939 7104
rect 12875 7044 12879 7100
rect 12879 7044 12935 7100
rect 12935 7044 12939 7100
rect 12875 7040 12939 7044
rect 12955 7100 13019 7104
rect 12955 7044 12959 7100
rect 12959 7044 13015 7100
rect 13015 7044 13019 7100
rect 12955 7040 13019 7044
rect 20557 7100 20621 7104
rect 20557 7044 20561 7100
rect 20561 7044 20617 7100
rect 20617 7044 20621 7100
rect 20557 7040 20621 7044
rect 20637 7100 20701 7104
rect 20637 7044 20641 7100
rect 20641 7044 20697 7100
rect 20697 7044 20701 7100
rect 20637 7040 20701 7044
rect 20717 7100 20781 7104
rect 20717 7044 20721 7100
rect 20721 7044 20777 7100
rect 20777 7044 20781 7100
rect 20717 7040 20781 7044
rect 20797 7100 20861 7104
rect 20797 7044 20801 7100
rect 20801 7044 20857 7100
rect 20857 7044 20861 7100
rect 20797 7040 20861 7044
rect 28399 7100 28463 7104
rect 28399 7044 28403 7100
rect 28403 7044 28459 7100
rect 28459 7044 28463 7100
rect 28399 7040 28463 7044
rect 28479 7100 28543 7104
rect 28479 7044 28483 7100
rect 28483 7044 28539 7100
rect 28539 7044 28543 7100
rect 28479 7040 28543 7044
rect 28559 7100 28623 7104
rect 28559 7044 28563 7100
rect 28563 7044 28619 7100
rect 28619 7044 28623 7100
rect 28559 7040 28623 7044
rect 28639 7100 28703 7104
rect 28639 7044 28643 7100
rect 28643 7044 28699 7100
rect 28699 7044 28703 7100
rect 28639 7040 28703 7044
rect 8794 6556 8858 6560
rect 8794 6500 8798 6556
rect 8798 6500 8854 6556
rect 8854 6500 8858 6556
rect 8794 6496 8858 6500
rect 8874 6556 8938 6560
rect 8874 6500 8878 6556
rect 8878 6500 8934 6556
rect 8934 6500 8938 6556
rect 8874 6496 8938 6500
rect 8954 6556 9018 6560
rect 8954 6500 8958 6556
rect 8958 6500 9014 6556
rect 9014 6500 9018 6556
rect 8954 6496 9018 6500
rect 9034 6556 9098 6560
rect 9034 6500 9038 6556
rect 9038 6500 9094 6556
rect 9094 6500 9098 6556
rect 9034 6496 9098 6500
rect 16636 6556 16700 6560
rect 16636 6500 16640 6556
rect 16640 6500 16696 6556
rect 16696 6500 16700 6556
rect 16636 6496 16700 6500
rect 16716 6556 16780 6560
rect 16716 6500 16720 6556
rect 16720 6500 16776 6556
rect 16776 6500 16780 6556
rect 16716 6496 16780 6500
rect 16796 6556 16860 6560
rect 16796 6500 16800 6556
rect 16800 6500 16856 6556
rect 16856 6500 16860 6556
rect 16796 6496 16860 6500
rect 16876 6556 16940 6560
rect 16876 6500 16880 6556
rect 16880 6500 16936 6556
rect 16936 6500 16940 6556
rect 16876 6496 16940 6500
rect 24478 6556 24542 6560
rect 24478 6500 24482 6556
rect 24482 6500 24538 6556
rect 24538 6500 24542 6556
rect 24478 6496 24542 6500
rect 24558 6556 24622 6560
rect 24558 6500 24562 6556
rect 24562 6500 24618 6556
rect 24618 6500 24622 6556
rect 24558 6496 24622 6500
rect 24638 6556 24702 6560
rect 24638 6500 24642 6556
rect 24642 6500 24698 6556
rect 24698 6500 24702 6556
rect 24638 6496 24702 6500
rect 24718 6556 24782 6560
rect 24718 6500 24722 6556
rect 24722 6500 24778 6556
rect 24778 6500 24782 6556
rect 24718 6496 24782 6500
rect 32320 6556 32384 6560
rect 32320 6500 32324 6556
rect 32324 6500 32380 6556
rect 32380 6500 32384 6556
rect 32320 6496 32384 6500
rect 32400 6556 32464 6560
rect 32400 6500 32404 6556
rect 32404 6500 32460 6556
rect 32460 6500 32464 6556
rect 32400 6496 32464 6500
rect 32480 6556 32544 6560
rect 32480 6500 32484 6556
rect 32484 6500 32540 6556
rect 32540 6500 32544 6556
rect 32480 6496 32544 6500
rect 32560 6556 32624 6560
rect 32560 6500 32564 6556
rect 32564 6500 32620 6556
rect 32620 6500 32624 6556
rect 32560 6496 32624 6500
rect 4873 6012 4937 6016
rect 4873 5956 4877 6012
rect 4877 5956 4933 6012
rect 4933 5956 4937 6012
rect 4873 5952 4937 5956
rect 4953 6012 5017 6016
rect 4953 5956 4957 6012
rect 4957 5956 5013 6012
rect 5013 5956 5017 6012
rect 4953 5952 5017 5956
rect 5033 6012 5097 6016
rect 5033 5956 5037 6012
rect 5037 5956 5093 6012
rect 5093 5956 5097 6012
rect 5033 5952 5097 5956
rect 5113 6012 5177 6016
rect 5113 5956 5117 6012
rect 5117 5956 5173 6012
rect 5173 5956 5177 6012
rect 5113 5952 5177 5956
rect 12715 6012 12779 6016
rect 12715 5956 12719 6012
rect 12719 5956 12775 6012
rect 12775 5956 12779 6012
rect 12715 5952 12779 5956
rect 12795 6012 12859 6016
rect 12795 5956 12799 6012
rect 12799 5956 12855 6012
rect 12855 5956 12859 6012
rect 12795 5952 12859 5956
rect 12875 6012 12939 6016
rect 12875 5956 12879 6012
rect 12879 5956 12935 6012
rect 12935 5956 12939 6012
rect 12875 5952 12939 5956
rect 12955 6012 13019 6016
rect 12955 5956 12959 6012
rect 12959 5956 13015 6012
rect 13015 5956 13019 6012
rect 12955 5952 13019 5956
rect 20557 6012 20621 6016
rect 20557 5956 20561 6012
rect 20561 5956 20617 6012
rect 20617 5956 20621 6012
rect 20557 5952 20621 5956
rect 20637 6012 20701 6016
rect 20637 5956 20641 6012
rect 20641 5956 20697 6012
rect 20697 5956 20701 6012
rect 20637 5952 20701 5956
rect 20717 6012 20781 6016
rect 20717 5956 20721 6012
rect 20721 5956 20777 6012
rect 20777 5956 20781 6012
rect 20717 5952 20781 5956
rect 20797 6012 20861 6016
rect 20797 5956 20801 6012
rect 20801 5956 20857 6012
rect 20857 5956 20861 6012
rect 20797 5952 20861 5956
rect 28399 6012 28463 6016
rect 28399 5956 28403 6012
rect 28403 5956 28459 6012
rect 28459 5956 28463 6012
rect 28399 5952 28463 5956
rect 28479 6012 28543 6016
rect 28479 5956 28483 6012
rect 28483 5956 28539 6012
rect 28539 5956 28543 6012
rect 28479 5952 28543 5956
rect 28559 6012 28623 6016
rect 28559 5956 28563 6012
rect 28563 5956 28619 6012
rect 28619 5956 28623 6012
rect 28559 5952 28623 5956
rect 28639 6012 28703 6016
rect 28639 5956 28643 6012
rect 28643 5956 28699 6012
rect 28699 5956 28703 6012
rect 28639 5952 28703 5956
rect 8794 5468 8858 5472
rect 8794 5412 8798 5468
rect 8798 5412 8854 5468
rect 8854 5412 8858 5468
rect 8794 5408 8858 5412
rect 8874 5468 8938 5472
rect 8874 5412 8878 5468
rect 8878 5412 8934 5468
rect 8934 5412 8938 5468
rect 8874 5408 8938 5412
rect 8954 5468 9018 5472
rect 8954 5412 8958 5468
rect 8958 5412 9014 5468
rect 9014 5412 9018 5468
rect 8954 5408 9018 5412
rect 9034 5468 9098 5472
rect 9034 5412 9038 5468
rect 9038 5412 9094 5468
rect 9094 5412 9098 5468
rect 9034 5408 9098 5412
rect 16636 5468 16700 5472
rect 16636 5412 16640 5468
rect 16640 5412 16696 5468
rect 16696 5412 16700 5468
rect 16636 5408 16700 5412
rect 16716 5468 16780 5472
rect 16716 5412 16720 5468
rect 16720 5412 16776 5468
rect 16776 5412 16780 5468
rect 16716 5408 16780 5412
rect 16796 5468 16860 5472
rect 16796 5412 16800 5468
rect 16800 5412 16856 5468
rect 16856 5412 16860 5468
rect 16796 5408 16860 5412
rect 16876 5468 16940 5472
rect 16876 5412 16880 5468
rect 16880 5412 16936 5468
rect 16936 5412 16940 5468
rect 16876 5408 16940 5412
rect 24478 5468 24542 5472
rect 24478 5412 24482 5468
rect 24482 5412 24538 5468
rect 24538 5412 24542 5468
rect 24478 5408 24542 5412
rect 24558 5468 24622 5472
rect 24558 5412 24562 5468
rect 24562 5412 24618 5468
rect 24618 5412 24622 5468
rect 24558 5408 24622 5412
rect 24638 5468 24702 5472
rect 24638 5412 24642 5468
rect 24642 5412 24698 5468
rect 24698 5412 24702 5468
rect 24638 5408 24702 5412
rect 24718 5468 24782 5472
rect 24718 5412 24722 5468
rect 24722 5412 24778 5468
rect 24778 5412 24782 5468
rect 24718 5408 24782 5412
rect 32320 5468 32384 5472
rect 32320 5412 32324 5468
rect 32324 5412 32380 5468
rect 32380 5412 32384 5468
rect 32320 5408 32384 5412
rect 32400 5468 32464 5472
rect 32400 5412 32404 5468
rect 32404 5412 32460 5468
rect 32460 5412 32464 5468
rect 32400 5408 32464 5412
rect 32480 5468 32544 5472
rect 32480 5412 32484 5468
rect 32484 5412 32540 5468
rect 32540 5412 32544 5468
rect 32480 5408 32544 5412
rect 32560 5468 32624 5472
rect 32560 5412 32564 5468
rect 32564 5412 32620 5468
rect 32620 5412 32624 5468
rect 32560 5408 32624 5412
rect 4873 4924 4937 4928
rect 4873 4868 4877 4924
rect 4877 4868 4933 4924
rect 4933 4868 4937 4924
rect 4873 4864 4937 4868
rect 4953 4924 5017 4928
rect 4953 4868 4957 4924
rect 4957 4868 5013 4924
rect 5013 4868 5017 4924
rect 4953 4864 5017 4868
rect 5033 4924 5097 4928
rect 5033 4868 5037 4924
rect 5037 4868 5093 4924
rect 5093 4868 5097 4924
rect 5033 4864 5097 4868
rect 5113 4924 5177 4928
rect 5113 4868 5117 4924
rect 5117 4868 5173 4924
rect 5173 4868 5177 4924
rect 5113 4864 5177 4868
rect 12715 4924 12779 4928
rect 12715 4868 12719 4924
rect 12719 4868 12775 4924
rect 12775 4868 12779 4924
rect 12715 4864 12779 4868
rect 12795 4924 12859 4928
rect 12795 4868 12799 4924
rect 12799 4868 12855 4924
rect 12855 4868 12859 4924
rect 12795 4864 12859 4868
rect 12875 4924 12939 4928
rect 12875 4868 12879 4924
rect 12879 4868 12935 4924
rect 12935 4868 12939 4924
rect 12875 4864 12939 4868
rect 12955 4924 13019 4928
rect 12955 4868 12959 4924
rect 12959 4868 13015 4924
rect 13015 4868 13019 4924
rect 12955 4864 13019 4868
rect 20557 4924 20621 4928
rect 20557 4868 20561 4924
rect 20561 4868 20617 4924
rect 20617 4868 20621 4924
rect 20557 4864 20621 4868
rect 20637 4924 20701 4928
rect 20637 4868 20641 4924
rect 20641 4868 20697 4924
rect 20697 4868 20701 4924
rect 20637 4864 20701 4868
rect 20717 4924 20781 4928
rect 20717 4868 20721 4924
rect 20721 4868 20777 4924
rect 20777 4868 20781 4924
rect 20717 4864 20781 4868
rect 20797 4924 20861 4928
rect 20797 4868 20801 4924
rect 20801 4868 20857 4924
rect 20857 4868 20861 4924
rect 20797 4864 20861 4868
rect 28399 4924 28463 4928
rect 28399 4868 28403 4924
rect 28403 4868 28459 4924
rect 28459 4868 28463 4924
rect 28399 4864 28463 4868
rect 28479 4924 28543 4928
rect 28479 4868 28483 4924
rect 28483 4868 28539 4924
rect 28539 4868 28543 4924
rect 28479 4864 28543 4868
rect 28559 4924 28623 4928
rect 28559 4868 28563 4924
rect 28563 4868 28619 4924
rect 28619 4868 28623 4924
rect 28559 4864 28623 4868
rect 28639 4924 28703 4928
rect 28639 4868 28643 4924
rect 28643 4868 28699 4924
rect 28699 4868 28703 4924
rect 28639 4864 28703 4868
rect 8794 4380 8858 4384
rect 8794 4324 8798 4380
rect 8798 4324 8854 4380
rect 8854 4324 8858 4380
rect 8794 4320 8858 4324
rect 8874 4380 8938 4384
rect 8874 4324 8878 4380
rect 8878 4324 8934 4380
rect 8934 4324 8938 4380
rect 8874 4320 8938 4324
rect 8954 4380 9018 4384
rect 8954 4324 8958 4380
rect 8958 4324 9014 4380
rect 9014 4324 9018 4380
rect 8954 4320 9018 4324
rect 9034 4380 9098 4384
rect 9034 4324 9038 4380
rect 9038 4324 9094 4380
rect 9094 4324 9098 4380
rect 9034 4320 9098 4324
rect 16636 4380 16700 4384
rect 16636 4324 16640 4380
rect 16640 4324 16696 4380
rect 16696 4324 16700 4380
rect 16636 4320 16700 4324
rect 16716 4380 16780 4384
rect 16716 4324 16720 4380
rect 16720 4324 16776 4380
rect 16776 4324 16780 4380
rect 16716 4320 16780 4324
rect 16796 4380 16860 4384
rect 16796 4324 16800 4380
rect 16800 4324 16856 4380
rect 16856 4324 16860 4380
rect 16796 4320 16860 4324
rect 16876 4380 16940 4384
rect 16876 4324 16880 4380
rect 16880 4324 16936 4380
rect 16936 4324 16940 4380
rect 16876 4320 16940 4324
rect 24478 4380 24542 4384
rect 24478 4324 24482 4380
rect 24482 4324 24538 4380
rect 24538 4324 24542 4380
rect 24478 4320 24542 4324
rect 24558 4380 24622 4384
rect 24558 4324 24562 4380
rect 24562 4324 24618 4380
rect 24618 4324 24622 4380
rect 24558 4320 24622 4324
rect 24638 4380 24702 4384
rect 24638 4324 24642 4380
rect 24642 4324 24698 4380
rect 24698 4324 24702 4380
rect 24638 4320 24702 4324
rect 24718 4380 24782 4384
rect 24718 4324 24722 4380
rect 24722 4324 24778 4380
rect 24778 4324 24782 4380
rect 24718 4320 24782 4324
rect 32320 4380 32384 4384
rect 32320 4324 32324 4380
rect 32324 4324 32380 4380
rect 32380 4324 32384 4380
rect 32320 4320 32384 4324
rect 32400 4380 32464 4384
rect 32400 4324 32404 4380
rect 32404 4324 32460 4380
rect 32460 4324 32464 4380
rect 32400 4320 32464 4324
rect 32480 4380 32544 4384
rect 32480 4324 32484 4380
rect 32484 4324 32540 4380
rect 32540 4324 32544 4380
rect 32480 4320 32544 4324
rect 32560 4380 32624 4384
rect 32560 4324 32564 4380
rect 32564 4324 32620 4380
rect 32620 4324 32624 4380
rect 32560 4320 32624 4324
rect 4873 3836 4937 3840
rect 4873 3780 4877 3836
rect 4877 3780 4933 3836
rect 4933 3780 4937 3836
rect 4873 3776 4937 3780
rect 4953 3836 5017 3840
rect 4953 3780 4957 3836
rect 4957 3780 5013 3836
rect 5013 3780 5017 3836
rect 4953 3776 5017 3780
rect 5033 3836 5097 3840
rect 5033 3780 5037 3836
rect 5037 3780 5093 3836
rect 5093 3780 5097 3836
rect 5033 3776 5097 3780
rect 5113 3836 5177 3840
rect 5113 3780 5117 3836
rect 5117 3780 5173 3836
rect 5173 3780 5177 3836
rect 5113 3776 5177 3780
rect 12715 3836 12779 3840
rect 12715 3780 12719 3836
rect 12719 3780 12775 3836
rect 12775 3780 12779 3836
rect 12715 3776 12779 3780
rect 12795 3836 12859 3840
rect 12795 3780 12799 3836
rect 12799 3780 12855 3836
rect 12855 3780 12859 3836
rect 12795 3776 12859 3780
rect 12875 3836 12939 3840
rect 12875 3780 12879 3836
rect 12879 3780 12935 3836
rect 12935 3780 12939 3836
rect 12875 3776 12939 3780
rect 12955 3836 13019 3840
rect 12955 3780 12959 3836
rect 12959 3780 13015 3836
rect 13015 3780 13019 3836
rect 12955 3776 13019 3780
rect 20557 3836 20621 3840
rect 20557 3780 20561 3836
rect 20561 3780 20617 3836
rect 20617 3780 20621 3836
rect 20557 3776 20621 3780
rect 20637 3836 20701 3840
rect 20637 3780 20641 3836
rect 20641 3780 20697 3836
rect 20697 3780 20701 3836
rect 20637 3776 20701 3780
rect 20717 3836 20781 3840
rect 20717 3780 20721 3836
rect 20721 3780 20777 3836
rect 20777 3780 20781 3836
rect 20717 3776 20781 3780
rect 20797 3836 20861 3840
rect 20797 3780 20801 3836
rect 20801 3780 20857 3836
rect 20857 3780 20861 3836
rect 20797 3776 20861 3780
rect 28399 3836 28463 3840
rect 28399 3780 28403 3836
rect 28403 3780 28459 3836
rect 28459 3780 28463 3836
rect 28399 3776 28463 3780
rect 28479 3836 28543 3840
rect 28479 3780 28483 3836
rect 28483 3780 28539 3836
rect 28539 3780 28543 3836
rect 28479 3776 28543 3780
rect 28559 3836 28623 3840
rect 28559 3780 28563 3836
rect 28563 3780 28619 3836
rect 28619 3780 28623 3836
rect 28559 3776 28623 3780
rect 28639 3836 28703 3840
rect 28639 3780 28643 3836
rect 28643 3780 28699 3836
rect 28699 3780 28703 3836
rect 28639 3776 28703 3780
rect 8794 3292 8858 3296
rect 8794 3236 8798 3292
rect 8798 3236 8854 3292
rect 8854 3236 8858 3292
rect 8794 3232 8858 3236
rect 8874 3292 8938 3296
rect 8874 3236 8878 3292
rect 8878 3236 8934 3292
rect 8934 3236 8938 3292
rect 8874 3232 8938 3236
rect 8954 3292 9018 3296
rect 8954 3236 8958 3292
rect 8958 3236 9014 3292
rect 9014 3236 9018 3292
rect 8954 3232 9018 3236
rect 9034 3292 9098 3296
rect 9034 3236 9038 3292
rect 9038 3236 9094 3292
rect 9094 3236 9098 3292
rect 9034 3232 9098 3236
rect 16636 3292 16700 3296
rect 16636 3236 16640 3292
rect 16640 3236 16696 3292
rect 16696 3236 16700 3292
rect 16636 3232 16700 3236
rect 16716 3292 16780 3296
rect 16716 3236 16720 3292
rect 16720 3236 16776 3292
rect 16776 3236 16780 3292
rect 16716 3232 16780 3236
rect 16796 3292 16860 3296
rect 16796 3236 16800 3292
rect 16800 3236 16856 3292
rect 16856 3236 16860 3292
rect 16796 3232 16860 3236
rect 16876 3292 16940 3296
rect 16876 3236 16880 3292
rect 16880 3236 16936 3292
rect 16936 3236 16940 3292
rect 16876 3232 16940 3236
rect 24478 3292 24542 3296
rect 24478 3236 24482 3292
rect 24482 3236 24538 3292
rect 24538 3236 24542 3292
rect 24478 3232 24542 3236
rect 24558 3292 24622 3296
rect 24558 3236 24562 3292
rect 24562 3236 24618 3292
rect 24618 3236 24622 3292
rect 24558 3232 24622 3236
rect 24638 3292 24702 3296
rect 24638 3236 24642 3292
rect 24642 3236 24698 3292
rect 24698 3236 24702 3292
rect 24638 3232 24702 3236
rect 24718 3292 24782 3296
rect 24718 3236 24722 3292
rect 24722 3236 24778 3292
rect 24778 3236 24782 3292
rect 24718 3232 24782 3236
rect 32320 3292 32384 3296
rect 32320 3236 32324 3292
rect 32324 3236 32380 3292
rect 32380 3236 32384 3292
rect 32320 3232 32384 3236
rect 32400 3292 32464 3296
rect 32400 3236 32404 3292
rect 32404 3236 32460 3292
rect 32460 3236 32464 3292
rect 32400 3232 32464 3236
rect 32480 3292 32544 3296
rect 32480 3236 32484 3292
rect 32484 3236 32540 3292
rect 32540 3236 32544 3292
rect 32480 3232 32544 3236
rect 32560 3292 32624 3296
rect 32560 3236 32564 3292
rect 32564 3236 32620 3292
rect 32620 3236 32624 3292
rect 32560 3232 32624 3236
rect 4873 2748 4937 2752
rect 4873 2692 4877 2748
rect 4877 2692 4933 2748
rect 4933 2692 4937 2748
rect 4873 2688 4937 2692
rect 4953 2748 5017 2752
rect 4953 2692 4957 2748
rect 4957 2692 5013 2748
rect 5013 2692 5017 2748
rect 4953 2688 5017 2692
rect 5033 2748 5097 2752
rect 5033 2692 5037 2748
rect 5037 2692 5093 2748
rect 5093 2692 5097 2748
rect 5033 2688 5097 2692
rect 5113 2748 5177 2752
rect 5113 2692 5117 2748
rect 5117 2692 5173 2748
rect 5173 2692 5177 2748
rect 5113 2688 5177 2692
rect 12715 2748 12779 2752
rect 12715 2692 12719 2748
rect 12719 2692 12775 2748
rect 12775 2692 12779 2748
rect 12715 2688 12779 2692
rect 12795 2748 12859 2752
rect 12795 2692 12799 2748
rect 12799 2692 12855 2748
rect 12855 2692 12859 2748
rect 12795 2688 12859 2692
rect 12875 2748 12939 2752
rect 12875 2692 12879 2748
rect 12879 2692 12935 2748
rect 12935 2692 12939 2748
rect 12875 2688 12939 2692
rect 12955 2748 13019 2752
rect 12955 2692 12959 2748
rect 12959 2692 13015 2748
rect 13015 2692 13019 2748
rect 12955 2688 13019 2692
rect 20557 2748 20621 2752
rect 20557 2692 20561 2748
rect 20561 2692 20617 2748
rect 20617 2692 20621 2748
rect 20557 2688 20621 2692
rect 20637 2748 20701 2752
rect 20637 2692 20641 2748
rect 20641 2692 20697 2748
rect 20697 2692 20701 2748
rect 20637 2688 20701 2692
rect 20717 2748 20781 2752
rect 20717 2692 20721 2748
rect 20721 2692 20777 2748
rect 20777 2692 20781 2748
rect 20717 2688 20781 2692
rect 20797 2748 20861 2752
rect 20797 2692 20801 2748
rect 20801 2692 20857 2748
rect 20857 2692 20861 2748
rect 20797 2688 20861 2692
rect 28399 2748 28463 2752
rect 28399 2692 28403 2748
rect 28403 2692 28459 2748
rect 28459 2692 28463 2748
rect 28399 2688 28463 2692
rect 28479 2748 28543 2752
rect 28479 2692 28483 2748
rect 28483 2692 28539 2748
rect 28539 2692 28543 2748
rect 28479 2688 28543 2692
rect 28559 2748 28623 2752
rect 28559 2692 28563 2748
rect 28563 2692 28619 2748
rect 28619 2692 28623 2748
rect 28559 2688 28623 2692
rect 28639 2748 28703 2752
rect 28639 2692 28643 2748
rect 28643 2692 28699 2748
rect 28699 2692 28703 2748
rect 28639 2688 28703 2692
rect 8794 2204 8858 2208
rect 8794 2148 8798 2204
rect 8798 2148 8854 2204
rect 8854 2148 8858 2204
rect 8794 2144 8858 2148
rect 8874 2204 8938 2208
rect 8874 2148 8878 2204
rect 8878 2148 8934 2204
rect 8934 2148 8938 2204
rect 8874 2144 8938 2148
rect 8954 2204 9018 2208
rect 8954 2148 8958 2204
rect 8958 2148 9014 2204
rect 9014 2148 9018 2204
rect 8954 2144 9018 2148
rect 9034 2204 9098 2208
rect 9034 2148 9038 2204
rect 9038 2148 9094 2204
rect 9094 2148 9098 2204
rect 9034 2144 9098 2148
rect 16636 2204 16700 2208
rect 16636 2148 16640 2204
rect 16640 2148 16696 2204
rect 16696 2148 16700 2204
rect 16636 2144 16700 2148
rect 16716 2204 16780 2208
rect 16716 2148 16720 2204
rect 16720 2148 16776 2204
rect 16776 2148 16780 2204
rect 16716 2144 16780 2148
rect 16796 2204 16860 2208
rect 16796 2148 16800 2204
rect 16800 2148 16856 2204
rect 16856 2148 16860 2204
rect 16796 2144 16860 2148
rect 16876 2204 16940 2208
rect 16876 2148 16880 2204
rect 16880 2148 16936 2204
rect 16936 2148 16940 2204
rect 16876 2144 16940 2148
rect 24478 2204 24542 2208
rect 24478 2148 24482 2204
rect 24482 2148 24538 2204
rect 24538 2148 24542 2204
rect 24478 2144 24542 2148
rect 24558 2204 24622 2208
rect 24558 2148 24562 2204
rect 24562 2148 24618 2204
rect 24618 2148 24622 2204
rect 24558 2144 24622 2148
rect 24638 2204 24702 2208
rect 24638 2148 24642 2204
rect 24642 2148 24698 2204
rect 24698 2148 24702 2204
rect 24638 2144 24702 2148
rect 24718 2204 24782 2208
rect 24718 2148 24722 2204
rect 24722 2148 24778 2204
rect 24778 2148 24782 2204
rect 24718 2144 24782 2148
rect 32320 2204 32384 2208
rect 32320 2148 32324 2204
rect 32324 2148 32380 2204
rect 32380 2148 32384 2204
rect 32320 2144 32384 2148
rect 32400 2204 32464 2208
rect 32400 2148 32404 2204
rect 32404 2148 32460 2204
rect 32460 2148 32464 2204
rect 32400 2144 32464 2148
rect 32480 2204 32544 2208
rect 32480 2148 32484 2204
rect 32484 2148 32540 2204
rect 32540 2148 32544 2204
rect 32480 2144 32544 2148
rect 32560 2204 32624 2208
rect 32560 2148 32564 2204
rect 32564 2148 32620 2204
rect 32620 2148 32624 2204
rect 32560 2144 32624 2148
rect 4873 1660 4937 1664
rect 4873 1604 4877 1660
rect 4877 1604 4933 1660
rect 4933 1604 4937 1660
rect 4873 1600 4937 1604
rect 4953 1660 5017 1664
rect 4953 1604 4957 1660
rect 4957 1604 5013 1660
rect 5013 1604 5017 1660
rect 4953 1600 5017 1604
rect 5033 1660 5097 1664
rect 5033 1604 5037 1660
rect 5037 1604 5093 1660
rect 5093 1604 5097 1660
rect 5033 1600 5097 1604
rect 5113 1660 5177 1664
rect 5113 1604 5117 1660
rect 5117 1604 5173 1660
rect 5173 1604 5177 1660
rect 5113 1600 5177 1604
rect 12715 1660 12779 1664
rect 12715 1604 12719 1660
rect 12719 1604 12775 1660
rect 12775 1604 12779 1660
rect 12715 1600 12779 1604
rect 12795 1660 12859 1664
rect 12795 1604 12799 1660
rect 12799 1604 12855 1660
rect 12855 1604 12859 1660
rect 12795 1600 12859 1604
rect 12875 1660 12939 1664
rect 12875 1604 12879 1660
rect 12879 1604 12935 1660
rect 12935 1604 12939 1660
rect 12875 1600 12939 1604
rect 12955 1660 13019 1664
rect 12955 1604 12959 1660
rect 12959 1604 13015 1660
rect 13015 1604 13019 1660
rect 12955 1600 13019 1604
rect 20557 1660 20621 1664
rect 20557 1604 20561 1660
rect 20561 1604 20617 1660
rect 20617 1604 20621 1660
rect 20557 1600 20621 1604
rect 20637 1660 20701 1664
rect 20637 1604 20641 1660
rect 20641 1604 20697 1660
rect 20697 1604 20701 1660
rect 20637 1600 20701 1604
rect 20717 1660 20781 1664
rect 20717 1604 20721 1660
rect 20721 1604 20777 1660
rect 20777 1604 20781 1660
rect 20717 1600 20781 1604
rect 20797 1660 20861 1664
rect 20797 1604 20801 1660
rect 20801 1604 20857 1660
rect 20857 1604 20861 1660
rect 20797 1600 20861 1604
rect 28399 1660 28463 1664
rect 28399 1604 28403 1660
rect 28403 1604 28459 1660
rect 28459 1604 28463 1660
rect 28399 1600 28463 1604
rect 28479 1660 28543 1664
rect 28479 1604 28483 1660
rect 28483 1604 28539 1660
rect 28539 1604 28543 1660
rect 28479 1600 28543 1604
rect 28559 1660 28623 1664
rect 28559 1604 28563 1660
rect 28563 1604 28619 1660
rect 28619 1604 28623 1660
rect 28559 1600 28623 1604
rect 28639 1660 28703 1664
rect 28639 1604 28643 1660
rect 28643 1604 28699 1660
rect 28699 1604 28703 1660
rect 28639 1600 28703 1604
rect 8794 1116 8858 1120
rect 8794 1060 8798 1116
rect 8798 1060 8854 1116
rect 8854 1060 8858 1116
rect 8794 1056 8858 1060
rect 8874 1116 8938 1120
rect 8874 1060 8878 1116
rect 8878 1060 8934 1116
rect 8934 1060 8938 1116
rect 8874 1056 8938 1060
rect 8954 1116 9018 1120
rect 8954 1060 8958 1116
rect 8958 1060 9014 1116
rect 9014 1060 9018 1116
rect 8954 1056 9018 1060
rect 9034 1116 9098 1120
rect 9034 1060 9038 1116
rect 9038 1060 9094 1116
rect 9094 1060 9098 1116
rect 9034 1056 9098 1060
rect 16636 1116 16700 1120
rect 16636 1060 16640 1116
rect 16640 1060 16696 1116
rect 16696 1060 16700 1116
rect 16636 1056 16700 1060
rect 16716 1116 16780 1120
rect 16716 1060 16720 1116
rect 16720 1060 16776 1116
rect 16776 1060 16780 1116
rect 16716 1056 16780 1060
rect 16796 1116 16860 1120
rect 16796 1060 16800 1116
rect 16800 1060 16856 1116
rect 16856 1060 16860 1116
rect 16796 1056 16860 1060
rect 16876 1116 16940 1120
rect 16876 1060 16880 1116
rect 16880 1060 16936 1116
rect 16936 1060 16940 1116
rect 16876 1056 16940 1060
rect 24478 1116 24542 1120
rect 24478 1060 24482 1116
rect 24482 1060 24538 1116
rect 24538 1060 24542 1116
rect 24478 1056 24542 1060
rect 24558 1116 24622 1120
rect 24558 1060 24562 1116
rect 24562 1060 24618 1116
rect 24618 1060 24622 1116
rect 24558 1056 24622 1060
rect 24638 1116 24702 1120
rect 24638 1060 24642 1116
rect 24642 1060 24698 1116
rect 24698 1060 24702 1116
rect 24638 1056 24702 1060
rect 24718 1116 24782 1120
rect 24718 1060 24722 1116
rect 24722 1060 24778 1116
rect 24778 1060 24782 1116
rect 24718 1056 24782 1060
rect 32320 1116 32384 1120
rect 32320 1060 32324 1116
rect 32324 1060 32380 1116
rect 32380 1060 32384 1116
rect 32320 1056 32384 1060
rect 32400 1116 32464 1120
rect 32400 1060 32404 1116
rect 32404 1060 32460 1116
rect 32460 1060 32464 1116
rect 32400 1056 32464 1060
rect 32480 1116 32544 1120
rect 32480 1060 32484 1116
rect 32484 1060 32540 1116
rect 32540 1060 32544 1116
rect 32480 1056 32544 1060
rect 32560 1116 32624 1120
rect 32560 1060 32564 1116
rect 32564 1060 32620 1116
rect 32620 1060 32624 1116
rect 32560 1056 32624 1060
<< metal4 >>
rect 1534 19549 1594 21760
rect 2270 20093 2330 21760
rect 3006 20093 3066 21760
rect 2267 20092 2333 20093
rect 2267 20028 2268 20092
rect 2332 20028 2333 20092
rect 2267 20027 2333 20028
rect 3003 20092 3069 20093
rect 3003 20028 3004 20092
rect 3068 20028 3069 20092
rect 3003 20027 3069 20028
rect 3742 19549 3802 21760
rect 4478 20093 4538 21760
rect 5214 20909 5274 21760
rect 5211 20908 5277 20909
rect 5211 20844 5212 20908
rect 5276 20844 5277 20908
rect 5211 20843 5277 20844
rect 4865 20160 5185 20720
rect 4865 20096 4873 20160
rect 4937 20096 4953 20160
rect 5017 20096 5033 20160
rect 5097 20096 5113 20160
rect 5177 20096 5185 20160
rect 4475 20092 4541 20093
rect 4475 20028 4476 20092
rect 4540 20028 4541 20092
rect 4475 20027 4541 20028
rect 1531 19548 1597 19549
rect 1531 19484 1532 19548
rect 1596 19484 1597 19548
rect 1531 19483 1597 19484
rect 3739 19548 3805 19549
rect 3739 19484 3740 19548
rect 3804 19484 3805 19548
rect 3739 19483 3805 19484
rect 4865 19072 5185 20096
rect 5950 20093 6010 21760
rect 6686 20093 6746 21760
rect 5947 20092 6013 20093
rect 5947 20028 5948 20092
rect 6012 20028 6013 20092
rect 5947 20027 6013 20028
rect 6683 20092 6749 20093
rect 6683 20028 6684 20092
rect 6748 20028 6749 20092
rect 6683 20027 6749 20028
rect 7422 19957 7482 21760
rect 8158 20501 8218 21760
rect 8894 20909 8954 21760
rect 8891 20908 8957 20909
rect 8891 20844 8892 20908
rect 8956 20844 8957 20908
rect 8891 20843 8957 20844
rect 8786 20704 9106 20720
rect 8786 20640 8794 20704
rect 8858 20640 8874 20704
rect 8938 20640 8954 20704
rect 9018 20640 9034 20704
rect 9098 20640 9106 20704
rect 8155 20500 8221 20501
rect 8155 20436 8156 20500
rect 8220 20436 8221 20500
rect 8155 20435 8221 20436
rect 7419 19956 7485 19957
rect 7419 19892 7420 19956
rect 7484 19892 7485 19956
rect 7419 19891 7485 19892
rect 4865 19008 4873 19072
rect 4937 19008 4953 19072
rect 5017 19008 5033 19072
rect 5097 19008 5113 19072
rect 5177 19008 5185 19072
rect 4865 17984 5185 19008
rect 4865 17920 4873 17984
rect 4937 17920 4953 17984
rect 5017 17920 5033 17984
rect 5097 17920 5113 17984
rect 5177 17920 5185 17984
rect 4865 16896 5185 17920
rect 4865 16832 4873 16896
rect 4937 16832 4953 16896
rect 5017 16832 5033 16896
rect 5097 16832 5113 16896
rect 5177 16832 5185 16896
rect 4865 15808 5185 16832
rect 4865 15744 4873 15808
rect 4937 15744 4953 15808
rect 5017 15744 5033 15808
rect 5097 15744 5113 15808
rect 5177 15744 5185 15808
rect 4865 14720 5185 15744
rect 4865 14656 4873 14720
rect 4937 14656 4953 14720
rect 5017 14656 5033 14720
rect 5097 14656 5113 14720
rect 5177 14656 5185 14720
rect 4865 13632 5185 14656
rect 4865 13568 4873 13632
rect 4937 13568 4953 13632
rect 5017 13568 5033 13632
rect 5097 13568 5113 13632
rect 5177 13568 5185 13632
rect 4865 12544 5185 13568
rect 4865 12480 4873 12544
rect 4937 12480 4953 12544
rect 5017 12480 5033 12544
rect 5097 12480 5113 12544
rect 5177 12480 5185 12544
rect 4865 11456 5185 12480
rect 4865 11392 4873 11456
rect 4937 11392 4953 11456
rect 5017 11392 5033 11456
rect 5097 11392 5113 11456
rect 5177 11392 5185 11456
rect 4865 10368 5185 11392
rect 4865 10304 4873 10368
rect 4937 10304 4953 10368
rect 5017 10304 5033 10368
rect 5097 10304 5113 10368
rect 5177 10304 5185 10368
rect 4865 9280 5185 10304
rect 4865 9216 4873 9280
rect 4937 9216 4953 9280
rect 5017 9216 5033 9280
rect 5097 9216 5113 9280
rect 5177 9216 5185 9280
rect 4865 8192 5185 9216
rect 4865 8128 4873 8192
rect 4937 8128 4953 8192
rect 5017 8128 5033 8192
rect 5097 8128 5113 8192
rect 5177 8128 5185 8192
rect 4865 7104 5185 8128
rect 4865 7040 4873 7104
rect 4937 7040 4953 7104
rect 5017 7040 5033 7104
rect 5097 7040 5113 7104
rect 5177 7040 5185 7104
rect 4865 6016 5185 7040
rect 4865 5952 4873 6016
rect 4937 5952 4953 6016
rect 5017 5952 5033 6016
rect 5097 5952 5113 6016
rect 5177 5952 5185 6016
rect 4865 4928 5185 5952
rect 4865 4864 4873 4928
rect 4937 4864 4953 4928
rect 5017 4864 5033 4928
rect 5097 4864 5113 4928
rect 5177 4864 5185 4928
rect 4865 3840 5185 4864
rect 4865 3776 4873 3840
rect 4937 3776 4953 3840
rect 5017 3776 5033 3840
rect 5097 3776 5113 3840
rect 5177 3776 5185 3840
rect 4865 2752 5185 3776
rect 4865 2688 4873 2752
rect 4937 2688 4953 2752
rect 5017 2688 5033 2752
rect 5097 2688 5113 2752
rect 5177 2688 5185 2752
rect 4865 1664 5185 2688
rect 4865 1600 4873 1664
rect 4937 1600 4953 1664
rect 5017 1600 5033 1664
rect 5097 1600 5113 1664
rect 5177 1600 5185 1664
rect 4865 1040 5185 1600
rect 8786 19616 9106 20640
rect 8786 19552 8794 19616
rect 8858 19552 8874 19616
rect 8938 19552 8954 19616
rect 9018 19552 9034 19616
rect 9098 19552 9106 19616
rect 8786 18528 9106 19552
rect 9630 19549 9690 21760
rect 9627 19548 9693 19549
rect 9627 19484 9628 19548
rect 9692 19484 9693 19548
rect 9627 19483 9693 19484
rect 10366 19005 10426 21760
rect 11102 20637 11162 21760
rect 11099 20636 11165 20637
rect 11099 20572 11100 20636
rect 11164 20572 11165 20636
rect 11099 20571 11165 20572
rect 11838 19549 11898 21760
rect 12574 20637 12634 21760
rect 12571 20636 12637 20637
rect 12571 20572 12572 20636
rect 12636 20572 12637 20636
rect 12571 20571 12637 20572
rect 12707 20160 13027 20720
rect 12707 20096 12715 20160
rect 12779 20096 12795 20160
rect 12859 20096 12875 20160
rect 12939 20096 12955 20160
rect 13019 20096 13027 20160
rect 11835 19548 11901 19549
rect 11835 19484 11836 19548
rect 11900 19484 11901 19548
rect 11835 19483 11901 19484
rect 12707 19072 13027 20096
rect 13310 19277 13370 21760
rect 14046 20093 14106 21760
rect 14782 20637 14842 21760
rect 14779 20636 14845 20637
rect 14779 20572 14780 20636
rect 14844 20572 14845 20636
rect 14779 20571 14845 20572
rect 14043 20092 14109 20093
rect 14043 20028 14044 20092
rect 14108 20028 14109 20092
rect 14043 20027 14109 20028
rect 13307 19276 13373 19277
rect 13307 19212 13308 19276
rect 13372 19212 13373 19276
rect 13307 19211 13373 19212
rect 12707 19008 12715 19072
rect 12779 19008 12795 19072
rect 12859 19008 12875 19072
rect 12939 19008 12955 19072
rect 13019 19008 13027 19072
rect 10363 19004 10429 19005
rect 10363 18940 10364 19004
rect 10428 18940 10429 19004
rect 10363 18939 10429 18940
rect 8786 18464 8794 18528
rect 8858 18464 8874 18528
rect 8938 18464 8954 18528
rect 9018 18464 9034 18528
rect 9098 18464 9106 18528
rect 8786 17440 9106 18464
rect 8786 17376 8794 17440
rect 8858 17376 8874 17440
rect 8938 17376 8954 17440
rect 9018 17376 9034 17440
rect 9098 17376 9106 17440
rect 8786 16352 9106 17376
rect 8786 16288 8794 16352
rect 8858 16288 8874 16352
rect 8938 16288 8954 16352
rect 9018 16288 9034 16352
rect 9098 16288 9106 16352
rect 8786 15264 9106 16288
rect 8786 15200 8794 15264
rect 8858 15200 8874 15264
rect 8938 15200 8954 15264
rect 9018 15200 9034 15264
rect 9098 15200 9106 15264
rect 8786 14176 9106 15200
rect 8786 14112 8794 14176
rect 8858 14112 8874 14176
rect 8938 14112 8954 14176
rect 9018 14112 9034 14176
rect 9098 14112 9106 14176
rect 8786 13088 9106 14112
rect 8786 13024 8794 13088
rect 8858 13024 8874 13088
rect 8938 13024 8954 13088
rect 9018 13024 9034 13088
rect 9098 13024 9106 13088
rect 8786 12000 9106 13024
rect 8786 11936 8794 12000
rect 8858 11936 8874 12000
rect 8938 11936 8954 12000
rect 9018 11936 9034 12000
rect 9098 11936 9106 12000
rect 8786 10912 9106 11936
rect 8786 10848 8794 10912
rect 8858 10848 8874 10912
rect 8938 10848 8954 10912
rect 9018 10848 9034 10912
rect 9098 10848 9106 10912
rect 8786 9824 9106 10848
rect 8786 9760 8794 9824
rect 8858 9760 8874 9824
rect 8938 9760 8954 9824
rect 9018 9760 9034 9824
rect 9098 9760 9106 9824
rect 8786 8736 9106 9760
rect 8786 8672 8794 8736
rect 8858 8672 8874 8736
rect 8938 8672 8954 8736
rect 9018 8672 9034 8736
rect 9098 8672 9106 8736
rect 8786 7648 9106 8672
rect 8786 7584 8794 7648
rect 8858 7584 8874 7648
rect 8938 7584 8954 7648
rect 9018 7584 9034 7648
rect 9098 7584 9106 7648
rect 8786 6560 9106 7584
rect 8786 6496 8794 6560
rect 8858 6496 8874 6560
rect 8938 6496 8954 6560
rect 9018 6496 9034 6560
rect 9098 6496 9106 6560
rect 8786 5472 9106 6496
rect 8786 5408 8794 5472
rect 8858 5408 8874 5472
rect 8938 5408 8954 5472
rect 9018 5408 9034 5472
rect 9098 5408 9106 5472
rect 8786 4384 9106 5408
rect 8786 4320 8794 4384
rect 8858 4320 8874 4384
rect 8938 4320 8954 4384
rect 9018 4320 9034 4384
rect 9098 4320 9106 4384
rect 8786 3296 9106 4320
rect 8786 3232 8794 3296
rect 8858 3232 8874 3296
rect 8938 3232 8954 3296
rect 9018 3232 9034 3296
rect 9098 3232 9106 3296
rect 8786 2208 9106 3232
rect 8786 2144 8794 2208
rect 8858 2144 8874 2208
rect 8938 2144 8954 2208
rect 9018 2144 9034 2208
rect 9098 2144 9106 2208
rect 8786 1120 9106 2144
rect 8786 1056 8794 1120
rect 8858 1056 8874 1120
rect 8938 1056 8954 1120
rect 9018 1056 9034 1120
rect 9098 1056 9106 1120
rect 8786 1040 9106 1056
rect 12707 17984 13027 19008
rect 15518 19005 15578 21760
rect 16254 19549 16314 21760
rect 16990 20909 17050 21760
rect 16987 20908 17053 20909
rect 16987 20844 16988 20908
rect 17052 20844 17053 20908
rect 16987 20843 17053 20844
rect 16628 20704 16948 20720
rect 16628 20640 16636 20704
rect 16700 20640 16716 20704
rect 16780 20640 16796 20704
rect 16860 20640 16876 20704
rect 16940 20640 16948 20704
rect 16628 19616 16948 20640
rect 16628 19552 16636 19616
rect 16700 19552 16716 19616
rect 16780 19552 16796 19616
rect 16860 19552 16876 19616
rect 16940 19552 16948 19616
rect 16251 19548 16317 19549
rect 16251 19484 16252 19548
rect 16316 19484 16317 19548
rect 16251 19483 16317 19484
rect 15515 19004 15581 19005
rect 15515 18940 15516 19004
rect 15580 18940 15581 19004
rect 15515 18939 15581 18940
rect 12707 17920 12715 17984
rect 12779 17920 12795 17984
rect 12859 17920 12875 17984
rect 12939 17920 12955 17984
rect 13019 17920 13027 17984
rect 12707 16896 13027 17920
rect 12707 16832 12715 16896
rect 12779 16832 12795 16896
rect 12859 16832 12875 16896
rect 12939 16832 12955 16896
rect 13019 16832 13027 16896
rect 12707 15808 13027 16832
rect 12707 15744 12715 15808
rect 12779 15744 12795 15808
rect 12859 15744 12875 15808
rect 12939 15744 12955 15808
rect 13019 15744 13027 15808
rect 12707 14720 13027 15744
rect 12707 14656 12715 14720
rect 12779 14656 12795 14720
rect 12859 14656 12875 14720
rect 12939 14656 12955 14720
rect 13019 14656 13027 14720
rect 12707 13632 13027 14656
rect 12707 13568 12715 13632
rect 12779 13568 12795 13632
rect 12859 13568 12875 13632
rect 12939 13568 12955 13632
rect 13019 13568 13027 13632
rect 12707 12544 13027 13568
rect 12707 12480 12715 12544
rect 12779 12480 12795 12544
rect 12859 12480 12875 12544
rect 12939 12480 12955 12544
rect 13019 12480 13027 12544
rect 12707 11456 13027 12480
rect 12707 11392 12715 11456
rect 12779 11392 12795 11456
rect 12859 11392 12875 11456
rect 12939 11392 12955 11456
rect 13019 11392 13027 11456
rect 12707 10368 13027 11392
rect 12707 10304 12715 10368
rect 12779 10304 12795 10368
rect 12859 10304 12875 10368
rect 12939 10304 12955 10368
rect 13019 10304 13027 10368
rect 12707 9280 13027 10304
rect 12707 9216 12715 9280
rect 12779 9216 12795 9280
rect 12859 9216 12875 9280
rect 12939 9216 12955 9280
rect 13019 9216 13027 9280
rect 12707 8192 13027 9216
rect 12707 8128 12715 8192
rect 12779 8128 12795 8192
rect 12859 8128 12875 8192
rect 12939 8128 12955 8192
rect 13019 8128 13027 8192
rect 12707 7104 13027 8128
rect 12707 7040 12715 7104
rect 12779 7040 12795 7104
rect 12859 7040 12875 7104
rect 12939 7040 12955 7104
rect 13019 7040 13027 7104
rect 12707 6016 13027 7040
rect 12707 5952 12715 6016
rect 12779 5952 12795 6016
rect 12859 5952 12875 6016
rect 12939 5952 12955 6016
rect 13019 5952 13027 6016
rect 12707 4928 13027 5952
rect 12707 4864 12715 4928
rect 12779 4864 12795 4928
rect 12859 4864 12875 4928
rect 12939 4864 12955 4928
rect 13019 4864 13027 4928
rect 12707 3840 13027 4864
rect 12707 3776 12715 3840
rect 12779 3776 12795 3840
rect 12859 3776 12875 3840
rect 12939 3776 12955 3840
rect 13019 3776 13027 3840
rect 12707 2752 13027 3776
rect 12707 2688 12715 2752
rect 12779 2688 12795 2752
rect 12859 2688 12875 2752
rect 12939 2688 12955 2752
rect 13019 2688 13027 2752
rect 12707 1664 13027 2688
rect 12707 1600 12715 1664
rect 12779 1600 12795 1664
rect 12859 1600 12875 1664
rect 12939 1600 12955 1664
rect 13019 1600 13027 1664
rect 12707 1040 13027 1600
rect 16628 18528 16948 19552
rect 17726 19413 17786 21760
rect 18462 20637 18522 21760
rect 19198 20773 19258 21760
rect 19934 21181 19994 21760
rect 19931 21180 19997 21181
rect 19931 21116 19932 21180
rect 19996 21116 19997 21180
rect 19931 21115 19997 21116
rect 20670 20909 20730 21760
rect 20667 20908 20733 20909
rect 20667 20844 20668 20908
rect 20732 20844 20733 20908
rect 20667 20843 20733 20844
rect 19195 20772 19261 20773
rect 19195 20708 19196 20772
rect 19260 20708 19261 20772
rect 19195 20707 19261 20708
rect 18459 20636 18525 20637
rect 18459 20572 18460 20636
rect 18524 20572 18525 20636
rect 18459 20571 18525 20572
rect 20549 20160 20869 20720
rect 21406 20501 21466 21760
rect 22142 21045 22202 21760
rect 22878 21045 22938 21760
rect 23614 21181 23674 21760
rect 23611 21180 23677 21181
rect 23611 21116 23612 21180
rect 23676 21116 23677 21180
rect 23611 21115 23677 21116
rect 22139 21044 22205 21045
rect 22139 20980 22140 21044
rect 22204 20980 22205 21044
rect 22139 20979 22205 20980
rect 22875 21044 22941 21045
rect 22875 20980 22876 21044
rect 22940 20980 22941 21044
rect 22875 20979 22941 20980
rect 21403 20500 21469 20501
rect 21403 20436 21404 20500
rect 21468 20436 21469 20500
rect 21403 20435 21469 20436
rect 20549 20096 20557 20160
rect 20621 20096 20637 20160
rect 20701 20096 20717 20160
rect 20781 20096 20797 20160
rect 20861 20096 20869 20160
rect 17723 19412 17789 19413
rect 17723 19348 17724 19412
rect 17788 19348 17789 19412
rect 17723 19347 17789 19348
rect 16628 18464 16636 18528
rect 16700 18464 16716 18528
rect 16780 18464 16796 18528
rect 16860 18464 16876 18528
rect 16940 18464 16948 18528
rect 16628 17440 16948 18464
rect 16628 17376 16636 17440
rect 16700 17376 16716 17440
rect 16780 17376 16796 17440
rect 16860 17376 16876 17440
rect 16940 17376 16948 17440
rect 16628 16352 16948 17376
rect 16628 16288 16636 16352
rect 16700 16288 16716 16352
rect 16780 16288 16796 16352
rect 16860 16288 16876 16352
rect 16940 16288 16948 16352
rect 16628 15264 16948 16288
rect 16628 15200 16636 15264
rect 16700 15200 16716 15264
rect 16780 15200 16796 15264
rect 16860 15200 16876 15264
rect 16940 15200 16948 15264
rect 16628 14176 16948 15200
rect 16628 14112 16636 14176
rect 16700 14112 16716 14176
rect 16780 14112 16796 14176
rect 16860 14112 16876 14176
rect 16940 14112 16948 14176
rect 16628 13088 16948 14112
rect 16628 13024 16636 13088
rect 16700 13024 16716 13088
rect 16780 13024 16796 13088
rect 16860 13024 16876 13088
rect 16940 13024 16948 13088
rect 16628 12000 16948 13024
rect 16628 11936 16636 12000
rect 16700 11936 16716 12000
rect 16780 11936 16796 12000
rect 16860 11936 16876 12000
rect 16940 11936 16948 12000
rect 16628 10912 16948 11936
rect 16628 10848 16636 10912
rect 16700 10848 16716 10912
rect 16780 10848 16796 10912
rect 16860 10848 16876 10912
rect 16940 10848 16948 10912
rect 16628 9824 16948 10848
rect 16628 9760 16636 9824
rect 16700 9760 16716 9824
rect 16780 9760 16796 9824
rect 16860 9760 16876 9824
rect 16940 9760 16948 9824
rect 16628 8736 16948 9760
rect 16628 8672 16636 8736
rect 16700 8672 16716 8736
rect 16780 8672 16796 8736
rect 16860 8672 16876 8736
rect 16940 8672 16948 8736
rect 16628 7648 16948 8672
rect 16628 7584 16636 7648
rect 16700 7584 16716 7648
rect 16780 7584 16796 7648
rect 16860 7584 16876 7648
rect 16940 7584 16948 7648
rect 16628 6560 16948 7584
rect 16628 6496 16636 6560
rect 16700 6496 16716 6560
rect 16780 6496 16796 6560
rect 16860 6496 16876 6560
rect 16940 6496 16948 6560
rect 16628 5472 16948 6496
rect 16628 5408 16636 5472
rect 16700 5408 16716 5472
rect 16780 5408 16796 5472
rect 16860 5408 16876 5472
rect 16940 5408 16948 5472
rect 16628 4384 16948 5408
rect 16628 4320 16636 4384
rect 16700 4320 16716 4384
rect 16780 4320 16796 4384
rect 16860 4320 16876 4384
rect 16940 4320 16948 4384
rect 16628 3296 16948 4320
rect 16628 3232 16636 3296
rect 16700 3232 16716 3296
rect 16780 3232 16796 3296
rect 16860 3232 16876 3296
rect 16940 3232 16948 3296
rect 16628 2208 16948 3232
rect 16628 2144 16636 2208
rect 16700 2144 16716 2208
rect 16780 2144 16796 2208
rect 16860 2144 16876 2208
rect 16940 2144 16948 2208
rect 16628 1120 16948 2144
rect 16628 1056 16636 1120
rect 16700 1056 16716 1120
rect 16780 1056 16796 1120
rect 16860 1056 16876 1120
rect 16940 1056 16948 1120
rect 16628 1040 16948 1056
rect 20549 19072 20869 20096
rect 24350 20090 24410 21760
rect 25086 21560 25146 21760
rect 25822 21560 25882 21760
rect 26558 21560 26618 21760
rect 27294 21560 27354 21760
rect 28030 21560 28090 21760
rect 28766 21560 28826 21760
rect 29502 21560 29562 21760
rect 24166 20030 24410 20090
rect 24470 20704 24790 20720
rect 24470 20640 24478 20704
rect 24542 20640 24558 20704
rect 24622 20640 24638 20704
rect 24702 20640 24718 20704
rect 24782 20640 24790 20704
rect 24166 19277 24226 20030
rect 24470 19616 24790 20640
rect 24470 19552 24478 19616
rect 24542 19552 24558 19616
rect 24622 19552 24638 19616
rect 24702 19552 24718 19616
rect 24782 19552 24790 19616
rect 24163 19276 24229 19277
rect 24163 19212 24164 19276
rect 24228 19212 24229 19276
rect 24163 19211 24229 19212
rect 20549 19008 20557 19072
rect 20621 19008 20637 19072
rect 20701 19008 20717 19072
rect 20781 19008 20797 19072
rect 20861 19008 20869 19072
rect 20549 17984 20869 19008
rect 20549 17920 20557 17984
rect 20621 17920 20637 17984
rect 20701 17920 20717 17984
rect 20781 17920 20797 17984
rect 20861 17920 20869 17984
rect 20549 16896 20869 17920
rect 20549 16832 20557 16896
rect 20621 16832 20637 16896
rect 20701 16832 20717 16896
rect 20781 16832 20797 16896
rect 20861 16832 20869 16896
rect 20549 15808 20869 16832
rect 20549 15744 20557 15808
rect 20621 15744 20637 15808
rect 20701 15744 20717 15808
rect 20781 15744 20797 15808
rect 20861 15744 20869 15808
rect 20549 14720 20869 15744
rect 20549 14656 20557 14720
rect 20621 14656 20637 14720
rect 20701 14656 20717 14720
rect 20781 14656 20797 14720
rect 20861 14656 20869 14720
rect 20549 13632 20869 14656
rect 20549 13568 20557 13632
rect 20621 13568 20637 13632
rect 20701 13568 20717 13632
rect 20781 13568 20797 13632
rect 20861 13568 20869 13632
rect 20549 12544 20869 13568
rect 20549 12480 20557 12544
rect 20621 12480 20637 12544
rect 20701 12480 20717 12544
rect 20781 12480 20797 12544
rect 20861 12480 20869 12544
rect 20549 11456 20869 12480
rect 20549 11392 20557 11456
rect 20621 11392 20637 11456
rect 20701 11392 20717 11456
rect 20781 11392 20797 11456
rect 20861 11392 20869 11456
rect 20549 10368 20869 11392
rect 20549 10304 20557 10368
rect 20621 10304 20637 10368
rect 20701 10304 20717 10368
rect 20781 10304 20797 10368
rect 20861 10304 20869 10368
rect 20549 9280 20869 10304
rect 20549 9216 20557 9280
rect 20621 9216 20637 9280
rect 20701 9216 20717 9280
rect 20781 9216 20797 9280
rect 20861 9216 20869 9280
rect 20549 8192 20869 9216
rect 20549 8128 20557 8192
rect 20621 8128 20637 8192
rect 20701 8128 20717 8192
rect 20781 8128 20797 8192
rect 20861 8128 20869 8192
rect 20549 7104 20869 8128
rect 20549 7040 20557 7104
rect 20621 7040 20637 7104
rect 20701 7040 20717 7104
rect 20781 7040 20797 7104
rect 20861 7040 20869 7104
rect 20549 6016 20869 7040
rect 20549 5952 20557 6016
rect 20621 5952 20637 6016
rect 20701 5952 20717 6016
rect 20781 5952 20797 6016
rect 20861 5952 20869 6016
rect 20549 4928 20869 5952
rect 20549 4864 20557 4928
rect 20621 4864 20637 4928
rect 20701 4864 20717 4928
rect 20781 4864 20797 4928
rect 20861 4864 20869 4928
rect 20549 3840 20869 4864
rect 20549 3776 20557 3840
rect 20621 3776 20637 3840
rect 20701 3776 20717 3840
rect 20781 3776 20797 3840
rect 20861 3776 20869 3840
rect 20549 2752 20869 3776
rect 20549 2688 20557 2752
rect 20621 2688 20637 2752
rect 20701 2688 20717 2752
rect 20781 2688 20797 2752
rect 20861 2688 20869 2752
rect 20549 1664 20869 2688
rect 20549 1600 20557 1664
rect 20621 1600 20637 1664
rect 20701 1600 20717 1664
rect 20781 1600 20797 1664
rect 20861 1600 20869 1664
rect 20549 1040 20869 1600
rect 24470 18528 24790 19552
rect 24470 18464 24478 18528
rect 24542 18464 24558 18528
rect 24622 18464 24638 18528
rect 24702 18464 24718 18528
rect 24782 18464 24790 18528
rect 24470 17440 24790 18464
rect 24470 17376 24478 17440
rect 24542 17376 24558 17440
rect 24622 17376 24638 17440
rect 24702 17376 24718 17440
rect 24782 17376 24790 17440
rect 24470 16352 24790 17376
rect 24470 16288 24478 16352
rect 24542 16288 24558 16352
rect 24622 16288 24638 16352
rect 24702 16288 24718 16352
rect 24782 16288 24790 16352
rect 24470 15264 24790 16288
rect 24470 15200 24478 15264
rect 24542 15200 24558 15264
rect 24622 15200 24638 15264
rect 24702 15200 24718 15264
rect 24782 15200 24790 15264
rect 24470 14176 24790 15200
rect 24470 14112 24478 14176
rect 24542 14112 24558 14176
rect 24622 14112 24638 14176
rect 24702 14112 24718 14176
rect 24782 14112 24790 14176
rect 24470 13088 24790 14112
rect 24470 13024 24478 13088
rect 24542 13024 24558 13088
rect 24622 13024 24638 13088
rect 24702 13024 24718 13088
rect 24782 13024 24790 13088
rect 24470 12000 24790 13024
rect 24470 11936 24478 12000
rect 24542 11936 24558 12000
rect 24622 11936 24638 12000
rect 24702 11936 24718 12000
rect 24782 11936 24790 12000
rect 24470 10912 24790 11936
rect 24470 10848 24478 10912
rect 24542 10848 24558 10912
rect 24622 10848 24638 10912
rect 24702 10848 24718 10912
rect 24782 10848 24790 10912
rect 24470 9824 24790 10848
rect 24470 9760 24478 9824
rect 24542 9760 24558 9824
rect 24622 9760 24638 9824
rect 24702 9760 24718 9824
rect 24782 9760 24790 9824
rect 24470 8736 24790 9760
rect 24470 8672 24478 8736
rect 24542 8672 24558 8736
rect 24622 8672 24638 8736
rect 24702 8672 24718 8736
rect 24782 8672 24790 8736
rect 24470 7648 24790 8672
rect 24470 7584 24478 7648
rect 24542 7584 24558 7648
rect 24622 7584 24638 7648
rect 24702 7584 24718 7648
rect 24782 7584 24790 7648
rect 24470 6560 24790 7584
rect 24470 6496 24478 6560
rect 24542 6496 24558 6560
rect 24622 6496 24638 6560
rect 24702 6496 24718 6560
rect 24782 6496 24790 6560
rect 24470 5472 24790 6496
rect 24470 5408 24478 5472
rect 24542 5408 24558 5472
rect 24622 5408 24638 5472
rect 24702 5408 24718 5472
rect 24782 5408 24790 5472
rect 24470 4384 24790 5408
rect 24470 4320 24478 4384
rect 24542 4320 24558 4384
rect 24622 4320 24638 4384
rect 24702 4320 24718 4384
rect 24782 4320 24790 4384
rect 24470 3296 24790 4320
rect 24470 3232 24478 3296
rect 24542 3232 24558 3296
rect 24622 3232 24638 3296
rect 24702 3232 24718 3296
rect 24782 3232 24790 3296
rect 24470 2208 24790 3232
rect 24470 2144 24478 2208
rect 24542 2144 24558 2208
rect 24622 2144 24638 2208
rect 24702 2144 24718 2208
rect 24782 2144 24790 2208
rect 24470 1120 24790 2144
rect 24470 1056 24478 1120
rect 24542 1056 24558 1120
rect 24622 1056 24638 1120
rect 24702 1056 24718 1120
rect 24782 1056 24790 1120
rect 24470 1040 24790 1056
rect 28391 20160 28711 20720
rect 28391 20096 28399 20160
rect 28463 20096 28479 20160
rect 28543 20096 28559 20160
rect 28623 20096 28639 20160
rect 28703 20096 28711 20160
rect 28391 19072 28711 20096
rect 28391 19008 28399 19072
rect 28463 19008 28479 19072
rect 28543 19008 28559 19072
rect 28623 19008 28639 19072
rect 28703 19008 28711 19072
rect 28391 17984 28711 19008
rect 28391 17920 28399 17984
rect 28463 17920 28479 17984
rect 28543 17920 28559 17984
rect 28623 17920 28639 17984
rect 28703 17920 28711 17984
rect 28391 16896 28711 17920
rect 30238 17917 30298 21760
rect 30974 19685 31034 21760
rect 31710 20773 31770 21760
rect 32446 21560 32506 21760
rect 31707 20772 31773 20773
rect 31707 20708 31708 20772
rect 31772 20708 31773 20772
rect 31707 20707 31773 20708
rect 32312 20704 32632 20720
rect 32312 20640 32320 20704
rect 32384 20640 32400 20704
rect 32464 20640 32480 20704
rect 32544 20640 32560 20704
rect 32624 20640 32632 20704
rect 30971 19684 31037 19685
rect 30971 19620 30972 19684
rect 31036 19620 31037 19684
rect 30971 19619 31037 19620
rect 32312 19616 32632 20640
rect 32312 19552 32320 19616
rect 32384 19552 32400 19616
rect 32464 19552 32480 19616
rect 32544 19552 32560 19616
rect 32624 19552 32632 19616
rect 32312 18528 32632 19552
rect 32312 18464 32320 18528
rect 32384 18464 32400 18528
rect 32464 18464 32480 18528
rect 32544 18464 32560 18528
rect 32624 18464 32632 18528
rect 30235 17916 30301 17917
rect 30235 17852 30236 17916
rect 30300 17852 30301 17916
rect 30235 17851 30301 17852
rect 28391 16832 28399 16896
rect 28463 16832 28479 16896
rect 28543 16832 28559 16896
rect 28623 16832 28639 16896
rect 28703 16832 28711 16896
rect 28391 15808 28711 16832
rect 28391 15744 28399 15808
rect 28463 15744 28479 15808
rect 28543 15744 28559 15808
rect 28623 15744 28639 15808
rect 28703 15744 28711 15808
rect 28391 14720 28711 15744
rect 28391 14656 28399 14720
rect 28463 14656 28479 14720
rect 28543 14656 28559 14720
rect 28623 14656 28639 14720
rect 28703 14656 28711 14720
rect 28391 13632 28711 14656
rect 28391 13568 28399 13632
rect 28463 13568 28479 13632
rect 28543 13568 28559 13632
rect 28623 13568 28639 13632
rect 28703 13568 28711 13632
rect 28391 12544 28711 13568
rect 28391 12480 28399 12544
rect 28463 12480 28479 12544
rect 28543 12480 28559 12544
rect 28623 12480 28639 12544
rect 28703 12480 28711 12544
rect 28391 11456 28711 12480
rect 28391 11392 28399 11456
rect 28463 11392 28479 11456
rect 28543 11392 28559 11456
rect 28623 11392 28639 11456
rect 28703 11392 28711 11456
rect 28391 10368 28711 11392
rect 28391 10304 28399 10368
rect 28463 10304 28479 10368
rect 28543 10304 28559 10368
rect 28623 10304 28639 10368
rect 28703 10304 28711 10368
rect 28391 9280 28711 10304
rect 28391 9216 28399 9280
rect 28463 9216 28479 9280
rect 28543 9216 28559 9280
rect 28623 9216 28639 9280
rect 28703 9216 28711 9280
rect 28391 8192 28711 9216
rect 28391 8128 28399 8192
rect 28463 8128 28479 8192
rect 28543 8128 28559 8192
rect 28623 8128 28639 8192
rect 28703 8128 28711 8192
rect 28391 7104 28711 8128
rect 28391 7040 28399 7104
rect 28463 7040 28479 7104
rect 28543 7040 28559 7104
rect 28623 7040 28639 7104
rect 28703 7040 28711 7104
rect 28391 6016 28711 7040
rect 28391 5952 28399 6016
rect 28463 5952 28479 6016
rect 28543 5952 28559 6016
rect 28623 5952 28639 6016
rect 28703 5952 28711 6016
rect 28391 4928 28711 5952
rect 28391 4864 28399 4928
rect 28463 4864 28479 4928
rect 28543 4864 28559 4928
rect 28623 4864 28639 4928
rect 28703 4864 28711 4928
rect 28391 3840 28711 4864
rect 28391 3776 28399 3840
rect 28463 3776 28479 3840
rect 28543 3776 28559 3840
rect 28623 3776 28639 3840
rect 28703 3776 28711 3840
rect 28391 2752 28711 3776
rect 28391 2688 28399 2752
rect 28463 2688 28479 2752
rect 28543 2688 28559 2752
rect 28623 2688 28639 2752
rect 28703 2688 28711 2752
rect 28391 1664 28711 2688
rect 28391 1600 28399 1664
rect 28463 1600 28479 1664
rect 28543 1600 28559 1664
rect 28623 1600 28639 1664
rect 28703 1600 28711 1664
rect 28391 1040 28711 1600
rect 32312 17440 32632 18464
rect 32312 17376 32320 17440
rect 32384 17376 32400 17440
rect 32464 17376 32480 17440
rect 32544 17376 32560 17440
rect 32624 17376 32632 17440
rect 32312 16352 32632 17376
rect 32312 16288 32320 16352
rect 32384 16288 32400 16352
rect 32464 16288 32480 16352
rect 32544 16288 32560 16352
rect 32624 16288 32632 16352
rect 32312 15264 32632 16288
rect 32312 15200 32320 15264
rect 32384 15200 32400 15264
rect 32464 15200 32480 15264
rect 32544 15200 32560 15264
rect 32624 15200 32632 15264
rect 32312 14176 32632 15200
rect 32312 14112 32320 14176
rect 32384 14112 32400 14176
rect 32464 14112 32480 14176
rect 32544 14112 32560 14176
rect 32624 14112 32632 14176
rect 32312 13088 32632 14112
rect 32312 13024 32320 13088
rect 32384 13024 32400 13088
rect 32464 13024 32480 13088
rect 32544 13024 32560 13088
rect 32624 13024 32632 13088
rect 32312 12000 32632 13024
rect 32312 11936 32320 12000
rect 32384 11936 32400 12000
rect 32464 11936 32480 12000
rect 32544 11936 32560 12000
rect 32624 11936 32632 12000
rect 32312 10912 32632 11936
rect 32312 10848 32320 10912
rect 32384 10848 32400 10912
rect 32464 10848 32480 10912
rect 32544 10848 32560 10912
rect 32624 10848 32632 10912
rect 32312 9824 32632 10848
rect 32312 9760 32320 9824
rect 32384 9760 32400 9824
rect 32464 9760 32480 9824
rect 32544 9760 32560 9824
rect 32624 9760 32632 9824
rect 32312 8736 32632 9760
rect 32312 8672 32320 8736
rect 32384 8672 32400 8736
rect 32464 8672 32480 8736
rect 32544 8672 32560 8736
rect 32624 8672 32632 8736
rect 32312 7648 32632 8672
rect 32312 7584 32320 7648
rect 32384 7584 32400 7648
rect 32464 7584 32480 7648
rect 32544 7584 32560 7648
rect 32624 7584 32632 7648
rect 32312 6560 32632 7584
rect 32312 6496 32320 6560
rect 32384 6496 32400 6560
rect 32464 6496 32480 6560
rect 32544 6496 32560 6560
rect 32624 6496 32632 6560
rect 32312 5472 32632 6496
rect 32312 5408 32320 5472
rect 32384 5408 32400 5472
rect 32464 5408 32480 5472
rect 32544 5408 32560 5472
rect 32624 5408 32632 5472
rect 32312 4384 32632 5408
rect 32312 4320 32320 4384
rect 32384 4320 32400 4384
rect 32464 4320 32480 4384
rect 32544 4320 32560 4384
rect 32624 4320 32632 4384
rect 32312 3296 32632 4320
rect 32312 3232 32320 3296
rect 32384 3232 32400 3296
rect 32464 3232 32480 3296
rect 32544 3232 32560 3296
rect 32624 3232 32632 3296
rect 32312 2208 32632 3232
rect 32312 2144 32320 2208
rect 32384 2144 32400 2208
rect 32464 2144 32480 2208
rect 32544 2144 32560 2208
rect 32624 2144 32632 2208
rect 32312 1120 32632 2144
rect 32312 1056 32320 1120
rect 32384 1056 32400 1120
rect 32464 1056 32480 1120
rect 32544 1056 32560 1120
rect 32624 1056 32632 1120
rect 32312 1040 32632 1056
use sky130_fd_sc_hd__clkbuf_2  _035_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14812 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _036_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15272 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _037_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _038_
timestamp 1676037725
transform 1 0 14812 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _039_
timestamp 1676037725
transform -1 0 13800 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _040_
timestamp 1676037725
transform -1 0 17296 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _041_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17480 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _042_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 14812 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _043_
timestamp 1676037725
transform -1 0 12972 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _044_
timestamp 1676037725
transform -1 0 14444 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _045_
timestamp 1676037725
transform -1 0 12696 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _046_
timestamp 1676037725
transform -1 0 16284 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _047_
timestamp 1676037725
transform -1 0 12236 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _048_
timestamp 1676037725
transform -1 0 16100 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _049_
timestamp 1676037725
transform -1 0 11776 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _050_
timestamp 1676037725
transform -1 0 15456 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _051_
timestamp 1676037725
transform -1 0 11224 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _052_
timestamp 1676037725
transform -1 0 13616 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _053_
timestamp 1676037725
transform -1 0 10764 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _054_
timestamp 1676037725
transform -1 0 13800 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _055_
timestamp 1676037725
transform -1 0 11684 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _056_
timestamp 1676037725
transform -1 0 17296 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _057_
timestamp 1676037725
transform -1 0 12604 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _058_
timestamp 1676037725
transform 1 0 19688 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1676037725
transform -1 0 18952 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _060_
timestamp 1676037725
transform 1 0 19412 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1676037725
transform -1 0 18308 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _062_
timestamp 1676037725
transform 1 0 19228 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1676037725
transform -1 0 18032 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _064_
timestamp 1676037725
transform 1 0 20608 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1676037725
transform -1 0 16376 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _066_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25024 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _067_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 24380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _068_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 25024 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _069_
timestamp 1676037725
transform 1 0 23184 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _070_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 24656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _071_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23092 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _072_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19596 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _073_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23092 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _074_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22172 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1676037725
transform -1 0 25668 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _076_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23460 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _077_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 23276 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _078_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 24012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _079_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 24840 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _080_
timestamp 1676037725
transform 1 0 22448 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _081_
timestamp 1676037725
transform -1 0 20332 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _082_
timestamp 1676037725
transform 1 0 18308 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _083_
timestamp 1676037725
transform 1 0 20424 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1676037725
transform -1 0 17388 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_2  _085_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26312 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _086_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _087_
timestamp 1676037725
transform 1 0 27140 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _088_
timestamp 1676037725
transform -1 0 26680 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _089_
timestamp 1676037725
transform 1 0 26128 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _090_
timestamp 1676037725
transform -1 0 29440 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _091_
timestamp 1676037725
transform 1 0 29992 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _092_
timestamp 1676037725
transform 1 0 29900 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _093_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__conb_1  _093__13 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 29256 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1676037725
transform 1 0 6348 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1676037725
transform 1 0 5612 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1676037725
transform 1 0 4140 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1676037725
transform -1 0 4140 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1676037725
transform 1 0 2852 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1676037725
transform -1 0 2484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1676037725
transform -1 0 2668 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 31556 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1676037725
transform -1 0 27876 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1676037725
transform 1 0 29992 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  fanout11
timestamp 1676037725
transform -1 0 16376 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout12
timestamp 1676037725
transform -1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1676037725
transform 1 0 2484 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1676037725
transform 1 0 3772 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1676037725
transform 1 0 4876 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1676037725
transform 1 0 6348 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1676037725
transform 1 0 7452 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1676037725
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1676037725
transform 1 0 8924 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1676037725
transform 1 0 10028 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1676037725
transform 1 0 11132 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1676037725
transform 1 0 11500 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1676037725
transform 1 0 12604 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1676037725
transform 1 0 13708 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1676037725
transform 1 0 14076 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1676037725
transform 1 0 15180 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1676037725
transform 1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1676037725
transform 1 0 16652 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1676037725
transform 1 0 17756 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1676037725
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1676037725
transform 1 0 19228 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1676037725
transform 1 0 20332 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1676037725
transform 1 0 21436 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1676037725
transform 1 0 21804 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1676037725
transform 1 0 22908 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1676037725
transform 1 0 24012 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1676037725
transform 1 0 24380 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1676037725
transform 1 0 25484 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1676037725
transform 1 0 26588 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1676037725
transform 1 0 26956 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1676037725
transform 1 0 28060 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1676037725
transform 1 0 29164 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1676037725
transform 1 0 29532 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1676037725
transform 1 0 30636 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1676037725
transform 1 0 31740 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_337
timestamp 1676037725
transform 1 0 32108 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5796 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10764 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1676037725
transform 1 0 18860 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1676037725
transform 1 0 19964 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1676037725
transform 1 0 21068 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1676037725
transform 1 0 25116 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1676037725
transform 1 0 26220 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1676037725
transform 1 0 26772 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1676037725
transform 1 0 29164 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1676037725
transform 1 0 30268 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1676037725
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1676037725
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1676037725
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1676037725
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1676037725
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1676037725
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1676037725
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1676037725
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1676037725
transform 1 0 17388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1676037725
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1676037725
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1676037725
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1676037725
transform 1 0 21436 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1676037725
transform 1 0 22540 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1676037725
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1676037725
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1676037725
transform 1 0 26588 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1676037725
transform 1 0 27692 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1676037725
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1676037725
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_333
timestamp 1676037725
transform 1 0 31740 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1676037725
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1676037725
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_337
timestamp 1676037725
transform 1 0 32108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1676037725
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_337
timestamp 1676037725
transform 1 0 32108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1676037725
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_337
timestamp 1676037725
transform 1 0 32108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1676037725
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1676037725
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1676037725
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1676037725
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_337
timestamp 1676037725
transform 1 0 32108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1676037725
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1676037725
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1676037725
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1676037725
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1676037725
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1676037725
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1676037725
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1676037725
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1676037725
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_333
timestamp 1676037725
transform 1 0 31740 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_337
timestamp 1676037725
transform 1 0 32108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1676037725
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1676037725
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1676037725
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1676037725
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1676037725
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1676037725
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1676037725
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_329
timestamp 1676037725
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1676037725
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1676037725
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 1676037725
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 1676037725
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1676037725
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1676037725
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 1676037725
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 1676037725
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1676037725
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_321
timestamp 1676037725
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_333
timestamp 1676037725
transform 1 0 31740 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_337
timestamp 1676037725
transform 1 0 32108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 1676037725
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 1676037725
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 1676037725
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1676037725
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 1676037725
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 1676037725
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_261
timestamp 1676037725
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_273
timestamp 1676037725
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1676037725
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1676037725
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1676037725
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 1676037725
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_329
timestamp 1676037725
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 1676037725
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 1676037725
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1676037725
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 1676037725
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 1676037725
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 1676037725
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1676037725
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1676037725
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 1676037725
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1676037725
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1676037725
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_321
timestamp 1676037725
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_333
timestamp 1676037725
transform 1 0 31740 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_337
timestamp 1676037725
transform 1 0 32108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1676037725
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 1676037725
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 1676037725
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 1676037725
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1676037725
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 1676037725
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 1676037725
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 1676037725
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 1676037725
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1676037725
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1676037725
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1676037725
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 1676037725
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 1676037725
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 1676037725
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 1676037725
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 1676037725
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1676037725
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 1676037725
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 1676037725
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_233
timestamp 1676037725
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_245
timestamp 1676037725
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1676037725
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1676037725
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1676037725
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 1676037725
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 1676037725
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1676037725
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 1676037725
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_333
timestamp 1676037725
transform 1 0 31740 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_337
timestamp 1676037725
transform 1 0 32108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 1676037725
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1676037725
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_193
timestamp 1676037725
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_205
timestamp 1676037725
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 1676037725
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1676037725
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 1676037725
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 1676037725
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 1676037725
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_273
timestamp 1676037725
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1676037725
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1676037725
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1676037725
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 1676037725
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_329
timestamp 1676037725
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 1676037725
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1676037725
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1676037725
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 1676037725
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 1676037725
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1676037725
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 1676037725
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 1676037725
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_233
timestamp 1676037725
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_245
timestamp 1676037725
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1676037725
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1676037725
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 1676037725
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_289
timestamp 1676037725
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_301
timestamp 1676037725
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1676037725
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_321
timestamp 1676037725
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_333
timestamp 1676037725
transform 1 0 31740 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_337
timestamp 1676037725
transform 1 0 32108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1676037725
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 1676037725
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 1676037725
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_193
timestamp 1676037725
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_205
timestamp 1676037725
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_217
timestamp 1676037725
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1676037725
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1676037725
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1676037725
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 1676037725
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 1676037725
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1676037725
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1676037725
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 1676037725
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 1676037725
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_329
timestamp 1676037725
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_335
timestamp 1676037725
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1676037725
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1676037725
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1676037725
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 1676037725
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 1676037725
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1676037725
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 1676037725
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 1676037725
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 1676037725
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 1676037725
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1676037725
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1676037725
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1676037725
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1676037725
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 1676037725
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1676037725
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_321
timestamp 1676037725
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_333
timestamp 1676037725
transform 1 0 31740 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_337
timestamp 1676037725
transform 1 0 32108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1676037725
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1676037725
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1676037725
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1676037725
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1676037725
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1676037725
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 1676037725
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 1676037725
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 1676037725
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1676037725
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1676037725
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 1676037725
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 1676037725
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 1676037725
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1676037725
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1676037725
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 1676037725
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 1676037725
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_329
timestamp 1676037725
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 1676037725
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1676037725
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1676037725
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1676037725
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1676037725
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 1676037725
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 1676037725
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 1676037725
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 1676037725
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1676037725
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 1676037725
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 1676037725
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_233
timestamp 1676037725
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 1676037725
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1676037725
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 1676037725
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 1676037725
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 1676037725
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 1676037725
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1676037725
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_321
timestamp 1676037725
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_333
timestamp 1676037725
transform 1 0 31740 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_337
timestamp 1676037725
transform 1 0 32108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1676037725
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1676037725
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1676037725
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1676037725
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1676037725
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 1676037725
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1676037725
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 1676037725
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1676037725
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 1676037725
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 1676037725
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_261
timestamp 1676037725
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 1676037725
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1676037725
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1676037725
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 1676037725
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 1676037725
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_329
timestamp 1676037725
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_335
timestamp 1676037725
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1676037725
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1676037725
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1676037725
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1676037725
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 1676037725
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1676037725
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1676037725
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 1676037725
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 1676037725
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 1676037725
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1676037725
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 1676037725
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 1676037725
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 1676037725
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 1676037725
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1676037725
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_321
timestamp 1676037725
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_333
timestamp 1676037725
transform 1 0 31740 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_337
timestamp 1676037725
transform 1 0 32108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1676037725
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1676037725
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1676037725
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1676037725
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 1676037725
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 1676037725
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 1676037725
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 1676037725
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1676037725
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 1676037725
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 1676037725
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 1676037725
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 1676037725
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1676037725
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1676037725
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1676037725
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 1676037725
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_329
timestamp 1676037725
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 1676037725
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1676037725
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1676037725
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1676037725
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1676037725
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1676037725
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 1676037725
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1676037725
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1676037725
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1676037725
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 1676037725
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 1676037725
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 1676037725
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1676037725
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1676037725
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 1676037725
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_289
timestamp 1676037725
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 1676037725
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1676037725
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_321
timestamp 1676037725
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_333
timestamp 1676037725
transform 1 0 31740 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_337
timestamp 1676037725
transform 1 0 32108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 1676037725
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1676037725
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1676037725
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 1676037725
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 1676037725
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 1676037725
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1676037725
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1676037725
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1676037725
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1676037725
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 1676037725
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1676037725
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1676037725
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 1676037725
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 1676037725
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_329
timestamp 1676037725
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 1676037725
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1676037725
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1676037725
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 1676037725
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 1676037725
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 1676037725
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1676037725
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 1676037725
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 1676037725
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 1676037725
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1676037725
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1676037725
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_265
timestamp 1676037725
transform 1 0 25484 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_291
timestamp 1676037725
transform 1 0 27876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_303
timestamp 1676037725
transform 1 0 28980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1676037725
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_321 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30636 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_326
timestamp 1676037725
transform 1 0 31096 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_333
timestamp 1676037725
transform 1 0 31740 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_337
timestamp 1676037725
transform 1 0 32108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_149 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_157
timestamp 1676037725
transform 1 0 15548 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_163
timestamp 1676037725
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1676037725
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1676037725
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_193
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_208
timestamp 1676037725
transform 1 0 20240 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_220
timestamp 1676037725
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_233
timestamp 1676037725
transform 1 0 22540 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_241
timestamp 1676037725
transform 1 0 23276 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_249
timestamp 1676037725
transform 1 0 24012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_256
timestamp 1676037725
transform 1 0 24656 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_263
timestamp 1676037725
transform 1 0 25300 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_275
timestamp 1676037725
transform 1 0 26404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1676037725
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_287
timestamp 1676037725
transform 1 0 27508 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_308
timestamp 1676037725
transform 1 0 29440 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_334
timestamp 1676037725
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1676037725
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_109
timestamp 1676037725
transform 1 0 11132 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_116
timestamp 1676037725
transform 1 0 11776 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_128
timestamp 1676037725
transform 1 0 12880 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_132
timestamp 1676037725
transform 1 0 13248 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_138
timestamp 1676037725
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_149
timestamp 1676037725
transform 1 0 14812 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_156
timestamp 1676037725
transform 1 0 15456 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_165
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 1676037725
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 1676037725
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1676037725
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_201
timestamp 1676037725
transform 1 0 19596 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_209
timestamp 1676037725
transform 1 0 20332 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_216
timestamp 1676037725
transform 1 0 20976 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_228
timestamp 1676037725
transform 1 0 22080 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_239
timestamp 1676037725
transform 1 0 23092 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_250
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_258
timestamp 1676037725
transform 1 0 24840 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_265
timestamp 1676037725
transform 1 0 25484 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_273
timestamp 1676037725
transform 1 0 26220 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_295
timestamp 1676037725
transform 1 0 28244 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_306
timestamp 1676037725
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_313
timestamp 1676037725
transform 1 0 29900 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_334
timestamp 1676037725
transform 1 0 31832 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_11
timestamp 1676037725
transform 1 0 2116 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_17
timestamp 1676037725
transform 1 0 2668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_33
timestamp 1676037725
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_45
timestamp 1676037725
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_53
timestamp 1676037725
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 1676037725
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_105
timestamp 1676037725
transform 1 0 10764 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_121
timestamp 1676037725
transform 1 0 12236 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_126
timestamp 1676037725
transform 1 0 12696 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_130
timestamp 1676037725
transform 1 0 13064 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_136
timestamp 1676037725
transform 1 0 13616 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_145
timestamp 1676037725
transform 1 0 14444 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_158
timestamp 1676037725
transform 1 0 15640 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_166
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_178
timestamp 1676037725
transform 1 0 17480 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_182
timestamp 1676037725
transform 1 0 17848 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_187
timestamp 1676037725
transform 1 0 18308 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_195
timestamp 1676037725
transform 1 0 19044 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_206
timestamp 1676037725
transform 1 0 20056 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_219
timestamp 1676037725
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_230
timestamp 1676037725
transform 1 0 22264 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_238
timestamp 1676037725
transform 1 0 23000 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_246
timestamp 1676037725
transform 1 0 23736 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_253
timestamp 1676037725
transform 1 0 24380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_257
timestamp 1676037725
transform 1 0 24748 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_278
timestamp 1676037725
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_303
timestamp 1676037725
transform 1 0 28980 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_334
timestamp 1676037725
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_15
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_23
timestamp 1676037725
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_37
timestamp 1676037725
transform 1 0 4508 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_45
timestamp 1676037725
transform 1 0 5244 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_61
timestamp 1676037725
transform 1 0 6716 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_73
timestamp 1676037725
transform 1 0 7820 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_81
timestamp 1676037725
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_105
timestamp 1676037725
transform 1 0 10764 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_115
timestamp 1676037725
transform 1 0 11684 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_125
timestamp 1676037725
transform 1 0 12604 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_133
timestamp 1676037725
transform 1 0 13340 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_138
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_149
timestamp 1676037725
transform 1 0 14812 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_153
timestamp 1676037725
transform 1 0 15180 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_163
timestamp 1676037725
transform 1 0 16100 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_176
timestamp 1676037725
transform 1 0 17296 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_183
timestamp 1676037725
transform 1 0 17940 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_208
timestamp 1676037725
transform 1 0 20240 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_221
timestamp 1676037725
transform 1 0 21436 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_235
timestamp 1676037725
transform 1 0 22724 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_246
timestamp 1676037725
transform 1 0 23736 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_260
timestamp 1676037725
transform 1 0 25024 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_267
timestamp 1676037725
transform 1 0 25668 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_271
timestamp 1676037725
transform 1 0 26036 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_293
timestamp 1676037725
transform 1 0 28060 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_297
timestamp 1676037725
transform 1 0 28428 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_306
timestamp 1676037725
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_331
timestamp 1676037725
transform 1 0 31556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_337
timestamp 1676037725
transform 1 0 32108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_27
timestamp 1676037725
transform 1 0 3588 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_29
timestamp 1676037725
transform 1 0 3772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_41
timestamp 1676037725
transform 1 0 4876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_53
timestamp 1676037725
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_81
timestamp 1676037725
transform 1 0 8556 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_85
timestamp 1676037725
transform 1 0 8924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_97
timestamp 1676037725
transform 1 0 10028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_109
timestamp 1676037725
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_121
timestamp 1676037725
transform 1 0 12236 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_129
timestamp 1676037725
transform 1 0 12972 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_137
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_141
timestamp 1676037725
transform 1 0 14076 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_149
timestamp 1676037725
transform 1 0 14812 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_157
timestamp 1676037725
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_161
timestamp 1676037725
transform 1 0 15916 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_166
timestamp 1676037725
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_176
timestamp 1676037725
transform 1 0 17296 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_184
timestamp 1676037725
transform 1 0 18032 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_194
timestamp 1676037725
transform 1 0 18952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_197
timestamp 1676037725
transform 1 0 19228 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_201
timestamp 1676037725
transform 1 0 19596 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_211
timestamp 1676037725
transform 1 0 20516 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_219
timestamp 1676037725
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1676037725
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_230
timestamp 1676037725
transform 1 0 22264 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_238
timestamp 1676037725
transform 1 0 23000 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_245
timestamp 1676037725
transform 1 0 23644 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_251
timestamp 1676037725
transform 1 0 24196 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_253
timestamp 1676037725
transform 1 0 24380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_258
timestamp 1676037725
transform 1 0 24840 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_265
timestamp 1676037725
transform 1 0 25484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_272
timestamp 1676037725
transform 1 0 26128 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_303
timestamp 1676037725
transform 1 0 28980 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_307
timestamp 1676037725
transform 1 0 29348 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_309
timestamp 1676037725
transform 1 0 29532 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_333
timestamp 1676037725
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 29256 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 31464 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 30820 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 25208 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1676037725
transform 1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 25208 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 24564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1676037725
transform 1 0 20700 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 17664 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 32476 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 32476 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 32476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 32476 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 32476 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 32476 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 32476 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 32476 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 32476 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 32476 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 32476 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 32476 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 32476 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 32476 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 32476 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 32476 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 32476 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 32476 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 32476 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 32476 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 32476 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 32476 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 32476 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 32476 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 32476 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 32476 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 32476 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 32476 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 32476 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 32476 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 32476 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 32476 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 32476 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 32476 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 32476 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 32476 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 26864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 29440 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 32016 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 26864 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 32016 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 24288 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 29440 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
<< labels >>
flabel metal4 s 31710 21560 31770 21760 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 32446 21560 32506 21760 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30974 21560 31034 21760 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30238 21560 30298 21760 0 FreeSans 480 90 0 0 ui_in[0]
port 3 nsew signal input
flabel metal4 s 29502 21560 29562 21760 0 FreeSans 480 90 0 0 ui_in[1]
port 4 nsew signal input
flabel metal4 s 28766 21560 28826 21760 0 FreeSans 480 90 0 0 ui_in[2]
port 5 nsew signal input
flabel metal4 s 28030 21560 28090 21760 0 FreeSans 480 90 0 0 ui_in[3]
port 6 nsew signal input
flabel metal4 s 27294 21560 27354 21760 0 FreeSans 480 90 0 0 ui_in[4]
port 7 nsew signal input
flabel metal4 s 26558 21560 26618 21760 0 FreeSans 480 90 0 0 ui_in[5]
port 8 nsew signal input
flabel metal4 s 25822 21560 25882 21760 0 FreeSans 480 90 0 0 ui_in[6]
port 9 nsew signal input
flabel metal4 s 25086 21560 25146 21760 0 FreeSans 480 90 0 0 ui_in[7]
port 10 nsew signal input
flabel metal4 s 24350 21560 24410 21760 0 FreeSans 480 90 0 0 uio_in[0]
port 11 nsew signal input
flabel metal4 s 23614 21560 23674 21760 0 FreeSans 480 90 0 0 uio_in[1]
port 12 nsew signal input
flabel metal4 s 22878 21560 22938 21760 0 FreeSans 480 90 0 0 uio_in[2]
port 13 nsew signal input
flabel metal4 s 22142 21560 22202 21760 0 FreeSans 480 90 0 0 uio_in[3]
port 14 nsew signal input
flabel metal4 s 21406 21560 21466 21760 0 FreeSans 480 90 0 0 uio_in[4]
port 15 nsew signal input
flabel metal4 s 20670 21560 20730 21760 0 FreeSans 480 90 0 0 uio_in[5]
port 16 nsew signal input
flabel metal4 s 19934 21560 19994 21760 0 FreeSans 480 90 0 0 uio_in[6]
port 17 nsew signal input
flabel metal4 s 19198 21560 19258 21760 0 FreeSans 480 90 0 0 uio_in[7]
port 18 nsew signal input
flabel metal4 s 6686 21560 6746 21760 0 FreeSans 480 90 0 0 uio_oe[0]
port 19 nsew signal tristate
flabel metal4 s 5950 21560 6010 21760 0 FreeSans 480 90 0 0 uio_oe[1]
port 20 nsew signal tristate
flabel metal4 s 5214 21560 5274 21760 0 FreeSans 480 90 0 0 uio_oe[2]
port 21 nsew signal tristate
flabel metal4 s 4478 21560 4538 21760 0 FreeSans 480 90 0 0 uio_oe[3]
port 22 nsew signal tristate
flabel metal4 s 3742 21560 3802 21760 0 FreeSans 480 90 0 0 uio_oe[4]
port 23 nsew signal tristate
flabel metal4 s 3006 21560 3066 21760 0 FreeSans 480 90 0 0 uio_oe[5]
port 24 nsew signal tristate
flabel metal4 s 2270 21560 2330 21760 0 FreeSans 480 90 0 0 uio_oe[6]
port 25 nsew signal tristate
flabel metal4 s 1534 21560 1594 21760 0 FreeSans 480 90 0 0 uio_oe[7]
port 26 nsew signal tristate
flabel metal4 s 12574 21560 12634 21760 0 FreeSans 480 90 0 0 uio_out[0]
port 27 nsew signal tristate
flabel metal4 s 11838 21560 11898 21760 0 FreeSans 480 90 0 0 uio_out[1]
port 28 nsew signal tristate
flabel metal4 s 11102 21560 11162 21760 0 FreeSans 480 90 0 0 uio_out[2]
port 29 nsew signal tristate
flabel metal4 s 10366 21560 10426 21760 0 FreeSans 480 90 0 0 uio_out[3]
port 30 nsew signal tristate
flabel metal4 s 9630 21560 9690 21760 0 FreeSans 480 90 0 0 uio_out[4]
port 31 nsew signal tristate
flabel metal4 s 8894 21560 8954 21760 0 FreeSans 480 90 0 0 uio_out[5]
port 32 nsew signal tristate
flabel metal4 s 8158 21560 8218 21760 0 FreeSans 480 90 0 0 uio_out[6]
port 33 nsew signal tristate
flabel metal4 s 7422 21560 7482 21760 0 FreeSans 480 90 0 0 uio_out[7]
port 34 nsew signal tristate
flabel metal4 s 18462 21560 18522 21760 0 FreeSans 480 90 0 0 uo_out[0]
port 35 nsew signal tristate
flabel metal4 s 17726 21560 17786 21760 0 FreeSans 480 90 0 0 uo_out[1]
port 36 nsew signal tristate
flabel metal4 s 16990 21560 17050 21760 0 FreeSans 480 90 0 0 uo_out[2]
port 37 nsew signal tristate
flabel metal4 s 16254 21560 16314 21760 0 FreeSans 480 90 0 0 uo_out[3]
port 38 nsew signal tristate
flabel metal4 s 15518 21560 15578 21760 0 FreeSans 480 90 0 0 uo_out[4]
port 39 nsew signal tristate
flabel metal4 s 14782 21560 14842 21760 0 FreeSans 480 90 0 0 uo_out[5]
port 40 nsew signal tristate
flabel metal4 s 14046 21560 14106 21760 0 FreeSans 480 90 0 0 uo_out[6]
port 41 nsew signal tristate
flabel metal4 s 13310 21560 13370 21760 0 FreeSans 480 90 0 0 uo_out[7]
port 42 nsew signal tristate
flabel metal4 s 4865 1040 5185 20720 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 12707 1040 13027 20720 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 20549 1040 20869 20720 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 28391 1040 28711 20720 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 8786 1040 9106 20720 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 16628 1040 16948 20720 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 24470 1040 24790 20720 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 32312 1040 32632 20720 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
rlabel metal1 16790 20128 16790 20128 0 vccd1
rlabel via1 16868 20672 16868 20672 0 vssd1
rlabel metal1 25346 18394 25346 18394 0 _000_
rlabel metal1 25116 18122 25116 18122 0 _001_
rlabel metal1 24955 19958 24955 19958 0 _002_
rlabel metal2 26266 19482 26266 19482 0 _003_
rlabel metal1 24564 18870 24564 18870 0 _004_
rlabel metal1 25438 18632 25438 18632 0 _005_
rlabel metal1 28290 18836 28290 18836 0 _006_
rlabel metal2 30222 20672 30222 20672 0 _007_
rlabel metal1 16192 19890 16192 19890 0 _008_
rlabel metal2 15318 20230 15318 20230 0 _009_
rlabel metal1 14306 19482 14306 19482 0 _010_
rlabel metal2 17342 19550 17342 19550 0 _011_
rlabel metal2 14398 20230 14398 20230 0 _012_
rlabel metal1 12650 19380 12650 19380 0 _013_
rlabel metal1 12190 20468 12190 20468 0 _014_
rlabel metal2 11730 18564 11730 18564 0 _015_
rlabel metal1 14260 18938 14260 18938 0 _016_
rlabel metal2 13202 19652 13202 19652 0 _017_
rlabel metal1 12374 19720 12374 19720 0 _018_
rlabel metal1 14352 19754 14352 19754 0 _019_
rlabel metal1 19320 20434 19320 20434 0 _020_
rlabel metal2 18262 19516 18262 19516 0 _021_
rlabel metal1 19274 19278 19274 19278 0 _022_
rlabel metal1 17020 19346 17020 19346 0 _023_
rlabel metal2 23414 19686 23414 19686 0 _024_
rlabel metal2 24610 20230 24610 20230 0 _025_
rlabel metal2 24426 19244 24426 19244 0 _026_
rlabel metal1 23368 18258 23368 18258 0 _027_
rlabel metal2 23138 19720 23138 19720 0 _028_
rlabel metal1 24748 19822 24748 19822 0 _029_
rlabel metal1 23046 18802 23046 18802 0 _030_
rlabel metal1 24058 18122 24058 18122 0 _031_
rlabel metal2 19734 19380 19734 19380 0 _032_
rlabel metal1 17664 18734 17664 18734 0 _033_
rlabel metal4 31740 21185 31740 21185 0 clk
rlabel metal1 30130 18258 30130 18258 0 clknet_0_clk
rlabel metal2 26358 18292 26358 18292 0 clknet_1_0__leaf_clk
rlabel metal2 30038 18564 30038 18564 0 clknet_1_1__leaf_clk
rlabel metal1 23506 19244 23506 19244 0 cnt\[0\]
rlabel metal2 23460 19278 23460 19278 0 cnt\[1\]
rlabel metal1 23414 19822 23414 19822 0 cnt\[2\]
rlabel metal1 23598 19312 23598 19312 0 cnt\[3\]
rlabel metal1 23690 18802 23690 18802 0 cnt\[4\]
rlabel metal2 23230 18462 23230 18462 0 cnt\[5\]
rlabel metal1 22678 18768 22678 18768 0 cnt\[6\]
rlabel metal2 24886 20740 24886 20740 0 cnt\[7\]
rlabel metal2 31510 18632 31510 18632 0 net1
rlabel metal1 17296 19754 17296 19754 0 net10
rlabel metal1 6394 19856 6394 19856 0 net11
rlabel metal1 19964 19890 19964 19890 0 net12
rlabel metal1 29210 18870 29210 18870 0 net13
rlabel metal2 30774 19584 30774 19584 0 net14
rlabel metal2 30866 19312 30866 19312 0 net2
rlabel metal2 25254 19924 25254 19924 0 net3
rlabel metal2 24518 20128 24518 20128 0 net4
rlabel metal2 24886 19822 24886 19822 0 net5
rlabel metal1 23506 20264 23506 20264 0 net6
rlabel metal1 21436 19482 21436 19482 0 net7
rlabel metal1 20884 18938 20884 18938 0 net8
rlabel metal1 16146 19414 16146 19414 0 net9
rlabel metal4 31004 20641 31004 20641 0 rst_n
rlabel metal1 31740 19414 31740 19414 0 rst_n_i
rlabel metal4 30268 19757 30268 19757 0 ui_in[0]
rlabel metal4 24380 20845 24380 20845 0 uio_in[0]
rlabel metal4 23644 21389 23644 21389 0 uio_in[1]
rlabel metal4 22908 21321 22908 21321 0 uio_in[2]
rlabel metal4 22172 21321 22172 21321 0 uio_in[3]
rlabel metal4 21436 21049 21436 21049 0 uio_in[4]
rlabel metal4 20700 21253 20700 21253 0 uio_in[5]
rlabel metal1 22218 20468 22218 20468 0 uio_in[6]
rlabel metal4 19228 21185 19228 21185 0 uio_in[7]
rlabel via2 6578 20043 6578 20043 0 uio_oe[0]
rlabel via2 5842 20043 5842 20043 0 uio_oe[1]
rlabel metal1 5198 20026 5198 20026 0 uio_oe[2]
rlabel via2 4370 20043 4370 20043 0 uio_oe[3]
rlabel via2 3910 19499 3910 19499 0 uio_oe[4]
rlabel via2 3082 20043 3082 20043 0 uio_oe[5]
rlabel via2 2254 20043 2254 20043 0 uio_oe[6]
rlabel via2 2438 19499 2438 19499 0 uio_oe[7]
rlabel via2 12742 20587 12742 20587 0 uio_out[0]
rlabel via2 11914 19499 11914 19499 0 uio_out[1]
rlabel via2 12006 20587 12006 20587 0 uio_out[2]
rlabel metal1 11316 18938 11316 18938 0 uio_out[3]
rlabel via2 10994 19499 10994 19499 0 uio_out[4]
rlabel metal1 9844 20026 9844 20026 0 uio_out[5]
rlabel metal4 8188 21049 8188 21049 0 uio_out[6]
rlabel metal4 7452 20777 7452 20777 0 uio_out[7]
rlabel via2 18722 20587 18722 20587 0 uo_out[0]
rlabel metal1 18078 19278 18078 19278 0 uo_out[1]
rlabel metal2 17802 20723 17802 20723 0 uo_out[2]
rlabel via2 16146 19499 16146 19499 0 uo_out[3]
rlabel metal1 16882 18938 16882 18938 0 uo_out[4]
rlabel metal1 15088 20570 15088 20570 0 uo_out[5]
rlabel metal1 13662 20026 13662 20026 0 uo_out[6]
rlabel metal4 13340 20437 13340 20437 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 33580 21760
<< end >>
