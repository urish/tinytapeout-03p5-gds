magic
tech sky130A
magscale 1 2
timestamp 1685205181
<< nwell >>
rect 1066 19845 32514 20411
rect 1066 18757 32514 19323
rect 1066 17669 32514 18235
rect 1066 16581 32514 17147
rect 1066 15493 32514 16059
rect 1066 14405 32514 14971
rect 1066 13317 32514 13883
rect 1066 12229 32514 12795
rect 1066 11141 32514 11707
rect 1066 10053 32514 10619
rect 1066 8965 32514 9531
rect 1066 7877 32514 8443
rect 1066 6789 32514 7355
rect 1066 5701 32514 6267
rect 1066 4613 32514 5179
rect 1066 3525 32514 4091
rect 1066 2437 32514 3003
rect 1066 1349 32514 1915
<< obsli1 >>
rect 1104 1071 32476 20689
<< obsm1 >>
rect 1104 1040 32632 21072
<< obsm2 >>
rect 2226 1051 32626 21185
<< obsm3 >>
rect 1526 1055 32630 21181
<< metal4 >>
rect 1534 19548 1594 21760
rect 2270 20092 2330 21760
rect 3006 20092 3066 21760
rect 3742 19548 3802 21760
rect 4478 20092 4538 21760
rect 5214 20908 5274 21760
rect 4865 1040 5185 20720
rect 5950 20092 6010 21760
rect 6686 20092 6746 21760
rect 7422 19956 7482 21760
rect 8158 20500 8218 21760
rect 8894 20908 8954 21760
rect 8786 1040 9106 20720
rect 9630 19548 9690 21760
rect 10366 19004 10426 21760
rect 11102 20636 11162 21760
rect 11838 19548 11898 21760
rect 12574 20636 12634 21760
rect 12707 1040 13027 20720
rect 13310 19276 13370 21760
rect 14046 20092 14106 21760
rect 14782 20636 14842 21760
rect 15518 19004 15578 21760
rect 16254 19548 16314 21760
rect 16990 20908 17050 21760
rect 16628 1040 16948 20720
rect 17726 19412 17786 21760
rect 18462 20636 18522 21760
rect 19198 20772 19258 21760
rect 19934 21180 19994 21760
rect 20670 20908 20730 21760
rect 20549 1040 20869 20720
rect 21406 20500 21466 21760
rect 22142 21044 22202 21760
rect 22878 21044 22938 21760
rect 23614 21180 23674 21760
rect 24350 20030 24410 21760
rect 25086 21560 25146 21760
rect 25822 21560 25882 21760
rect 26558 21560 26618 21760
rect 27294 21560 27354 21760
rect 28030 21560 28090 21760
rect 28766 21560 28826 21760
rect 29502 21560 29562 21760
rect 24470 1040 24790 20720
rect 28391 1040 28711 20720
rect 30238 17916 30298 21760
rect 30974 19684 31034 21760
rect 31710 20772 31770 21760
rect 32446 21560 32506 21760
rect 32312 1040 32632 20720
<< obsm4 >>
rect 1674 20012 2190 21181
rect 2410 20012 2926 21181
rect 3146 20012 3662 21181
rect 1674 19468 3662 20012
rect 3882 20012 4398 21181
rect 4618 20828 5134 21181
rect 5354 20828 5870 21181
rect 4618 20800 5870 20828
rect 4618 20012 4785 20800
rect 3882 19468 4785 20012
rect 1531 17851 4785 19468
rect 5265 20012 5870 20800
rect 6090 20012 6606 21181
rect 6826 20012 7342 21181
rect 5265 19876 7342 20012
rect 7562 20420 8078 21181
rect 8298 20828 8814 21181
rect 9034 20828 9550 21181
rect 8298 20800 9550 20828
rect 8298 20420 8706 20800
rect 7562 19876 8706 20420
rect 5265 17851 8706 19876
rect 9186 19468 9550 20800
rect 9770 19468 10286 21181
rect 9186 18924 10286 19468
rect 10506 20556 11022 21181
rect 11242 20556 11758 21181
rect 10506 19468 11758 20556
rect 11978 20556 12494 21181
rect 12714 20800 13230 21181
rect 11978 19468 12627 20556
rect 10506 18924 12627 19468
rect 9186 17851 12627 18924
rect 13107 19196 13230 20800
rect 13450 20012 13966 21181
rect 14186 20556 14702 21181
rect 14922 20556 15438 21181
rect 14186 20012 15438 20556
rect 13450 19196 15438 20012
rect 13107 18924 15438 19196
rect 15658 19468 16174 21181
rect 16394 20828 16910 21181
rect 17130 20828 17646 21181
rect 16394 20800 17646 20828
rect 16394 19468 16548 20800
rect 15658 18924 16548 19468
rect 13107 17851 16548 18924
rect 17028 19332 17646 20800
rect 17866 20556 18382 21181
rect 18602 20692 19118 21181
rect 19338 21100 19854 21181
rect 20074 21100 20590 21181
rect 19338 20828 20590 21100
rect 20810 20828 21326 21181
rect 19338 20800 21326 20828
rect 19338 20692 20469 20800
rect 18602 20556 20469 20692
rect 17866 19332 20469 20556
rect 17028 17851 20469 19332
rect 20949 20420 21326 20800
rect 21546 20964 22062 21181
rect 22282 20964 22798 21181
rect 23018 21100 23534 21181
rect 23754 21100 24270 21181
rect 23018 20964 24270 21100
rect 21546 20420 24270 20964
rect 20949 19950 24270 20420
rect 24490 20800 30158 21181
rect 20949 17851 24390 19950
rect 24870 17851 28311 20800
rect 28791 17851 30158 20800
rect 30378 19604 30894 21181
rect 31114 20692 31630 21181
rect 31114 19604 31773 20692
rect 30378 17851 31773 19604
<< labels >>
rlabel metal4 s 31710 20772 31770 21760 6 clk
port 1 nsew signal input
rlabel metal4 s 32446 21560 32506 21760 6 ena
port 2 nsew signal input
rlabel metal4 s 30974 19684 31034 21760 6 rst_n
port 3 nsew signal input
rlabel metal4 s 30238 17916 30298 21760 6 ui_in[0]
port 4 nsew signal input
rlabel metal4 s 29502 21560 29562 21760 6 ui_in[1]
port 5 nsew signal input
rlabel metal4 s 28766 21560 28826 21760 6 ui_in[2]
port 6 nsew signal input
rlabel metal4 s 28030 21560 28090 21760 6 ui_in[3]
port 7 nsew signal input
rlabel metal4 s 27294 21560 27354 21760 6 ui_in[4]
port 8 nsew signal input
rlabel metal4 s 26558 21560 26618 21760 6 ui_in[5]
port 9 nsew signal input
rlabel metal4 s 25822 21560 25882 21760 6 ui_in[6]
port 10 nsew signal input
rlabel metal4 s 25086 21560 25146 21760 6 ui_in[7]
port 11 nsew signal input
rlabel metal4 s 24350 20030 24410 21760 6 uio_in[0]
port 12 nsew signal input
rlabel metal4 s 23614 21180 23674 21760 6 uio_in[1]
port 13 nsew signal input
rlabel metal4 s 22878 21044 22938 21760 6 uio_in[2]
port 14 nsew signal input
rlabel metal4 s 22142 21044 22202 21760 6 uio_in[3]
port 15 nsew signal input
rlabel metal4 s 21406 20500 21466 21760 6 uio_in[4]
port 16 nsew signal input
rlabel metal4 s 20670 20908 20730 21760 6 uio_in[5]
port 17 nsew signal input
rlabel metal4 s 19934 21180 19994 21760 6 uio_in[6]
port 18 nsew signal input
rlabel metal4 s 19198 20772 19258 21760 6 uio_in[7]
port 19 nsew signal input
rlabel metal4 s 6686 20092 6746 21760 6 uio_oe[0]
port 20 nsew signal output
rlabel metal4 s 5950 20092 6010 21760 6 uio_oe[1]
port 21 nsew signal output
rlabel metal4 s 5214 20908 5274 21760 6 uio_oe[2]
port 22 nsew signal output
rlabel metal4 s 4478 20092 4538 21760 6 uio_oe[3]
port 23 nsew signal output
rlabel metal4 s 3742 19548 3802 21760 6 uio_oe[4]
port 24 nsew signal output
rlabel metal4 s 3006 20092 3066 21760 6 uio_oe[5]
port 25 nsew signal output
rlabel metal4 s 2270 20092 2330 21760 6 uio_oe[6]
port 26 nsew signal output
rlabel metal4 s 1534 19548 1594 21760 6 uio_oe[7]
port 27 nsew signal output
rlabel metal4 s 12574 20636 12634 21760 6 uio_out[0]
port 28 nsew signal output
rlabel metal4 s 11838 19548 11898 21760 6 uio_out[1]
port 29 nsew signal output
rlabel metal4 s 11102 20636 11162 21760 6 uio_out[2]
port 30 nsew signal output
rlabel metal4 s 10366 19004 10426 21760 6 uio_out[3]
port 31 nsew signal output
rlabel metal4 s 9630 19548 9690 21760 6 uio_out[4]
port 32 nsew signal output
rlabel metal4 s 8894 20908 8954 21760 6 uio_out[5]
port 33 nsew signal output
rlabel metal4 s 8158 20500 8218 21760 6 uio_out[6]
port 34 nsew signal output
rlabel metal4 s 7422 19956 7482 21760 6 uio_out[7]
port 35 nsew signal output
rlabel metal4 s 18462 20636 18522 21760 6 uo_out[0]
port 36 nsew signal output
rlabel metal4 s 17726 19412 17786 21760 6 uo_out[1]
port 37 nsew signal output
rlabel metal4 s 16990 20908 17050 21760 6 uo_out[2]
port 38 nsew signal output
rlabel metal4 s 16254 19548 16314 21760 6 uo_out[3]
port 39 nsew signal output
rlabel metal4 s 15518 19004 15578 21760 6 uo_out[4]
port 40 nsew signal output
rlabel metal4 s 14782 20636 14842 21760 6 uo_out[5]
port 41 nsew signal output
rlabel metal4 s 14046 20092 14106 21760 6 uo_out[6]
port 42 nsew signal output
rlabel metal4 s 13310 19276 13370 21760 6 uo_out[7]
port 43 nsew signal output
rlabel metal4 s 4865 1040 5185 20720 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s 12707 1040 13027 20720 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s 20549 1040 20869 20720 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s 28391 1040 28711 20720 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s 8786 1040 9106 20720 6 vssd1
port 45 nsew ground bidirectional
rlabel metal4 s 16628 1040 16948 20720 6 vssd1
port 45 nsew ground bidirectional
rlabel metal4 s 24470 1040 24790 20720 6 vssd1
port 45 nsew ground bidirectional
rlabel metal4 s 32312 1040 32632 20720 6 vssd1
port 45 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 33580 21760
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 627928
string GDS_FILE /home/uri/p/tinytapeout-03p5-gds/openlane/tt_um_test/runs/23_05_27_19_31/results/signoff/tt_um_test.magic.gds
string GDS_START 178412
<< end >>

