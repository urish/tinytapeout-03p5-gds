magic
tech sky130A
magscale 1 2
timestamp 1684775844
<< viali >>
rect 5917 9673 5951 9707
rect 7665 9673 7699 9707
rect 8493 9673 8527 9707
rect 16221 9673 16255 9707
rect 54677 9673 54711 9707
rect 58265 9673 58299 9707
rect 59277 9673 59311 9707
rect 60013 9673 60047 9707
rect 60841 9673 60875 9707
rect 63417 9673 63451 9707
rect 66177 9673 66211 9707
rect 66913 9673 66947 9707
rect 69811 9673 69845 9707
rect 90373 9673 90407 9707
rect 93501 9673 93535 9707
rect 95985 9673 96019 9707
rect 96905 9673 96939 9707
rect 98193 9673 98227 9707
rect 100677 9673 100711 9707
rect 103713 9673 103747 9707
rect 104725 9673 104759 9707
rect 105461 9673 105495 9707
rect 108865 9673 108899 9707
rect 111349 9673 111383 9707
rect 122665 9673 122699 9707
rect 125241 9673 125275 9707
rect 127909 9673 127943 9707
rect 128829 9673 128863 9707
rect 129565 9673 129599 9707
rect 131497 9673 131531 9707
rect 133521 9673 133555 9707
rect 134257 9673 134291 9707
rect 153393 9673 153427 9707
rect 156153 9673 156187 9707
rect 156889 9673 156923 9707
rect 157625 9673 157659 9707
rect 158729 9673 158763 9707
rect 160201 9673 160235 9707
rect 161949 9673 161983 9707
rect 165629 9673 165663 9707
rect 192585 9673 192619 9707
rect 193413 9673 193447 9707
rect 194885 9673 194919 9707
rect 196357 9673 196391 9707
rect 197369 9673 197403 9707
rect 198841 9673 198875 9707
rect 200037 9673 200071 9707
rect 202521 9673 202555 9707
rect 203257 9673 203291 9707
rect 207489 9673 207523 9707
rect 212641 9673 212675 9707
rect 225705 9673 225739 9707
rect 229845 9673 229879 9707
rect 233525 9673 233559 9707
rect 234353 9673 234387 9707
rect 235089 9673 235123 9707
rect 255697 9673 255731 9707
rect 260021 9673 260055 9707
rect 262413 9673 262447 9707
rect 262873 9673 262907 9707
rect 263333 9673 263367 9707
rect 267841 9673 267875 9707
rect 1685 9605 1719 9639
rect 2421 9605 2455 9639
rect 3249 9605 3283 9639
rect 4353 9605 4387 9639
rect 5089 9605 5123 9639
rect 5825 9605 5859 9639
rect 6837 9605 6871 9639
rect 7573 9605 7607 9639
rect 8401 9605 8435 9639
rect 11989 9605 12023 9639
rect 12725 9605 12759 9639
rect 13553 9605 13587 9639
rect 14657 9605 14691 9639
rect 15393 9605 15427 9639
rect 16129 9605 16163 9639
rect 17141 9605 17175 9639
rect 17325 9605 17359 9639
rect 17877 9605 17911 9639
rect 18613 9605 18647 9639
rect 18797 9605 18831 9639
rect 25513 9605 25547 9639
rect 26617 9605 26651 9639
rect 130577 9605 130611 9639
rect 172345 9605 172379 9639
rect 172529 9605 172563 9639
rect 173081 9605 173115 9639
rect 175841 9605 175875 9639
rect 176669 9605 176703 9639
rect 240241 9605 240275 9639
rect 261033 9605 261067 9639
rect 4537 9537 4571 9571
rect 9689 9537 9723 9571
rect 23765 9537 23799 9571
rect 23857 9537 23891 9571
rect 25145 9537 25179 9571
rect 26433 9537 26467 9571
rect 27997 9537 28031 9571
rect 28641 9537 28675 9571
rect 29745 9537 29779 9571
rect 32413 9537 32447 9571
rect 35633 9537 35667 9571
rect 36277 9537 36311 9571
rect 36921 9537 36955 9571
rect 38117 9537 38151 9571
rect 38853 9537 38887 9571
rect 39497 9537 39531 9571
rect 40785 9537 40819 9571
rect 41429 9537 41463 9571
rect 42073 9537 42107 9571
rect 43269 9537 43303 9571
rect 44005 9537 44039 9571
rect 44649 9537 44683 9571
rect 45937 9537 45971 9571
rect 46581 9537 46615 9571
rect 47225 9537 47259 9571
rect 48421 9537 48455 9571
rect 49157 9537 49191 9571
rect 49801 9537 49835 9571
rect 50629 9537 50663 9571
rect 51365 9537 51399 9571
rect 52101 9537 52135 9571
rect 53021 9537 53055 9571
rect 53849 9537 53883 9571
rect 54493 9537 54527 9571
rect 58081 9537 58115 9571
rect 59093 9537 59127 9571
rect 59829 9537 59863 9571
rect 60657 9537 60691 9571
rect 63233 9537 63267 9571
rect 65993 9537 66027 9571
rect 66729 9537 66763 9571
rect 69121 9537 69155 9571
rect 69581 9537 69615 9571
rect 72157 9537 72191 9571
rect 72433 9537 72467 9571
rect 74733 9537 74767 9571
rect 77309 9537 77343 9571
rect 79885 9537 79919 9571
rect 82461 9537 82495 9571
rect 84577 9537 84611 9571
rect 86785 9537 86819 9571
rect 89269 9537 89303 9571
rect 90189 9537 90223 9571
rect 93317 9537 93351 9571
rect 94789 9537 94823 9571
rect 95801 9537 95835 9571
rect 96721 9537 96755 9571
rect 98009 9537 98043 9571
rect 99297 9537 99331 9571
rect 99481 9537 99515 9571
rect 100493 9537 100527 9571
rect 103253 9537 103287 9571
rect 103897 9537 103931 9571
rect 104909 9537 104943 9571
rect 105645 9537 105679 9571
rect 106381 9537 106415 9571
rect 107761 9537 107795 9571
rect 108405 9537 108439 9571
rect 109049 9537 109083 9571
rect 110061 9537 110095 9571
rect 110797 9537 110831 9571
rect 111533 9537 111567 9571
rect 112913 9537 112947 9571
rect 113557 9537 113591 9571
rect 114201 9537 114235 9571
rect 115213 9537 115247 9571
rect 115949 9537 115983 9571
rect 116685 9537 116719 9571
rect 118065 9537 118099 9571
rect 118709 9537 118743 9571
rect 119353 9537 119387 9571
rect 120365 9537 120399 9571
rect 121101 9537 121135 9571
rect 121745 9537 121779 9571
rect 122481 9537 122515 9571
rect 125057 9537 125091 9571
rect 127725 9537 127759 9571
rect 128645 9537 128679 9571
rect 129381 9537 129415 9571
rect 130209 9537 130243 9571
rect 130393 9537 130427 9571
rect 131313 9537 131347 9571
rect 133337 9537 133371 9571
rect 134073 9537 134107 9571
rect 138121 9537 138155 9571
rect 138765 9537 138799 9571
rect 139409 9537 139443 9571
rect 140697 9537 140731 9571
rect 141341 9537 141375 9571
rect 141985 9537 142019 9571
rect 143273 9537 143307 9571
rect 143917 9537 143951 9571
rect 144561 9537 144595 9571
rect 145849 9537 145883 9571
rect 146493 9537 146527 9571
rect 147137 9537 147171 9571
rect 148425 9537 148459 9571
rect 149069 9537 149103 9571
rect 149713 9537 149747 9571
rect 151001 9537 151035 9571
rect 151645 9537 151679 9571
rect 152289 9537 152323 9571
rect 153577 9537 153611 9571
rect 154221 9537 154255 9571
rect 154865 9537 154899 9571
rect 155969 9537 156003 9571
rect 156705 9537 156739 9571
rect 157441 9537 157475 9571
rect 158545 9537 158579 9571
rect 159281 9537 159315 9571
rect 160017 9537 160051 9571
rect 161305 9537 161339 9571
rect 162317 9537 162351 9571
rect 163973 9537 164007 9571
rect 164341 9537 164375 9571
rect 165445 9537 165479 9571
rect 166457 9537 166491 9571
rect 167285 9537 167319 9571
rect 168113 9537 168147 9571
rect 171701 9537 171735 9571
rect 174461 9537 174495 9571
rect 177773 9537 177807 9571
rect 179153 9537 179187 9571
rect 179429 9537 179463 9571
rect 181729 9537 181763 9571
rect 182005 9537 182039 9571
rect 184305 9537 184339 9571
rect 186881 9537 186915 9571
rect 189457 9537 189491 9571
rect 190837 9537 190871 9571
rect 192401 9537 192435 9571
rect 193229 9537 193263 9571
rect 194701 9537 194735 9571
rect 196173 9537 196207 9571
rect 197185 9537 197219 9571
rect 197921 9537 197955 9571
rect 198657 9537 198691 9571
rect 199853 9537 199887 9571
rect 202337 9537 202371 9571
rect 203073 9537 203107 9571
rect 205833 9537 205867 9571
rect 206569 9537 206603 9571
rect 207673 9537 207707 9571
rect 208317 9537 208351 9571
rect 208961 9537 208995 9571
rect 210249 9537 210283 9571
rect 210893 9537 210927 9571
rect 211537 9537 211571 9571
rect 212825 9537 212859 9571
rect 213469 9537 213503 9571
rect 214113 9537 214147 9571
rect 215401 9537 215435 9571
rect 216045 9537 216079 9571
rect 216689 9537 216723 9571
rect 217977 9537 218011 9571
rect 218621 9537 218655 9571
rect 219265 9537 219299 9571
rect 220553 9537 220587 9571
rect 221197 9537 221231 9571
rect 221841 9537 221875 9571
rect 223129 9537 223163 9571
rect 223773 9537 223807 9571
rect 224601 9537 224635 9571
rect 224785 9537 224819 9571
rect 224969 9537 225003 9571
rect 225521 9537 225555 9571
rect 228189 9537 228223 9571
rect 229661 9537 229695 9571
rect 230765 9537 230799 9571
rect 231409 9537 231443 9571
rect 233341 9537 233375 9571
rect 234169 9537 234203 9571
rect 234905 9537 234939 9571
rect 235825 9537 235859 9571
rect 236009 9537 236043 9571
rect 239689 9537 239723 9571
rect 241253 9537 241287 9571
rect 243553 9537 243587 9571
rect 246129 9537 246163 9571
rect 248705 9537 248739 9571
rect 251281 9537 251315 9571
rect 253857 9537 253891 9571
rect 255881 9537 255915 9571
rect 257905 9537 257939 9571
rect 257997 9537 258031 9571
rect 259193 9537 259227 9571
rect 259377 9537 259411 9571
rect 259837 9537 259871 9571
rect 260665 9537 260699 9571
rect 260849 9537 260883 9571
rect 261769 9537 261803 9571
rect 262229 9537 262263 9571
rect 263241 9537 263275 9571
rect 264161 9537 264195 9571
rect 264345 9537 264379 9571
rect 265173 9537 265207 9571
rect 266001 9537 266035 9571
rect 267105 9537 267139 9571
rect 268209 9537 268243 9571
rect 269497 9537 269531 9571
rect 270141 9537 270175 9571
rect 9965 9469 9999 9503
rect 12173 9469 12207 9503
rect 14841 9469 14875 9503
rect 26249 9469 26283 9503
rect 27813 9469 27847 9503
rect 53389 9469 53423 9503
rect 53665 9469 53699 9503
rect 75009 9469 75043 9503
rect 77585 9469 77619 9503
rect 80161 9469 80195 9503
rect 82737 9469 82771 9503
rect 84853 9469 84887 9503
rect 87061 9469 87095 9503
rect 89085 9469 89119 9503
rect 89821 9469 89855 9503
rect 161121 9469 161155 9503
rect 162777 9469 162811 9503
rect 164617 9469 164651 9503
rect 166273 9469 166307 9503
rect 167101 9469 167135 9503
rect 167929 9469 167963 9503
rect 169125 9469 169159 9503
rect 169401 9469 169435 9503
rect 174737 9469 174771 9503
rect 178049 9469 178083 9503
rect 184581 9469 184615 9503
rect 187157 9469 187191 9503
rect 189733 9469 189767 9503
rect 241529 9469 241563 9503
rect 243829 9469 243863 9503
rect 246405 9469 246439 9503
rect 248981 9469 249015 9503
rect 251557 9469 251591 9503
rect 254133 9469 254167 9503
rect 256433 9469 256467 9503
rect 256709 9469 256743 9503
rect 259009 9469 259043 9503
rect 261585 9469 261619 9503
rect 264989 9469 265023 9503
rect 265817 9469 265851 9503
rect 269313 9469 269347 9503
rect 270417 9469 270451 9503
rect 3433 9401 3467 9435
rect 5273 9401 5307 9435
rect 13737 9401 13771 9435
rect 15577 9401 15611 9435
rect 18061 9401 18095 9435
rect 28825 9401 28859 9435
rect 32597 9401 32631 9435
rect 48973 9401 49007 9435
rect 114017 9401 114051 9435
rect 117881 9401 117915 9435
rect 138581 9401 138615 9435
rect 141157 9401 141191 9435
rect 143733 9401 143767 9435
rect 146953 9401 146987 9435
rect 148885 9401 148919 9435
rect 154037 9401 154071 9435
rect 159465 9401 159499 9435
rect 176853 9401 176887 9435
rect 198105 9401 198139 9435
rect 218437 9401 218471 9435
rect 221013 9401 221047 9435
rect 1777 9333 1811 9367
rect 2513 9333 2547 9367
rect 6929 9333 6963 9367
rect 12817 9333 12851 9367
rect 24041 9333 24075 9367
rect 28181 9333 28215 9367
rect 29929 9333 29963 9367
rect 35449 9333 35483 9367
rect 36093 9333 36127 9367
rect 36737 9333 36771 9367
rect 37933 9333 37967 9367
rect 38669 9333 38703 9367
rect 39313 9333 39347 9367
rect 40601 9333 40635 9367
rect 41245 9333 41279 9367
rect 41889 9333 41923 9367
rect 43085 9333 43119 9367
rect 43821 9333 43855 9367
rect 44465 9333 44499 9367
rect 45753 9333 45787 9367
rect 46397 9333 46431 9367
rect 47041 9333 47075 9367
rect 48237 9333 48271 9367
rect 49617 9333 49651 9367
rect 50445 9333 50479 9367
rect 51181 9333 51215 9367
rect 51917 9333 51951 9367
rect 52837 9333 52871 9367
rect 54033 9333 54067 9367
rect 89453 9333 89487 9367
rect 94881 9333 94915 9367
rect 99665 9333 99699 9367
rect 106197 9333 106231 9367
rect 107577 9333 107611 9367
rect 108221 9333 108255 9367
rect 109877 9333 109911 9367
rect 110613 9333 110647 9367
rect 112729 9333 112763 9367
rect 113373 9333 113407 9367
rect 115029 9333 115063 9367
rect 115765 9333 115799 9367
rect 116501 9333 116535 9367
rect 118525 9333 118559 9367
rect 119169 9333 119203 9367
rect 120181 9333 120215 9367
rect 120917 9333 120951 9367
rect 121837 9333 121871 9367
rect 139225 9333 139259 9367
rect 140513 9333 140547 9367
rect 141801 9333 141835 9367
rect 143089 9333 143123 9367
rect 144377 9333 144411 9367
rect 145665 9333 145699 9367
rect 146309 9333 146343 9367
rect 148241 9333 148275 9367
rect 149529 9333 149563 9367
rect 150817 9333 150851 9367
rect 151461 9333 151495 9367
rect 152105 9333 152139 9367
rect 154681 9333 154715 9367
rect 161489 9333 161523 9367
rect 166641 9333 166675 9367
rect 167469 9333 167503 9367
rect 168297 9333 168331 9367
rect 173173 9333 173207 9367
rect 175933 9333 175967 9367
rect 190929 9333 190963 9367
rect 206385 9333 206419 9367
rect 208133 9333 208167 9367
rect 208777 9333 208811 9367
rect 210065 9333 210099 9367
rect 210709 9333 210743 9367
rect 211353 9333 211387 9367
rect 213285 9333 213319 9367
rect 213929 9333 213963 9367
rect 215217 9333 215251 9367
rect 215861 9333 215895 9367
rect 216505 9333 216539 9367
rect 217793 9333 217827 9367
rect 219081 9333 219115 9367
rect 220369 9333 220403 9367
rect 221657 9333 221691 9367
rect 222945 9333 222979 9367
rect 223589 9333 223623 9367
rect 228373 9333 228407 9367
rect 230857 9333 230891 9367
rect 231593 9333 231627 9367
rect 236193 9333 236227 9367
rect 236561 9333 236595 9367
rect 240333 9333 240367 9367
rect 258181 9333 258215 9367
rect 261953 9333 261987 9367
rect 264529 9333 264563 9367
rect 265357 9333 265391 9367
rect 266185 9333 266219 9367
rect 267197 9333 267231 9367
rect 268485 9333 268519 9367
rect 269681 9333 269715 9367
rect 1777 9129 1811 9163
rect 23213 9129 23247 9163
rect 33609 9129 33643 9163
rect 35173 9129 35207 9163
rect 53205 9129 53239 9163
rect 57529 9129 57563 9163
rect 59185 9129 59219 9163
rect 60013 9129 60047 9163
rect 62773 9129 62807 9163
rect 66361 9129 66395 9163
rect 88441 9129 88475 9163
rect 90189 9129 90223 9163
rect 96169 9129 96203 9163
rect 98009 9129 98043 9163
rect 121009 9129 121043 9163
rect 121929 9129 121963 9163
rect 123217 9129 123251 9163
rect 124597 9129 124631 9163
rect 127817 9129 127851 9163
rect 131405 9129 131439 9163
rect 156153 9129 156187 9163
rect 156981 9129 157015 9163
rect 157809 9129 157843 9163
rect 164801 9129 164835 9163
rect 170505 9129 170539 9163
rect 193597 9129 193631 9163
rect 195805 9129 195839 9163
rect 198933 9129 198967 9163
rect 200957 9129 200991 9163
rect 204085 9129 204119 9163
rect 228373 9129 228407 9163
rect 234077 9129 234111 9163
rect 234905 9129 234939 9163
rect 236837 9129 236871 9163
rect 237573 9129 237607 9163
rect 260205 9129 260239 9163
rect 261769 9129 261803 9163
rect 269083 9129 269117 9163
rect 112177 9061 112211 9095
rect 133429 9061 133463 9095
rect 134257 9061 134291 9095
rect 134901 9061 134935 9095
rect 154957 9061 154991 9095
rect 223405 9061 223439 9095
rect 264805 9061 264839 9095
rect 268393 9061 268427 9095
rect 22845 8993 22879 9027
rect 23673 8993 23707 9027
rect 27169 8993 27203 9027
rect 69581 8993 69615 9027
rect 72065 8993 72099 9027
rect 73445 8993 73479 9027
rect 74733 8993 74767 9027
rect 75009 8993 75043 9027
rect 77217 8993 77251 9027
rect 77493 8993 77527 9027
rect 78597 8993 78631 9027
rect 79885 8993 79919 9027
rect 82369 8993 82403 9027
rect 83841 8993 83875 9027
rect 89361 8993 89395 9027
rect 94973 8993 95007 9027
rect 95801 8993 95835 9027
rect 96813 8993 96847 9027
rect 97641 8993 97675 9027
rect 98469 8993 98503 9027
rect 99297 8993 99331 9027
rect 100401 8993 100435 9027
rect 128737 8993 128771 9027
rect 129289 8993 129323 9027
rect 165353 8993 165387 9027
rect 179613 8993 179647 9027
rect 180901 8993 180935 9027
rect 182189 8993 182223 9027
rect 182465 8993 182499 9027
rect 184305 8993 184339 9027
rect 185593 8993 185627 9027
rect 186881 8993 186915 9027
rect 189457 8993 189491 9027
rect 197277 8993 197311 9027
rect 224325 8993 224359 9027
rect 230029 8993 230063 9027
rect 231041 8993 231075 9027
rect 241989 8993 242023 9027
rect 243461 8993 243495 9027
rect 254133 8993 254167 9027
rect 256433 8993 256467 9027
rect 257721 8993 257755 9027
rect 263977 8993 264011 9027
rect 267933 8993 267967 9027
rect 268853 8993 268887 9027
rect 3157 8925 3191 8959
rect 8309 8925 8343 8959
rect 10517 8925 10551 8959
rect 11253 8925 11287 8959
rect 13461 8925 13495 8959
rect 23029 8925 23063 8959
rect 23857 8925 23891 8959
rect 26893 8925 26927 8959
rect 28917 8925 28951 8959
rect 29009 8925 29043 8959
rect 30113 8925 30147 8959
rect 30205 8925 30239 8959
rect 31125 8925 31159 8959
rect 31217 8925 31251 8959
rect 31953 8925 31987 8959
rect 32045 8925 32079 8959
rect 32229 8925 32263 8959
rect 33425 8925 33459 8959
rect 40325 8925 40359 8959
rect 45477 8925 45511 8959
rect 53021 8925 53055 8959
rect 53757 8925 53791 8959
rect 53941 8925 53975 8959
rect 54585 8925 54619 8959
rect 54769 8925 54803 8959
rect 55505 8925 55539 8959
rect 55689 8925 55723 8959
rect 56425 8925 56459 8959
rect 56517 8925 56551 8959
rect 57161 8925 57195 8959
rect 57345 8925 57379 8959
rect 58081 8925 58115 8959
rect 58173 8925 58207 8959
rect 58909 8925 58943 8959
rect 59001 8925 59035 8959
rect 59645 8925 59679 8959
rect 59829 8925 59863 8959
rect 60749 8925 60783 8959
rect 60933 8925 60967 8959
rect 61577 8925 61611 8959
rect 61761 8925 61795 8959
rect 62405 8925 62439 8959
rect 62589 8925 62623 8959
rect 63233 8925 63267 8959
rect 63417 8925 63451 8959
rect 64061 8925 64095 8959
rect 64245 8925 64279 8959
rect 64981 8925 65015 8959
rect 65073 8925 65107 8959
rect 65993 8925 66027 8959
rect 66177 8925 66211 8959
rect 66821 8925 66855 8959
rect 67097 8925 67131 8959
rect 69857 8925 69891 8959
rect 72341 8925 72375 8959
rect 73721 8925 73755 8959
rect 78873 8925 78907 8959
rect 80161 8925 80195 8959
rect 82645 8925 82679 8959
rect 84117 8925 84151 8959
rect 85405 8925 85439 8959
rect 86509 8925 86543 8959
rect 88257 8925 88291 8959
rect 88993 8925 89027 8959
rect 89177 8925 89211 8959
rect 89913 8925 89947 8959
rect 90005 8925 90039 8959
rect 90741 8925 90775 8959
rect 90833 8925 90867 8959
rect 91661 8925 91695 8959
rect 91845 8925 91879 8959
rect 92489 8925 92523 8959
rect 92673 8925 92707 8959
rect 93409 8925 93443 8959
rect 93501 8925 93535 8959
rect 93685 8925 93719 8959
rect 94145 8925 94179 8959
rect 94329 8925 94363 8959
rect 95157 8925 95191 8959
rect 95985 8925 96019 8959
rect 96997 8925 97031 8959
rect 97825 8925 97859 8959
rect 98653 8925 98687 8959
rect 99481 8925 99515 8959
rect 100125 8925 100159 8959
rect 107209 8925 107243 8959
rect 112361 8925 112395 8959
rect 117513 8925 117547 8959
rect 120825 8925 120859 8959
rect 121653 8925 121687 8959
rect 121745 8925 121779 8959
rect 122665 8925 122699 8959
rect 122757 8925 122791 8959
rect 123401 8925 123435 8959
rect 123585 8925 123619 8959
rect 124229 8925 124263 8959
rect 124413 8925 124447 8959
rect 125057 8925 125091 8959
rect 125241 8925 125275 8959
rect 125885 8925 125919 8959
rect 126069 8925 126103 8959
rect 126713 8925 126747 8959
rect 126897 8925 126931 8959
rect 127633 8925 127667 8959
rect 128369 8925 128403 8959
rect 128553 8925 128587 8959
rect 129565 8925 129599 8959
rect 131037 8925 131071 8959
rect 131221 8925 131255 8959
rect 131865 8925 131899 8959
rect 132049 8925 132083 8959
rect 133061 8925 133095 8959
rect 133245 8925 133279 8959
rect 133981 8925 134015 8959
rect 134073 8925 134107 8959
rect 134717 8925 134751 8959
rect 139777 8925 139811 8959
rect 144929 8925 144963 8959
rect 150081 8925 150115 8959
rect 155141 8925 155175 8959
rect 155785 8925 155819 8959
rect 155969 8925 156003 8959
rect 156705 8925 156739 8959
rect 156797 8925 156831 8959
rect 157533 8925 157567 8959
rect 157625 8925 157659 8959
rect 158637 8925 158671 8959
rect 159833 8925 159867 8959
rect 160201 8925 160235 8959
rect 160845 8925 160879 8959
rect 161213 8925 161247 8959
rect 161857 8925 161891 8959
rect 162225 8925 162259 8959
rect 162593 8925 162627 8959
rect 163789 8925 163823 8959
rect 165169 8925 165203 8959
rect 166641 8925 166675 8959
rect 167929 8925 167963 8959
rect 168113 8925 168147 8959
rect 169033 8925 169067 8959
rect 170321 8925 170355 8959
rect 174093 8925 174127 8959
rect 177497 8925 177531 8959
rect 179889 8925 179923 8959
rect 181177 8925 181211 8959
rect 184581 8925 184615 8959
rect 185869 8925 185903 8959
rect 187157 8925 187191 8959
rect 189733 8925 189767 8959
rect 190653 8925 190687 8959
rect 190745 8925 190779 8959
rect 191573 8925 191607 8959
rect 191757 8925 191791 8959
rect 192493 8925 192527 8959
rect 192585 8925 192619 8959
rect 193321 8925 193355 8959
rect 193413 8925 193447 8959
rect 194609 8925 194643 8959
rect 194793 8925 194827 8959
rect 195529 8925 195563 8959
rect 195621 8925 195655 8959
rect 196265 8925 196299 8959
rect 196449 8925 196483 8959
rect 197553 8925 197587 8959
rect 198657 8925 198691 8959
rect 198749 8925 198783 8959
rect 199761 8925 199795 8959
rect 199945 8925 199979 8959
rect 200589 8925 200623 8959
rect 200773 8925 200807 8959
rect 201417 8925 201451 8959
rect 201601 8925 201635 8959
rect 202061 8925 202095 8959
rect 202245 8925 202279 8959
rect 203073 8925 203107 8959
rect 203257 8925 203291 8959
rect 203441 8925 203475 8959
rect 203901 8925 203935 8959
rect 211721 8925 211755 8959
rect 216873 8925 216907 8959
rect 222025 8925 222059 8959
rect 223221 8925 223255 8959
rect 224049 8925 224083 8959
rect 224141 8925 224175 8959
rect 225613 8925 225647 8959
rect 225705 8925 225739 8959
rect 226441 8925 226475 8959
rect 226533 8925 226567 8959
rect 227269 8925 227303 8959
rect 227361 8925 227395 8959
rect 228097 8925 228131 8959
rect 228189 8925 228223 8959
rect 228833 8925 228867 8959
rect 229017 8925 229051 8959
rect 229661 8925 229695 8959
rect 229845 8925 229879 8959
rect 230765 8925 230799 8959
rect 232053 8925 232087 8959
rect 232237 8925 232271 8959
rect 232881 8925 232915 8959
rect 233065 8925 233099 8959
rect 233709 8925 233743 8959
rect 233893 8925 233927 8959
rect 234537 8925 234571 8959
rect 234721 8925 234755 8959
rect 235825 8925 235859 8959
rect 236009 8925 236043 8959
rect 236193 8925 236227 8959
rect 236653 8925 236687 8959
rect 237389 8925 237423 8959
rect 242265 8925 242299 8959
rect 243737 8925 243771 8959
rect 244749 8925 244783 8959
rect 245025 8925 245059 8959
rect 246129 8925 246163 8959
rect 246405 8925 246439 8959
rect 247417 8925 247451 8959
rect 247693 8925 247727 8959
rect 248705 8925 248739 8959
rect 248981 8925 249015 8959
rect 251281 8925 251315 8959
rect 251557 8925 251591 8959
rect 252569 8925 252603 8959
rect 252845 8925 252879 8959
rect 253857 8925 253891 8959
rect 256709 8925 256743 8959
rect 257997 8925 258031 8959
rect 263701 8925 263735 8959
rect 268025 8925 268059 8959
rect 270141 8925 270175 8959
rect 270417 8925 270451 8959
rect 3341 8857 3375 8891
rect 8493 8857 8527 8891
rect 10701 8857 10735 8891
rect 25145 8857 25179 8891
rect 26065 8857 26099 8891
rect 32781 8857 32815 8891
rect 85589 8857 85623 8891
rect 159189 8857 159223 8891
rect 164157 8857 164191 8891
rect 167285 8857 167319 8891
rect 169677 8857 169711 8891
rect 176761 8857 176795 8891
rect 259101 8857 259135 8891
rect 260113 8857 260147 8891
rect 261677 8857 261711 8891
rect 262597 8857 262631 8891
rect 265265 8857 265299 8891
rect 266829 8857 266863 8891
rect 11345 8789 11379 8823
rect 13553 8789 13587 8823
rect 24041 8789 24075 8823
rect 25237 8789 25271 8823
rect 26157 8789 26191 8823
rect 29193 8789 29227 8823
rect 30389 8789 30423 8823
rect 31401 8789 31435 8823
rect 32873 8789 32907 8823
rect 40141 8789 40175 8823
rect 45293 8789 45327 8823
rect 54125 8789 54159 8823
rect 54953 8789 54987 8823
rect 55873 8789 55907 8823
rect 56701 8789 56735 8823
rect 58357 8789 58391 8823
rect 61117 8789 61151 8823
rect 61945 8789 61979 8823
rect 63601 8789 63635 8823
rect 64429 8789 64463 8823
rect 65257 8789 65291 8823
rect 86601 8789 86635 8823
rect 91017 8789 91051 8823
rect 92029 8789 92063 8823
rect 92857 8789 92891 8823
rect 94513 8789 94547 8823
rect 95341 8789 95375 8823
rect 97181 8789 97215 8823
rect 98837 8789 98871 8823
rect 99665 8789 99699 8823
rect 107025 8789 107059 8823
rect 117329 8789 117363 8823
rect 122941 8789 122975 8823
rect 123769 8789 123803 8823
rect 125425 8789 125459 8823
rect 126253 8789 126287 8823
rect 127081 8789 127115 8823
rect 132233 8789 132267 8823
rect 135453 8789 135487 8823
rect 139593 8789 139627 8823
rect 144745 8789 144779 8823
rect 149897 8789 149931 8823
rect 155509 8789 155543 8823
rect 168297 8789 168331 8823
rect 170229 8789 170263 8823
rect 174185 8789 174219 8823
rect 176853 8789 176887 8823
rect 177589 8789 177623 8823
rect 190929 8789 190963 8823
rect 191205 8789 191239 8823
rect 191941 8789 191975 8823
rect 192769 8789 192803 8823
rect 194977 8789 195011 8823
rect 196633 8789 196667 8823
rect 200129 8789 200163 8823
rect 201785 8789 201819 8823
rect 202429 8789 202463 8823
rect 202705 8789 202739 8823
rect 211537 8789 211571 8823
rect 216689 8789 216723 8823
rect 221841 8789 221875 8823
rect 225889 8789 225923 8823
rect 226717 8789 226751 8823
rect 227545 8789 227579 8823
rect 229201 8789 229235 8823
rect 232421 8789 232455 8823
rect 233249 8789 233283 8823
rect 236561 8789 236595 8823
rect 259193 8789 259227 8823
rect 262689 8789 262723 8823
rect 265357 8789 265391 8823
rect 266921 8789 266955 8823
rect 23489 8585 23523 8619
rect 25237 8585 25271 8619
rect 28733 8585 28767 8619
rect 29653 8585 29687 8619
rect 30481 8585 30515 8619
rect 31309 8585 31343 8619
rect 32689 8585 32723 8619
rect 54125 8585 54159 8619
rect 54769 8585 54803 8619
rect 55505 8585 55539 8619
rect 56241 8585 56275 8619
rect 57069 8585 57103 8619
rect 58633 8585 58667 8619
rect 59829 8585 59863 8619
rect 60749 8585 60783 8619
rect 61577 8585 61611 8619
rect 62313 8585 62347 8619
rect 63785 8585 63819 8619
rect 64613 8585 64647 8619
rect 88993 8585 89027 8619
rect 91109 8585 91143 8619
rect 91845 8585 91879 8619
rect 92581 8585 92615 8619
rect 94605 8585 94639 8619
rect 95341 8585 95375 8619
rect 96813 8585 96847 8619
rect 97457 8585 97491 8619
rect 98653 8585 98687 8619
rect 100217 8585 100251 8619
rect 100861 8585 100895 8619
rect 121929 8585 121963 8619
rect 123217 8585 123251 8619
rect 123953 8585 123987 8619
rect 125609 8585 125643 8619
rect 126345 8585 126379 8619
rect 127081 8585 127115 8619
rect 128001 8585 128035 8619
rect 129473 8585 129507 8619
rect 131589 8585 131623 8619
rect 132325 8585 132359 8619
rect 134533 8585 134567 8619
rect 156889 8585 156923 8619
rect 158361 8585 158395 8619
rect 159373 8585 159407 8619
rect 165169 8585 165203 8619
rect 169953 8585 169987 8619
rect 190561 8585 190595 8619
rect 191297 8585 191331 8619
rect 192217 8585 192251 8619
rect 193597 8585 193631 8619
rect 194241 8585 194275 8619
rect 195621 8585 195655 8619
rect 196633 8585 196667 8619
rect 197553 8585 197587 8619
rect 197921 8585 197955 8619
rect 198841 8585 198875 8619
rect 199485 8585 199519 8619
rect 200865 8585 200899 8619
rect 201601 8585 201635 8619
rect 202705 8585 202739 8619
rect 203533 8585 203567 8619
rect 225981 8585 226015 8619
rect 226717 8585 226751 8619
rect 228281 8585 228315 8619
rect 229109 8585 229143 8619
rect 231041 8585 231075 8619
rect 231961 8585 231995 8619
rect 233433 8585 233467 8619
rect 234905 8585 234939 8619
rect 236009 8585 236043 8619
rect 236653 8585 236687 8619
rect 258273 8585 258307 8619
rect 262597 8585 262631 8619
rect 263241 8585 263275 8619
rect 268393 8585 268427 8619
rect 25789 8517 25823 8551
rect 26157 8517 26191 8551
rect 27261 8517 27295 8551
rect 67005 8517 67039 8551
rect 266093 8517 266127 8551
rect 266737 8517 266771 8551
rect 23305 8449 23339 8483
rect 23857 8449 23891 8483
rect 24041 8449 24075 8483
rect 25053 8449 25087 8483
rect 26433 8449 26467 8483
rect 26617 8449 26651 8483
rect 28457 8449 28491 8483
rect 28549 8449 28583 8483
rect 29469 8449 29503 8483
rect 30297 8449 30331 8483
rect 31125 8449 31159 8483
rect 32505 8449 32539 8483
rect 53941 8449 53975 8483
rect 54585 8449 54619 8483
rect 55321 8449 55355 8483
rect 56057 8449 56091 8483
rect 56885 8449 56919 8483
rect 58449 8449 58483 8483
rect 59737 8449 59771 8483
rect 60565 8449 60599 8483
rect 61393 8449 61427 8483
rect 62129 8449 62163 8483
rect 63601 8449 63635 8483
rect 64429 8449 64463 8483
rect 65257 8449 65291 8483
rect 66821 8449 66855 8483
rect 71329 8449 71363 8483
rect 74273 8449 74307 8483
rect 76481 8449 76515 8483
rect 76757 8449 76791 8483
rect 79425 8449 79459 8483
rect 81633 8449 81667 8483
rect 88809 8449 88843 8483
rect 89913 8449 89947 8483
rect 90925 8449 90959 8483
rect 91661 8449 91695 8483
rect 92397 8449 92431 8483
rect 93225 8449 93259 8483
rect 93317 8449 93351 8483
rect 94421 8449 94455 8483
rect 95157 8449 95191 8483
rect 96445 8449 96479 8483
rect 96629 8449 96663 8483
rect 97273 8449 97307 8483
rect 98469 8449 98503 8483
rect 99941 8449 99975 8483
rect 100033 8449 100067 8483
rect 100677 8449 100711 8483
rect 121285 8449 121319 8483
rect 121561 8449 121595 8483
rect 121745 8449 121779 8483
rect 123033 8449 123067 8483
rect 123769 8449 123803 8483
rect 125425 8449 125459 8483
rect 126161 8449 126195 8483
rect 126897 8449 126931 8483
rect 127633 8449 127667 8483
rect 127817 8449 127851 8483
rect 129105 8449 129139 8483
rect 129289 8449 129323 8483
rect 130761 8449 130795 8483
rect 130945 8449 130979 8483
rect 131405 8449 131439 8483
rect 132141 8449 132175 8483
rect 132969 8449 133003 8483
rect 133153 8449 133187 8483
rect 134257 8449 134291 8483
rect 134349 8449 134383 8483
rect 156705 8449 156739 8483
rect 158177 8449 158211 8483
rect 159189 8449 159223 8483
rect 160017 8449 160051 8483
rect 161213 8449 161247 8483
rect 162501 8449 162535 8483
rect 163329 8449 163363 8483
rect 163697 8449 163731 8483
rect 164985 8449 165019 8483
rect 166825 8449 166859 8483
rect 168297 8449 168331 8483
rect 169769 8449 169803 8483
rect 183293 8449 183327 8483
rect 186973 8449 187007 8483
rect 187249 8449 187283 8483
rect 188445 8449 188479 8483
rect 188721 8449 188755 8483
rect 190377 8449 190411 8483
rect 191113 8449 191147 8483
rect 192033 8449 192067 8483
rect 193229 8449 193263 8483
rect 193413 8449 193447 8483
rect 194057 8449 194091 8483
rect 195437 8449 195471 8483
rect 196449 8449 196483 8483
rect 197369 8449 197403 8483
rect 198657 8449 198691 8483
rect 199301 8449 199335 8483
rect 200681 8449 200715 8483
rect 201417 8449 201451 8483
rect 202521 8449 202555 8483
rect 203349 8449 203383 8483
rect 224417 8449 224451 8483
rect 224601 8449 224635 8483
rect 225061 8449 225095 8483
rect 225797 8449 225831 8483
rect 226533 8449 226567 8483
rect 228097 8449 228131 8483
rect 228925 8449 228959 8483
rect 230029 8449 230063 8483
rect 230673 8449 230707 8483
rect 230857 8449 230891 8483
rect 231777 8449 231811 8483
rect 233249 8449 233283 8483
rect 234537 8449 234571 8483
rect 234721 8449 234755 8483
rect 235733 8449 235767 8483
rect 235825 8449 235859 8483
rect 236469 8449 236503 8483
rect 246405 8449 246439 8483
rect 246681 8449 246715 8483
rect 249349 8449 249383 8483
rect 251557 8449 251591 8483
rect 254501 8449 254535 8483
rect 256709 8449 256743 8483
rect 258089 8449 258123 8483
rect 259193 8449 259227 8483
rect 260205 8449 260239 8483
rect 261309 8449 261343 8483
rect 261677 8449 261711 8483
rect 262505 8449 262539 8483
rect 264253 8449 264287 8483
rect 265173 8449 265207 8483
rect 265541 8449 265575 8483
rect 266461 8449 266495 8483
rect 267381 8449 267415 8483
rect 267473 8449 267507 8483
rect 267749 8449 267783 8483
rect 268209 8449 268243 8483
rect 268301 8449 268335 8483
rect 268485 8449 268519 8483
rect 268577 8449 268611 8483
rect 268669 8449 268703 8483
rect 269497 8449 269531 8483
rect 24225 8381 24259 8415
rect 24593 8381 24627 8415
rect 24869 8381 24903 8415
rect 26249 8381 26283 8415
rect 32321 8381 32355 8415
rect 33149 8381 33183 8415
rect 53757 8381 53791 8415
rect 60381 8381 60415 8415
rect 66637 8381 66671 8415
rect 67465 8381 67499 8415
rect 71605 8381 71639 8415
rect 74549 8381 74583 8415
rect 79701 8381 79735 8415
rect 81909 8381 81943 8415
rect 89453 8381 89487 8415
rect 89729 8381 89763 8415
rect 130577 8381 130611 8415
rect 156521 8381 156555 8415
rect 157993 8381 158027 8415
rect 159005 8381 159039 8415
rect 159833 8381 159867 8415
rect 161673 8381 161707 8415
rect 162317 8381 162351 8415
rect 163973 8381 164007 8415
rect 164801 8381 164835 8415
rect 167101 8381 167135 8415
rect 168481 8381 168515 8415
rect 169585 8381 169619 8415
rect 183569 8381 183603 8415
rect 196265 8381 196299 8415
rect 197185 8381 197219 8415
rect 198473 8381 198507 8415
rect 202337 8381 202371 8415
rect 202981 8381 203015 8415
rect 203165 8381 203199 8415
rect 223865 8381 223899 8415
rect 224233 8381 224267 8415
rect 229845 8381 229879 8415
rect 249625 8381 249659 8415
rect 251833 8381 251867 8415
rect 254777 8381 254811 8415
rect 256985 8381 257019 8415
rect 259009 8381 259043 8415
rect 260021 8381 260055 8415
rect 263517 8381 263551 8415
rect 269313 8381 269347 8415
rect 269681 8381 269715 8415
rect 270141 8381 270175 8415
rect 270417 8381 270451 8415
rect 65441 8313 65475 8347
rect 162133 8313 162167 8347
rect 225245 8313 225279 8347
rect 230213 8313 230247 8347
rect 264437 8313 264471 8347
rect 27353 8245 27387 8279
rect 90097 8245 90131 8279
rect 93501 8245 93535 8279
rect 133337 8245 133371 8279
rect 160201 8245 160235 8279
rect 162685 8245 162719 8279
rect 259377 8245 259411 8279
rect 260389 8245 260423 8279
rect 267197 8245 267231 8279
rect 267657 8245 267691 8279
rect 25237 8041 25271 8075
rect 28365 8041 28399 8075
rect 133061 8041 133095 8075
rect 160293 8041 160327 8075
rect 162409 8041 162443 8075
rect 166365 8041 166399 8075
rect 167101 8041 167135 8075
rect 167837 8041 167871 8075
rect 169033 8041 169067 8075
rect 230857 8041 230891 8075
rect 259009 8041 259043 8075
rect 259653 8041 259687 8075
rect 260481 8041 260515 8075
rect 269681 8041 269715 8075
rect 93317 7973 93351 8007
rect 99573 7973 99607 8007
rect 107945 7973 107979 8007
rect 258365 7973 258399 8007
rect 100125 7905 100159 7939
rect 105185 7905 105219 7939
rect 105461 7905 105495 7939
rect 161397 7905 161431 7939
rect 169585 7905 169619 7939
rect 202797 7905 202831 7939
rect 216321 7905 216355 7939
rect 268209 7905 268243 7939
rect 268669 7905 268703 7939
rect 269221 7905 269255 7939
rect 270141 7905 270175 7939
rect 24961 7837 24995 7871
rect 25053 7837 25087 7871
rect 26157 7837 26191 7871
rect 26617 7837 26651 7871
rect 26709 7837 26743 7871
rect 27353 7837 27387 7871
rect 27537 7837 27571 7871
rect 28181 7837 28215 7871
rect 28917 7837 28951 7871
rect 89545 7837 89579 7871
rect 93133 7837 93167 7871
rect 99389 7837 99423 7871
rect 104541 7837 104575 7871
rect 104725 7837 104759 7871
rect 105599 7837 105633 7871
rect 105737 7837 105771 7871
rect 108957 7837 108991 7871
rect 109785 7837 109819 7871
rect 132877 7837 132911 7871
rect 160109 7837 160143 7871
rect 161584 7837 161618 7871
rect 161765 7837 161799 7871
rect 162225 7837 162259 7871
rect 163789 7837 163823 7871
rect 163881 7837 163915 7871
rect 164617 7837 164651 7871
rect 164709 7837 164743 7871
rect 165353 7837 165387 7871
rect 165537 7837 165571 7871
rect 166181 7837 166215 7871
rect 166917 7837 166951 7871
rect 167653 7837 167687 7871
rect 168849 7837 168883 7871
rect 215861 7837 215895 7871
rect 217793 7837 217827 7871
rect 219449 7837 219483 7871
rect 230673 7837 230707 7871
rect 235825 7837 235859 7871
rect 237021 7837 237055 7871
rect 237113 7837 237147 7871
rect 237849 7837 237883 7871
rect 237941 7837 237975 7871
rect 258825 7837 258859 7871
rect 259837 7837 259871 7871
rect 260297 7837 260331 7871
rect 261861 7837 261895 7871
rect 261953 7837 261987 7871
rect 262597 7837 262631 7871
rect 262781 7837 262815 7871
rect 263425 7837 263459 7871
rect 263609 7837 263643 7871
rect 264437 7837 264471 7871
rect 264989 7837 265023 7871
rect 265081 7837 265115 7871
rect 265817 7837 265851 7871
rect 265909 7837 265943 7871
rect 268301 7837 268335 7871
rect 269313 7837 269347 7871
rect 270417 7837 270451 7871
rect 107761 7769 107795 7803
rect 218713 7769 218747 7803
rect 238125 7769 238159 7803
rect 258181 7769 258215 7803
rect 267289 7769 267323 7803
rect 267657 7769 267691 7803
rect 25605 7701 25639 7735
rect 26893 7701 26927 7735
rect 27721 7701 27755 7735
rect 29101 7701 29135 7735
rect 89729 7701 89763 7735
rect 103805 7701 103839 7735
rect 104173 7701 104207 7735
rect 106381 7701 106415 7735
rect 109049 7701 109083 7735
rect 109969 7701 110003 7735
rect 164065 7701 164099 7735
rect 164893 7701 164927 7735
rect 165721 7701 165755 7735
rect 217885 7701 217919 7735
rect 218805 7701 218839 7735
rect 219541 7701 219575 7735
rect 237297 7701 237331 7735
rect 262137 7701 262171 7735
rect 262965 7701 262999 7735
rect 263793 7701 263827 7735
rect 264253 7701 264287 7735
rect 265265 7701 265299 7735
rect 266093 7701 266127 7735
rect 25605 7497 25639 7531
rect 26433 7497 26467 7531
rect 67373 7497 67407 7531
rect 109049 7497 109083 7531
rect 111717 7497 111751 7531
rect 121193 7497 121227 7531
rect 161305 7497 161339 7531
rect 162593 7497 162627 7531
rect 163329 7497 163363 7531
rect 164065 7497 164099 7531
rect 164801 7497 164835 7531
rect 165537 7497 165571 7531
rect 220369 7497 220403 7531
rect 259653 7497 259687 7531
rect 260297 7497 260331 7531
rect 261769 7497 261803 7531
rect 262505 7497 262539 7531
rect 263241 7497 263275 7531
rect 264345 7497 264379 7531
rect 265909 7497 265943 7531
rect 106105 7429 106139 7463
rect 268761 7429 268795 7463
rect 24501 7361 24535 7395
rect 25421 7361 25455 7395
rect 26249 7361 26283 7395
rect 27813 7361 27847 7395
rect 42809 7361 42843 7395
rect 67557 7361 67591 7395
rect 100217 7361 100251 7395
rect 106473 7361 106507 7395
rect 107393 7361 107427 7395
rect 108405 7361 108439 7395
rect 109601 7361 109635 7395
rect 109785 7361 109819 7395
rect 110521 7361 110555 7395
rect 112085 7361 112119 7395
rect 121377 7361 121411 7395
rect 145665 7361 145699 7395
rect 146723 7361 146757 7395
rect 151185 7361 151219 7395
rect 161121 7361 161155 7395
rect 162409 7361 162443 7395
rect 163237 7361 163271 7395
rect 163881 7361 163915 7395
rect 164617 7361 164651 7395
rect 165353 7361 165387 7395
rect 169309 7361 169343 7395
rect 214113 7361 214147 7395
rect 214481 7361 214515 7395
rect 215539 7361 215573 7395
rect 216413 7361 216447 7395
rect 217793 7361 217827 7395
rect 218713 7361 218747 7395
rect 218989 7361 219023 7395
rect 220553 7361 220587 7395
rect 221473 7361 221507 7395
rect 221590 7361 221624 7395
rect 221749 7361 221783 7395
rect 222945 7361 222979 7395
rect 223865 7361 223899 7395
rect 229753 7361 229787 7395
rect 230305 7361 230339 7395
rect 231225 7361 231259 7395
rect 232421 7361 232455 7395
rect 232605 7361 232639 7395
rect 235365 7361 235399 7395
rect 235457 7361 235491 7395
rect 236193 7361 236227 7395
rect 237297 7361 237331 7395
rect 237481 7361 237515 7395
rect 238585 7361 238619 7395
rect 259837 7361 259871 7395
rect 260481 7361 260515 7395
rect 261125 7361 261159 7395
rect 261585 7361 261619 7395
rect 262321 7361 262355 7395
rect 263057 7361 263091 7395
rect 264161 7361 264195 7395
rect 265081 7361 265115 7395
rect 265725 7361 265759 7395
rect 266553 7361 266587 7395
rect 267381 7361 267415 7395
rect 268393 7361 268427 7395
rect 269497 7361 269531 7395
rect 270141 7361 270175 7395
rect 25237 7293 25271 7327
rect 26065 7293 26099 7327
rect 106657 7293 106691 7327
rect 107531 7293 107565 7327
rect 107669 7293 107703 7327
rect 110638 7293 110672 7327
rect 110797 7293 110831 7327
rect 112637 7293 112671 7327
rect 145849 7293 145883 7327
rect 146585 7293 146619 7327
rect 146861 7293 146895 7327
rect 151369 7293 151403 7327
rect 153025 7293 153059 7327
rect 214665 7293 214699 7327
rect 215125 7293 215159 7327
rect 215401 7293 215435 7327
rect 215677 7293 215711 7327
rect 216597 7293 216631 7327
rect 217977 7293 218011 7327
rect 218851 7293 218885 7327
rect 220737 7293 220771 7327
rect 223129 7293 223163 7327
rect 223982 7293 224016 7327
rect 224141 7293 224175 7327
rect 225153 7293 225187 7327
rect 231501 7293 231535 7327
rect 236469 7293 236503 7327
rect 238401 7293 238435 7327
rect 265541 7293 265575 7327
rect 266369 7293 266403 7327
rect 267197 7293 267231 7327
rect 269313 7293 269347 7327
rect 270417 7293 270451 7327
rect 42625 7225 42659 7259
rect 43177 7225 43211 7259
rect 107117 7225 107151 7259
rect 108313 7225 108347 7259
rect 110245 7225 110279 7259
rect 111441 7225 111475 7259
rect 146309 7225 146343 7259
rect 147873 7225 147907 7259
rect 217241 7225 217275 7259
rect 218437 7225 218471 7259
rect 220001 7225 220035 7259
rect 221197 7225 221231 7259
rect 223589 7225 223623 7259
rect 224785 7225 224819 7259
rect 24685 7157 24719 7191
rect 27997 7157 28031 7191
rect 100033 7157 100067 7191
rect 108589 7157 108623 7191
rect 147505 7157 147539 7191
rect 150909 7157 150943 7191
rect 153393 7157 153427 7191
rect 169125 7157 169159 7191
rect 216321 7157 216355 7191
rect 219633 7157 219667 7191
rect 222393 7157 222427 7191
rect 229569 7157 229603 7191
rect 230397 7157 230431 7191
rect 235641 7157 235675 7191
rect 237665 7157 237699 7191
rect 238769 7157 238803 7191
rect 239137 7157 239171 7191
rect 260941 7157 260975 7191
rect 264897 7157 264931 7191
rect 266737 7157 266771 7191
rect 267565 7157 267599 7191
rect 269681 7157 269715 7191
rect 79241 6953 79275 6987
rect 79425 6953 79459 6987
rect 169585 6953 169619 6987
rect 229937 6953 229971 6987
rect 230121 6953 230155 6987
rect 100033 6885 100067 6919
rect 169769 6885 169803 6919
rect 190009 6885 190043 6919
rect 262689 6885 262723 6919
rect 93225 6817 93259 6851
rect 99573 6817 99607 6851
rect 100309 6817 100343 6851
rect 100447 6817 100481 6851
rect 108313 6817 108347 6851
rect 108773 6817 108807 6851
rect 110245 6817 110279 6851
rect 112453 6817 112487 6851
rect 113189 6817 113223 6851
rect 114569 6817 114603 6851
rect 114937 6817 114971 6851
rect 140697 6817 140731 6851
rect 141341 6817 141375 6851
rect 141617 6817 141651 6851
rect 141734 6817 141768 6851
rect 145849 6817 145883 6851
rect 146033 6817 146067 6851
rect 146493 6817 146527 6851
rect 148241 6817 148275 6851
rect 148885 6817 148919 6851
rect 149161 6817 149195 6851
rect 149299 6817 149333 6851
rect 150541 6817 150575 6851
rect 151185 6817 151219 6851
rect 151461 6817 151495 6851
rect 152381 6817 152415 6851
rect 210249 6817 210283 6851
rect 210893 6817 210927 6851
rect 212549 6817 212583 6851
rect 214389 6817 214423 6851
rect 215677 6817 215711 6851
rect 218621 6817 218655 6851
rect 219173 6817 219207 6851
rect 220185 6817 220219 6851
rect 220829 6817 220863 6851
rect 221105 6817 221139 6851
rect 221391 6817 221425 6851
rect 222669 6817 222703 6851
rect 223313 6817 223347 6851
rect 223589 6817 223623 6851
rect 225521 6817 225555 6851
rect 229569 6817 229603 6851
rect 236009 6817 236043 6851
rect 270877 6817 270911 6851
rect 25605 6749 25639 6783
rect 26525 6749 26559 6783
rect 92765 6749 92799 6783
rect 98653 6749 98687 6783
rect 99389 6749 99423 6783
rect 100585 6749 100619 6783
rect 102241 6749 102275 6783
rect 107761 6749 107795 6783
rect 108129 6749 108163 6783
rect 109049 6749 109083 6783
rect 109187 6749 109221 6783
rect 109325 6749 109359 6783
rect 140881 6749 140915 6783
rect 141893 6749 141927 6783
rect 146769 6749 146803 6783
rect 146907 6749 146941 6783
rect 147045 6749 147079 6783
rect 148425 6749 148459 6783
rect 149437 6749 149471 6783
rect 150725 6749 150759 6783
rect 151578 6749 151612 6783
rect 151737 6749 151771 6783
rect 169217 6749 169251 6783
rect 170321 6749 170355 6783
rect 190193 6749 190227 6783
rect 210433 6749 210467 6783
rect 211169 6749 211203 6783
rect 211307 6749 211341 6783
rect 211445 6749 211479 6783
rect 217977 6749 218011 6783
rect 218161 6749 218195 6783
rect 218897 6749 218931 6783
rect 219035 6749 219069 6783
rect 220369 6749 220403 6783
rect 221243 6749 221277 6783
rect 222393 6749 222427 6783
rect 222853 6749 222887 6783
rect 223727 6749 223761 6783
rect 223865 6749 223899 6783
rect 231133 6749 231167 6783
rect 235733 6749 235767 6783
rect 236745 6749 236779 6783
rect 237113 6749 237147 6783
rect 237205 6749 237239 6783
rect 261033 6749 261067 6783
rect 262229 6749 262263 6783
rect 262873 6749 262907 6783
rect 263333 6749 263367 6783
rect 264069 6749 264103 6783
rect 264805 6749 264839 6783
rect 265541 6749 265575 6783
rect 267197 6749 267231 6783
rect 267381 6749 267415 6783
rect 268117 6749 268151 6783
rect 269221 6749 269255 6783
rect 269497 6749 269531 6783
rect 270509 6749 270543 6783
rect 270693 6749 270727 6783
rect 79057 6681 79091 6715
rect 102793 6681 102827 6715
rect 112637 6681 112671 6715
rect 212733 6681 212767 6715
rect 215861 6681 215895 6715
rect 217517 6681 217551 6715
rect 225705 6681 225739 6715
rect 227361 6681 227395 6715
rect 231777 6681 231811 6715
rect 268485 6681 268519 6715
rect 25789 6613 25823 6647
rect 26709 6613 26743 6647
rect 44465 6613 44499 6647
rect 79267 6613 79301 6647
rect 99021 6613 99055 6647
rect 101229 6613 101263 6647
rect 109969 6613 110003 6647
rect 140421 6613 140455 6647
rect 142537 6613 142571 6647
rect 147689 6613 147723 6647
rect 150081 6613 150115 6647
rect 169585 6613 169619 6647
rect 170413 6613 170447 6647
rect 212089 6613 212123 6647
rect 215401 6613 215435 6647
rect 217793 6613 217827 6647
rect 219817 6613 219851 6647
rect 222025 6613 222059 6647
rect 224509 6613 224543 6647
rect 224969 6613 225003 6647
rect 227729 6613 227763 6647
rect 228097 6613 228131 6647
rect 229937 6613 229971 6647
rect 237389 6613 237423 6647
rect 260205 6613 260239 6647
rect 262045 6613 262079 6647
rect 263517 6613 263551 6647
rect 264253 6613 264287 6647
rect 264989 6613 265023 6647
rect 265725 6613 265759 6647
rect 267565 6613 267599 6647
rect 46121 6409 46155 6443
rect 46673 6409 46707 6443
rect 79609 6409 79643 6443
rect 100125 6409 100159 6443
rect 100309 6409 100343 6443
rect 181821 6409 181855 6443
rect 189197 6409 189231 6443
rect 189365 6409 189399 6443
rect 220001 6409 220035 6443
rect 263425 6409 263459 6443
rect 42809 6341 42843 6375
rect 43085 6341 43119 6375
rect 43913 6341 43947 6375
rect 45017 6341 45051 6375
rect 45293 6341 45327 6375
rect 45753 6341 45787 6375
rect 79425 6341 79459 6375
rect 119905 6341 119939 6375
rect 120105 6341 120139 6375
rect 121101 6341 121135 6375
rect 130301 6341 130335 6375
rect 152657 6341 152691 6375
rect 188997 6341 189031 6375
rect 270877 6341 270911 6375
rect 43177 6273 43211 6307
rect 43545 6273 43579 6307
rect 44465 6273 44499 6307
rect 45385 6273 45419 6307
rect 101781 6273 101815 6307
rect 106933 6273 106967 6307
rect 108773 6273 108807 6307
rect 110889 6273 110923 6307
rect 112729 6273 112763 6307
rect 120733 6273 120767 6307
rect 125149 6273 125183 6307
rect 130669 6273 130703 6307
rect 146493 6273 146527 6307
rect 148885 6273 148919 6307
rect 150817 6273 150851 6307
rect 156061 6273 156095 6307
rect 156889 6273 156923 6307
rect 181821 6273 181855 6307
rect 182005 6273 182039 6307
rect 182557 6273 182591 6307
rect 207581 6273 207615 6307
rect 214205 6273 214239 6307
rect 217793 6273 217827 6307
rect 221197 6273 221231 6307
rect 221335 6273 221369 6307
rect 221473 6273 221507 6307
rect 223037 6273 223071 6307
rect 223405 6273 223439 6307
rect 223681 6273 223715 6307
rect 225521 6273 225555 6307
rect 225889 6273 225923 6307
rect 230213 6273 230247 6307
rect 231317 6273 231351 6307
rect 236193 6273 236227 6307
rect 261217 6273 261251 6307
rect 262413 6273 262447 6307
rect 262505 6273 262539 6307
rect 263609 6273 263643 6307
rect 264253 6273 264287 6307
rect 264621 6273 264655 6307
rect 265449 6273 265483 6307
rect 266645 6273 266679 6307
rect 267841 6273 267875 6307
rect 268393 6273 268427 6307
rect 269405 6273 269439 6307
rect 270693 6273 270727 6307
rect 91569 6205 91603 6239
rect 91753 6205 91787 6239
rect 93409 6205 93443 6239
rect 101965 6205 101999 6239
rect 102241 6205 102275 6239
rect 107117 6205 107151 6239
rect 111073 6205 111107 6239
rect 119353 6205 119387 6239
rect 125425 6205 125459 6239
rect 146677 6205 146711 6239
rect 148149 6205 148183 6239
rect 149253 6205 149287 6239
rect 151001 6205 151035 6239
rect 157073 6205 157107 6239
rect 161581 6205 161615 6239
rect 207765 6205 207799 6239
rect 208409 6205 208443 6239
rect 214389 6205 214423 6239
rect 216045 6205 216079 6239
rect 217977 6205 218011 6239
rect 218437 6205 218471 6239
rect 218713 6205 218747 6239
rect 218830 6205 218864 6239
rect 218989 6205 219023 6239
rect 220277 6205 220311 6239
rect 220461 6205 220495 6239
rect 223865 6205 223899 6239
rect 231685 6205 231719 6239
rect 236469 6205 236503 6239
rect 261493 6205 261527 6239
rect 265725 6205 265759 6239
rect 266921 6205 266955 6239
rect 269681 6205 269715 6239
rect 270509 6205 270543 6239
rect 44097 6137 44131 6171
rect 46305 6137 46339 6171
rect 79057 6137 79091 6171
rect 90925 6137 90959 6171
rect 91293 6137 91327 6171
rect 99757 6137 99791 6171
rect 120273 6137 120307 6171
rect 220921 6137 220955 6171
rect 79425 6069 79459 6103
rect 100125 6069 100159 6103
rect 120089 6069 120123 6103
rect 121101 6069 121135 6103
rect 121285 6069 121319 6103
rect 156337 6069 156371 6103
rect 189181 6069 189215 6103
rect 219633 6069 219667 6103
rect 222117 6069 222151 6103
rect 230489 6069 230523 6103
rect 262689 6069 262723 6103
rect 47869 5865 47903 5899
rect 79333 5865 79367 5899
rect 180993 5865 181027 5899
rect 182925 5865 182959 5899
rect 217241 5865 217275 5899
rect 221105 5865 221139 5899
rect 221473 5865 221507 5899
rect 228465 5865 228499 5899
rect 230857 5865 230891 5899
rect 231041 5865 231075 5899
rect 232513 5865 232547 5899
rect 265541 5865 265575 5899
rect 79517 5797 79551 5831
rect 101045 5797 101079 5831
rect 111257 5797 111291 5831
rect 111533 5797 111567 5831
rect 112453 5797 112487 5831
rect 112821 5797 112855 5831
rect 115305 5797 115339 5831
rect 115673 5797 115707 5831
rect 224969 5797 225003 5831
rect 228649 5797 228683 5831
rect 270693 5797 270727 5831
rect 78965 5729 78999 5763
rect 81265 5729 81299 5763
rect 82001 5729 82035 5763
rect 87153 5729 87187 5763
rect 109049 5729 109083 5763
rect 120273 5729 120307 5763
rect 130209 5729 130243 5763
rect 143089 5729 143123 5763
rect 143273 5729 143307 5763
rect 143549 5729 143583 5763
rect 147689 5729 147723 5763
rect 148241 5729 148275 5763
rect 150081 5729 150115 5763
rect 150449 5729 150483 5763
rect 150817 5729 150851 5763
rect 153853 5729 153887 5763
rect 212825 5729 212859 5763
rect 215401 5729 215435 5763
rect 216045 5729 216079 5763
rect 216597 5729 216631 5763
rect 221841 5729 221875 5763
rect 222301 5729 222335 5763
rect 223957 5729 223991 5763
rect 224325 5729 224359 5763
rect 225521 5729 225555 5763
rect 226165 5729 226199 5763
rect 226441 5729 226475 5763
rect 229109 5729 229143 5763
rect 263149 5729 263183 5763
rect 269865 5729 269899 5763
rect 42717 5661 42751 5695
rect 43545 5661 43579 5695
rect 43637 5661 43671 5695
rect 44005 5661 44039 5695
rect 44387 5661 44421 5695
rect 46857 5661 46891 5695
rect 46949 5661 46983 5695
rect 47317 5661 47351 5695
rect 50813 5661 50847 5695
rect 51273 5661 51307 5695
rect 81449 5661 81483 5695
rect 83381 5661 83415 5695
rect 86877 5661 86911 5695
rect 92673 5661 92707 5695
rect 94513 5661 94547 5695
rect 100401 5661 100435 5695
rect 100677 5661 100711 5695
rect 100861 5661 100895 5695
rect 102149 5661 102183 5695
rect 110889 5661 110923 5695
rect 113189 5661 113223 5695
rect 115029 5661 115063 5695
rect 119077 5661 119111 5695
rect 120089 5661 120123 5695
rect 125057 5661 125091 5695
rect 129933 5661 129967 5695
rect 153393 5661 153427 5695
rect 155693 5661 155727 5695
rect 157533 5661 157567 5695
rect 157901 5661 157935 5695
rect 158637 5661 158671 5695
rect 159005 5661 159039 5695
rect 159373 5661 159407 5695
rect 161121 5661 161155 5695
rect 161213 5661 161247 5695
rect 161765 5661 161799 5695
rect 180625 5661 180659 5695
rect 180809 5661 180843 5695
rect 181637 5661 181671 5695
rect 182097 5661 182131 5695
rect 182373 5661 182407 5695
rect 212181 5661 212215 5695
rect 212549 5661 212583 5695
rect 214665 5661 214699 5695
rect 215585 5661 215619 5695
rect 216321 5661 216355 5695
rect 216459 5661 216493 5695
rect 225705 5661 225739 5695
rect 226558 5661 226592 5695
rect 226717 5661 226751 5695
rect 227729 5661 227763 5695
rect 228097 5661 228131 5695
rect 229385 5661 229419 5695
rect 231501 5661 231535 5695
rect 231685 5661 231719 5695
rect 232329 5661 232363 5695
rect 259009 5661 259043 5695
rect 260205 5661 260239 5695
rect 261677 5661 261711 5695
rect 262873 5661 262907 5695
rect 264069 5661 264103 5695
rect 264529 5661 264563 5695
rect 265265 5661 265299 5695
rect 265357 5661 265391 5695
rect 266001 5661 266035 5695
rect 266829 5661 266863 5695
rect 267197 5661 267231 5695
rect 268393 5661 268427 5695
rect 269497 5661 269531 5695
rect 269681 5661 269715 5695
rect 270325 5661 270359 5695
rect 270509 5661 270543 5695
rect 42073 5593 42107 5627
rect 50905 5593 50939 5627
rect 83565 5593 83599 5627
rect 85221 5593 85255 5627
rect 85589 5593 85623 5627
rect 92857 5593 92891 5627
rect 103161 5593 103195 5627
rect 108405 5593 108439 5627
rect 108773 5593 108807 5627
rect 109233 5593 109267 5627
rect 113373 5593 113407 5627
rect 119445 5593 119479 5627
rect 119813 5593 119847 5627
rect 121929 5593 121963 5627
rect 122573 5593 122607 5627
rect 148425 5593 148459 5627
rect 153577 5593 153611 5627
rect 155877 5593 155911 5627
rect 162133 5593 162167 5627
rect 162777 5593 162811 5627
rect 213009 5593 213043 5627
rect 222025 5593 222059 5627
rect 228465 5593 228499 5627
rect 230673 5593 230707 5627
rect 230873 5593 230907 5627
rect 231869 5593 231903 5627
rect 259377 5593 259411 5627
rect 260573 5593 260607 5627
rect 262045 5593 262079 5627
rect 268853 5593 268887 5627
rect 42165 5525 42199 5559
rect 43269 5525 43303 5559
rect 44557 5525 44591 5559
rect 46581 5525 46615 5559
rect 47685 5525 47719 5559
rect 50537 5525 50571 5559
rect 51641 5525 51675 5559
rect 51825 5525 51859 5559
rect 79333 5525 79367 5559
rect 81633 5525 81667 5559
rect 82737 5525 82771 5559
rect 83105 5525 83139 5559
rect 125149 5525 125183 5559
rect 152013 5525 152047 5559
rect 152381 5525 152415 5559
rect 152749 5525 152783 5559
rect 160201 5525 160235 5559
rect 160569 5525 160603 5559
rect 162869 5525 162903 5559
rect 180349 5525 180383 5559
rect 215309 5525 215343 5559
rect 227361 5525 227395 5559
rect 47133 5321 47167 5355
rect 53113 5321 53147 5355
rect 101137 5321 101171 5355
rect 119261 5321 119295 5355
rect 152473 5321 152507 5355
rect 157809 5321 157843 5355
rect 158177 5321 158211 5355
rect 163053 5321 163087 5355
rect 264897 5321 264931 5355
rect 267105 5321 267139 5355
rect 267749 5321 267783 5355
rect 268669 5321 268703 5355
rect 269681 5321 269715 5355
rect 37657 5253 37691 5287
rect 37933 5253 37967 5287
rect 38393 5253 38427 5287
rect 38761 5253 38795 5287
rect 43361 5253 43395 5287
rect 43637 5253 43671 5287
rect 43729 5253 43763 5287
rect 44465 5253 44499 5287
rect 45845 5253 45879 5287
rect 46121 5253 46155 5287
rect 46213 5253 46247 5287
rect 46949 5253 46983 5287
rect 50629 5253 50663 5287
rect 50905 5253 50939 5287
rect 51365 5253 51399 5287
rect 51733 5253 51767 5287
rect 80345 5253 80379 5287
rect 80713 5253 80747 5287
rect 81633 5253 81667 5287
rect 84945 5253 84979 5287
rect 86601 5253 86635 5287
rect 87705 5253 87739 5287
rect 88073 5253 88107 5287
rect 88441 5253 88475 5287
rect 89177 5253 89211 5287
rect 91293 5253 91327 5287
rect 91661 5253 91695 5287
rect 115305 5253 115339 5287
rect 150265 5253 150299 5287
rect 153301 5253 153335 5287
rect 162593 5253 162627 5287
rect 188445 5253 188479 5287
rect 189181 5253 189215 5287
rect 218253 5253 218287 5287
rect 218529 5253 218563 5287
rect 218897 5253 218931 5287
rect 219449 5253 219483 5287
rect 221105 5253 221139 5287
rect 221381 5253 221415 5287
rect 221749 5253 221783 5287
rect 224693 5253 224727 5287
rect 227545 5253 227579 5287
rect 228189 5253 228223 5287
rect 229937 5253 229971 5287
rect 231317 5253 231351 5287
rect 239413 5253 239447 5287
rect 261861 5253 261895 5287
rect 266277 5253 266311 5287
rect 270509 5253 270543 5287
rect 38025 5185 38059 5219
rect 41613 5185 41647 5219
rect 44097 5185 44131 5219
rect 46581 5185 46615 5219
rect 47961 5185 47995 5219
rect 50997 5185 51031 5219
rect 53021 5185 53055 5219
rect 80805 5185 80839 5219
rect 80897 5185 80931 5219
rect 81449 5185 81483 5219
rect 101045 5185 101079 5219
rect 107025 5185 107059 5219
rect 107163 5185 107197 5219
rect 107301 5185 107335 5219
rect 117421 5185 117455 5219
rect 120089 5185 120123 5219
rect 121009 5185 121043 5219
rect 122205 5185 122239 5219
rect 150633 5185 150667 5219
rect 161121 5185 161155 5219
rect 161581 5185 161615 5219
rect 163145 5185 163179 5219
rect 182005 5185 182039 5219
rect 182189 5185 182223 5219
rect 182557 5185 182591 5219
rect 188813 5185 188847 5219
rect 219265 5185 219299 5219
rect 222301 5185 222335 5219
rect 222853 5185 222887 5219
rect 225705 5185 225739 5219
rect 228465 5185 228499 5219
rect 230029 5185 230063 5219
rect 238677 5185 238711 5219
rect 238861 5185 238895 5219
rect 240241 5185 240275 5219
rect 260389 5185 260423 5219
rect 261677 5185 261711 5219
rect 262965 5185 262999 5219
rect 264713 5185 264747 5219
rect 266001 5185 266035 5219
rect 266093 5185 266127 5219
rect 266921 5185 266955 5219
rect 267565 5185 267599 5219
rect 268485 5185 268519 5219
rect 269497 5185 269531 5219
rect 270325 5185 270359 5219
rect 41797 5117 41831 5151
rect 42717 5117 42751 5151
rect 53757 5117 53791 5151
rect 79793 5117 79827 5151
rect 80161 5117 80195 5151
rect 83289 5117 83323 5151
rect 83841 5117 83875 5151
rect 84761 5117 84795 5151
rect 89453 5117 89487 5151
rect 89637 5117 89671 5151
rect 91753 5117 91787 5151
rect 91937 5117 91971 5151
rect 93593 5117 93627 5151
rect 106105 5117 106139 5151
rect 106289 5117 106323 5151
rect 108221 5117 108255 5151
rect 111809 5117 111843 5151
rect 111993 5117 112027 5151
rect 112729 5117 112763 5151
rect 112846 5117 112880 5151
rect 113005 5117 113039 5151
rect 115121 5117 115155 5151
rect 115581 5117 115615 5151
rect 117605 5117 117639 5151
rect 118359 5117 118393 5151
rect 118479 5117 118513 5151
rect 118617 5117 118651 5151
rect 120273 5117 120307 5151
rect 121126 5117 121160 5151
rect 121285 5117 121319 5151
rect 150817 5117 150851 5151
rect 151553 5117 151587 5151
rect 151691 5117 151725 5151
rect 151829 5117 151863 5151
rect 153117 5117 153151 5151
rect 153577 5117 153611 5151
rect 158269 5117 158303 5151
rect 158453 5117 158487 5151
rect 160017 5117 160051 5151
rect 214021 5117 214055 5151
rect 214205 5117 214239 5151
rect 215861 5117 215895 5151
rect 223037 5117 223071 5151
rect 225889 5117 225923 5151
rect 228741 5117 228775 5151
rect 260665 5117 260699 5151
rect 261493 5117 261527 5151
rect 263241 5117 263275 5151
rect 264529 5117 264563 5151
rect 266737 5117 266771 5151
rect 268301 5117 268335 5151
rect 269313 5117 269347 5151
rect 270141 5117 270175 5151
rect 38945 5049 38979 5083
rect 44649 5049 44683 5083
rect 94237 5049 94271 5083
rect 94605 5049 94639 5083
rect 94973 5049 95007 5083
rect 106749 5049 106783 5083
rect 111441 5049 111475 5083
rect 112453 5049 112487 5083
rect 118065 5049 118099 5083
rect 119905 5049 119939 5083
rect 120733 5049 120767 5083
rect 122389 5049 122423 5083
rect 151277 5049 151311 5083
rect 155417 5049 155451 5083
rect 162133 5049 162167 5083
rect 162593 5049 162627 5083
rect 182557 5049 182591 5083
rect 230949 5049 230983 5083
rect 240425 5049 240459 5083
rect 48145 4981 48179 5015
rect 51917 4981 51951 5015
rect 84301 4981 84335 5015
rect 84669 4981 84703 5015
rect 105737 4981 105771 5015
rect 107945 4981 107979 5015
rect 113649 4981 113683 5015
rect 114109 4981 114143 5015
rect 114753 4981 114787 5015
rect 121929 4981 121963 5015
rect 152749 4981 152783 5015
rect 160477 4981 160511 5015
rect 163329 4981 163363 5015
rect 189181 4981 189215 5015
rect 189365 4981 189399 5015
rect 225061 4981 225095 5015
rect 225429 4981 225463 5015
rect 231317 4981 231351 5015
rect 231501 4981 231535 5015
rect 239505 4981 239539 5015
rect 241989 4981 242023 5015
rect 242265 4981 242299 5015
rect 242633 4981 242667 5015
rect 259101 4981 259135 5015
rect 259469 4981 259503 5015
rect 259837 4981 259871 5015
rect 42625 4777 42659 4811
rect 48789 4777 48823 4811
rect 121837 4777 121871 4811
rect 155417 4777 155451 4811
rect 217057 4777 217091 4811
rect 219725 4777 219759 4811
rect 222761 4777 222795 4811
rect 223129 4777 223163 4811
rect 224693 4777 224727 4811
rect 225061 4777 225095 4811
rect 238309 4777 238343 4811
rect 238677 4777 238711 4811
rect 239965 4777 239999 4811
rect 240333 4777 240367 4811
rect 241897 4777 241931 4811
rect 253581 4777 253615 4811
rect 255789 4777 255823 4811
rect 256709 4777 256743 4811
rect 257997 4777 258031 4811
rect 263057 4777 263091 4811
rect 265173 4777 265207 4811
rect 266921 4777 266955 4811
rect 270325 4777 270359 4811
rect 270509 4777 270543 4811
rect 99481 4709 99515 4743
rect 107669 4709 107703 4743
rect 109417 4709 109451 4743
rect 110429 4709 110463 4743
rect 111625 4709 111659 4743
rect 153853 4709 153887 4743
rect 215861 4709 215895 4743
rect 217425 4709 217459 4743
rect 230765 4709 230799 4743
rect 259285 4709 259319 4743
rect 260757 4709 260791 4743
rect 269681 4709 269715 4743
rect 81725 4641 81759 4675
rect 92489 4641 92523 4675
rect 92673 4641 92707 4675
rect 94329 4641 94363 4675
rect 99941 4641 99975 4675
rect 100033 4641 100067 4675
rect 107209 4641 107243 4675
rect 107945 4641 107979 4675
rect 109785 4641 109819 4675
rect 110705 4641 110739 4675
rect 110843 4641 110877 4675
rect 114109 4641 114143 4675
rect 114293 4641 114327 4675
rect 114569 4641 114603 4675
rect 116225 4641 116259 4675
rect 118249 4641 118283 4675
rect 118893 4641 118927 4675
rect 120917 4641 120951 4675
rect 122481 4641 122515 4675
rect 122941 4641 122975 4675
rect 124597 4641 124631 4675
rect 143089 4641 143123 4675
rect 150541 4641 150575 4675
rect 151185 4641 151219 4675
rect 151737 4641 151771 4675
rect 153209 4641 153243 4675
rect 212549 4641 212583 4675
rect 215217 4641 215251 4675
rect 216413 4641 216447 4675
rect 220645 4641 220679 4675
rect 239045 4641 239079 4675
rect 241161 4641 241195 4675
rect 242817 4641 242851 4675
rect 244105 4641 244139 4675
rect 250637 4641 250671 4675
rect 251281 4641 251315 4675
rect 252201 4641 252235 4675
rect 254041 4641 254075 4675
rect 254409 4641 254443 4675
rect 259653 4641 259687 4675
rect 266185 4641 266219 4675
rect 43269 4573 43303 4607
rect 43361 4573 43395 4607
rect 47777 4573 47811 4607
rect 48619 4573 48653 4607
rect 52377 4573 52411 4607
rect 84025 4573 84059 4607
rect 85865 4573 85899 4607
rect 87889 4573 87923 4607
rect 94421 4573 94455 4607
rect 94513 4573 94547 4607
rect 94881 4573 94915 4607
rect 107025 4573 107059 4607
rect 108083 4573 108117 4607
rect 108221 4573 108255 4607
rect 109969 4573 110003 4607
rect 110981 4573 111015 4607
rect 118433 4573 118467 4607
rect 119169 4573 119203 4607
rect 119286 4573 119320 4607
rect 119445 4573 119479 4607
rect 120457 4573 120491 4607
rect 120733 4573 120767 4607
rect 150725 4573 150759 4607
rect 151461 4573 151495 4607
rect 151599 4573 151633 4607
rect 152381 4573 152415 4607
rect 153393 4573 153427 4607
rect 154129 4573 154163 4607
rect 154267 4573 154301 4607
rect 154405 4573 154439 4607
rect 155049 4573 155083 4607
rect 155969 4573 156003 4607
rect 158361 4573 158395 4607
rect 161029 4573 161063 4607
rect 212365 4573 212399 4607
rect 215401 4573 215435 4607
rect 216137 4573 216171 4607
rect 216275 4573 216309 4607
rect 222485 4573 222519 4607
rect 226533 4573 226567 4607
rect 228833 4573 228867 4607
rect 231225 4573 231259 4607
rect 231317 4573 231351 4607
rect 239229 4573 239263 4607
rect 240977 4573 241011 4607
rect 242265 4573 242299 4607
rect 242633 4573 242667 4607
rect 243921 4573 243955 4607
rect 251465 4573 251499 4607
rect 255053 4573 255087 4607
rect 257077 4573 257111 4607
rect 257261 4573 257295 4607
rect 258181 4573 258215 4607
rect 258365 4573 258399 4607
rect 259837 4573 259871 4607
rect 263241 4573 263275 4607
rect 263793 4573 263827 4607
rect 265357 4573 265391 4607
rect 265817 4573 265851 4607
rect 266001 4573 266035 4607
rect 266737 4573 266771 4607
rect 267473 4573 267507 4607
rect 267657 4573 267691 4607
rect 268209 4573 268243 4607
rect 269313 4573 269347 4607
rect 269497 4573 269531 4607
rect 41245 4505 41279 4539
rect 41337 4505 41371 4539
rect 41705 4505 41739 4539
rect 42073 4505 42107 4539
rect 43729 4505 43763 4539
rect 45201 4505 45235 4539
rect 47869 4505 47903 4539
rect 48237 4505 48271 4539
rect 52469 4505 52503 4539
rect 52837 4505 52871 4539
rect 81909 4505 81943 4539
rect 83565 4505 83599 4539
rect 84209 4505 84243 4539
rect 88073 4505 88107 4539
rect 89729 4505 89763 4539
rect 95249 4505 95283 4539
rect 99481 4505 99515 4539
rect 122665 4505 122699 4539
rect 143273 4505 143307 4539
rect 144929 4505 144963 4539
rect 145205 4505 145239 4539
rect 156153 4505 156187 4539
rect 157809 4505 157843 4539
rect 158545 4505 158579 4539
rect 160201 4505 160235 4539
rect 160569 4505 160603 4539
rect 160845 4505 160879 4539
rect 161213 4505 161247 4539
rect 162869 4505 162903 4539
rect 163145 4505 163179 4539
rect 214205 4505 214239 4539
rect 220829 4505 220863 4539
rect 225889 4505 225923 4539
rect 226257 4505 226291 4539
rect 226717 4505 226751 4539
rect 228373 4505 228407 4539
rect 228741 4505 228775 4539
rect 229569 4505 229603 4539
rect 230765 4505 230799 4539
rect 243553 4505 243587 4539
rect 244565 4505 244599 4539
rect 245117 4505 245151 4539
rect 254501 4505 254535 4539
rect 255329 4505 255363 4539
rect 258825 4505 258859 4539
rect 260481 4505 260515 4539
rect 264161 4505 264195 4539
rect 268577 4505 268611 4539
rect 270141 4505 270175 4539
rect 270341 4505 270375 4539
rect 40049 4437 40083 4471
rect 40417 4437 40451 4471
rect 40969 4437 41003 4471
rect 42257 4437 42291 4471
rect 42993 4437 43027 4471
rect 44097 4437 44131 4471
rect 44281 4437 44315 4471
rect 46949 4437 46983 4471
rect 47501 4437 47535 4471
rect 52101 4437 52135 4471
rect 53205 4437 53239 4471
rect 53389 4437 53423 4471
rect 80345 4437 80379 4471
rect 80713 4437 80747 4471
rect 81449 4437 81483 4471
rect 86509 4437 86543 4471
rect 86877 4437 86911 4471
rect 87245 4437 87279 4471
rect 87521 4437 87555 4471
rect 90097 4437 90131 4471
rect 90465 4437 90499 4471
rect 90833 4437 90867 4471
rect 100217 4437 100251 4471
rect 108865 4437 108899 4471
rect 113373 4437 113407 4471
rect 113741 4437 113775 4471
rect 120089 4437 120123 4471
rect 142445 4437 142479 4471
rect 158177 4437 158211 4471
rect 231501 4437 231535 4471
rect 239689 4437 239723 4471
rect 241621 4437 241655 4471
rect 243277 4437 243311 4471
rect 244841 4437 244875 4471
rect 245393 4437 245427 4471
rect 251925 4437 251959 4471
rect 257721 4437 257755 4471
rect 260297 4437 260331 4471
rect 267565 4437 267599 4471
rect 50077 4233 50111 4267
rect 50261 4233 50295 4267
rect 216781 4233 216815 4267
rect 265081 4233 265115 4267
rect 268761 4233 268795 4267
rect 40049 4165 40083 4199
rect 40601 4165 40635 4199
rect 40969 4165 41003 4199
rect 41337 4165 41371 4199
rect 41705 4165 41739 4199
rect 48145 4165 48179 4199
rect 48973 4165 49007 4199
rect 49249 4165 49283 4199
rect 49341 4165 49375 4199
rect 49709 4165 49743 4199
rect 50997 4165 51031 4199
rect 51733 4165 51767 4199
rect 52101 4165 52135 4199
rect 53021 4165 53055 4199
rect 81633 4165 81667 4199
rect 84945 4165 84979 4199
rect 147505 4165 147539 4199
rect 157809 4165 157843 4199
rect 158085 4165 158119 4199
rect 161305 4165 161339 4199
rect 190009 4165 190043 4199
rect 226717 4165 226751 4199
rect 235641 4165 235675 4199
rect 240425 4165 240459 4199
rect 242265 4165 242299 4199
rect 243921 4165 243955 4199
rect 252109 4165 252143 4199
rect 254041 4165 254075 4199
rect 255697 4165 255731 4199
rect 259653 4165 259687 4199
rect 260205 4165 260239 4199
rect 260941 4165 260975 4199
rect 25789 4097 25823 4131
rect 40877 4097 40911 4131
rect 47869 4097 47903 4131
rect 51273 4097 51307 4131
rect 51365 4097 51399 4131
rect 53205 4097 53239 4131
rect 84761 4097 84795 4131
rect 86601 4097 86635 4131
rect 86969 4097 87003 4131
rect 94329 4097 94363 4131
rect 104909 4097 104943 4131
rect 105829 4097 105863 4131
rect 107209 4097 107243 4131
rect 108405 4097 108439 4131
rect 112361 4097 112395 4131
rect 113557 4097 113591 4131
rect 114201 4097 114235 4131
rect 114661 4097 114695 4131
rect 115581 4097 115615 4131
rect 145021 4097 145055 4131
rect 151921 4097 151955 4131
rect 152657 4097 152691 4131
rect 154589 4097 154623 4131
rect 158453 4097 158487 4131
rect 159189 4097 159223 4131
rect 159465 4097 159499 4131
rect 190377 4097 190411 4131
rect 209329 4097 209363 4131
rect 209789 4097 209823 4131
rect 212825 4097 212859 4131
rect 214021 4097 214055 4131
rect 214941 4097 214975 4131
rect 215861 4097 215895 4131
rect 216137 4097 216171 4131
rect 224049 4097 224083 4131
rect 226165 4097 226199 4131
rect 230397 4097 230431 4131
rect 240793 4097 240827 4131
rect 254593 4097 254627 4131
rect 264621 4097 264655 4131
rect 265265 4097 265299 4131
rect 265909 4097 265943 4131
rect 266553 4097 266587 4131
rect 267197 4097 267231 4131
rect 267657 4097 267691 4131
rect 268577 4097 268611 4131
rect 269313 4097 269347 4131
rect 270049 4097 270083 4131
rect 270785 4097 270819 4131
rect 270877 4097 270911 4131
rect 81449 4029 81483 4063
rect 83289 4029 83323 4063
rect 94513 4029 94547 4063
rect 96169 4029 96203 4063
rect 99389 4029 99423 4063
rect 99573 4029 99607 4063
rect 101229 4029 101263 4063
rect 105093 4029 105127 4063
rect 105553 4029 105587 4063
rect 105967 4029 106001 4063
rect 106105 4029 106139 4063
rect 107393 4029 107427 4063
rect 108129 4029 108163 4063
rect 108267 4029 108301 4063
rect 112545 4029 112579 4063
rect 113281 4029 113315 4063
rect 113419 4029 113453 4063
rect 114845 4029 114879 4063
rect 115698 4029 115732 4063
rect 115857 4029 115891 4063
rect 117513 4029 117547 4063
rect 117697 4029 117731 4063
rect 117973 4029 118007 4063
rect 121745 4029 121779 4063
rect 121929 4029 121963 4063
rect 123585 4029 123619 4063
rect 141801 4029 141835 4063
rect 141985 4029 142019 4063
rect 142261 4029 142295 4063
rect 145665 4029 145699 4063
rect 145849 4029 145883 4063
rect 147965 4029 147999 4063
rect 148149 4029 148183 4063
rect 149805 4029 149839 4063
rect 151737 4029 151771 4063
rect 152381 4029 152415 4063
rect 152795 4029 152829 4063
rect 152933 4029 152967 4063
rect 153577 4029 153611 4063
rect 154865 4029 154899 4063
rect 158269 4029 158303 4063
rect 158913 4029 158947 4063
rect 159327 4029 159361 4063
rect 160109 4029 160143 4063
rect 161121 4029 161155 4063
rect 162961 4029 162995 4063
rect 163329 4029 163363 4063
rect 163697 4029 163731 4063
rect 207489 4029 207523 4063
rect 207673 4029 207707 4063
rect 209973 4029 210007 4063
rect 211629 4029 211663 4063
rect 213009 4029 213043 4063
rect 213469 4029 213503 4063
rect 213745 4029 213779 4063
rect 213862 4029 213896 4063
rect 215125 4029 215159 4063
rect 215585 4029 215619 4063
rect 215999 4029 216033 4063
rect 224325 4029 224359 4063
rect 224509 4029 224543 4063
rect 225245 4029 225279 4063
rect 225362 4029 225396 4063
rect 225521 4029 225555 4063
rect 228097 4029 228131 4063
rect 228281 4029 228315 4063
rect 229109 4029 229143 4063
rect 230213 4029 230247 4063
rect 252017 4029 252051 4063
rect 252937 4029 252971 4063
rect 253949 4029 253983 4063
rect 256525 4029 256559 4063
rect 256709 4029 256743 4063
rect 257629 4029 257663 4063
rect 257813 4029 257847 4063
rect 259101 4029 259135 4063
rect 261217 4029 261251 4063
rect 268393 4029 268427 4063
rect 80805 3961 80839 3995
rect 81173 3961 81207 3995
rect 84485 3961 84519 3995
rect 107853 3961 107887 3995
rect 113005 3961 113039 3995
rect 115305 3961 115339 3995
rect 121101 3961 121135 3995
rect 121469 3961 121503 3995
rect 143917 3961 143951 3995
rect 206477 3961 206511 3995
rect 206845 3961 206879 3995
rect 224969 3961 225003 3995
rect 230581 3961 230615 3995
rect 235917 3961 235951 3995
rect 244197 3961 244231 3995
rect 252569 3961 252603 3995
rect 254961 3961 254995 3995
rect 255329 3961 255363 3995
rect 256065 3961 256099 3995
rect 260481 3961 260515 3995
rect 265725 3961 265759 3995
rect 267013 3961 267047 3995
rect 267841 3961 267875 3995
rect 25973 3893 26007 3927
rect 41889 3893 41923 3927
rect 52285 3893 52319 3927
rect 83933 3893 83967 3927
rect 98653 3893 98687 3927
rect 101597 3893 101631 3927
rect 104081 3893 104115 3927
rect 104541 3893 104575 3927
rect 106749 3893 106783 3927
rect 109049 3893 109083 3927
rect 116501 3893 116535 3927
rect 116777 3893 116811 3927
rect 117145 3893 117179 3927
rect 119997 3893 120031 3927
rect 123953 3893 123987 3927
rect 141433 3893 141467 3927
rect 147873 3893 147907 3927
rect 155417 3893 155451 3927
rect 160569 3893 160603 3927
rect 211997 3893 212031 3927
rect 212733 3893 212767 3927
rect 214665 3893 214699 3927
rect 226809 3893 226843 3927
rect 227453 3893 227487 3927
rect 242541 3893 242575 3927
rect 250821 3893 250855 3927
rect 251189 3893 251223 3927
rect 251557 3893 251591 3927
rect 257169 3893 257203 3927
rect 258273 3893 258307 3927
rect 258549 3893 258583 3927
rect 259929 3893 259963 3927
rect 264437 3893 264471 3927
rect 266369 3893 266403 3927
rect 269497 3893 269531 3927
rect 270233 3893 270267 3927
rect 67189 3689 67223 3723
rect 88165 3689 88199 3723
rect 104265 3689 104299 3723
rect 116777 3689 116811 3723
rect 157533 3689 157567 3723
rect 160201 3689 160235 3723
rect 217057 3689 217091 3723
rect 222577 3689 222611 3723
rect 227361 3689 227395 3723
rect 260573 3689 260607 3723
rect 265357 3689 265391 3723
rect 266001 3689 266035 3723
rect 267197 3689 267231 3723
rect 268485 3689 268519 3723
rect 270049 3689 270083 3723
rect 270693 3689 270727 3723
rect 37749 3621 37783 3655
rect 42533 3621 42567 3655
rect 47961 3621 47995 3655
rect 99113 3621 99147 3655
rect 119813 3621 119847 3655
rect 121009 3621 121043 3655
rect 143733 3621 143767 3655
rect 144929 3621 144963 3655
rect 147229 3621 147263 3655
rect 159005 3621 159039 3655
rect 210065 3621 210099 3655
rect 215861 3621 215895 3655
rect 269313 3621 269347 3655
rect 24961 3553 24995 3587
rect 82829 3553 82863 3587
rect 83197 3553 83231 3587
rect 94053 3553 94087 3587
rect 96629 3553 96663 3587
rect 97273 3553 97307 3587
rect 97549 3553 97583 3587
rect 97687 3553 97721 3587
rect 101321 3553 101355 3587
rect 103805 3553 103839 3587
rect 104633 3553 104667 3587
rect 105369 3553 105403 3587
rect 107025 3553 107059 3587
rect 109141 3553 109175 3587
rect 110521 3553 110555 3587
rect 115581 3553 115615 3587
rect 115857 3553 115891 3587
rect 115995 3553 116029 3587
rect 119169 3553 119203 3587
rect 120089 3553 120123 3587
rect 120365 3553 120399 3587
rect 143089 3553 143123 3587
rect 144009 3553 144043 3587
rect 144147 3553 144181 3587
rect 145389 3553 145423 3587
rect 146033 3553 146067 3587
rect 146585 3553 146619 3587
rect 155693 3553 155727 3587
rect 156337 3553 156371 3587
rect 156613 3553 156647 3587
rect 156730 3553 156764 3587
rect 156889 3553 156923 3587
rect 158361 3553 158395 3587
rect 159281 3553 159315 3587
rect 159557 3553 159591 3587
rect 207213 3553 207247 3587
rect 207673 3553 207707 3587
rect 209329 3553 209363 3587
rect 210525 3553 210559 3587
rect 210709 3553 210743 3587
rect 212457 3553 212491 3587
rect 213101 3553 213135 3587
rect 215217 3553 215251 3587
rect 216137 3553 216171 3587
rect 216254 3553 216288 3587
rect 218897 3553 218931 3587
rect 225521 3553 225555 3587
rect 226165 3553 226199 3587
rect 226579 3553 226613 3587
rect 259285 3553 259319 3587
rect 25145 3485 25179 3519
rect 25789 3485 25823 3519
rect 26525 3485 26559 3519
rect 27261 3485 27295 3519
rect 36737 3485 36771 3519
rect 36829 3485 36863 3519
rect 67097 3485 67131 3519
rect 83473 3485 83507 3519
rect 87981 3485 88015 3519
rect 91753 3485 91787 3519
rect 95893 3485 95927 3519
rect 96813 3485 96847 3519
rect 97825 3485 97859 3519
rect 99481 3485 99515 3519
rect 101965 3485 101999 3519
rect 114937 3485 114971 3519
rect 115121 3485 115155 3519
rect 116133 3485 116167 3519
rect 119353 3485 119387 3519
rect 120206 3485 120240 3519
rect 122573 3485 122607 3519
rect 138949 3485 138983 3519
rect 143273 3485 143307 3519
rect 144285 3485 144319 3519
rect 145573 3485 145607 3519
rect 146309 3485 146343 3519
rect 146447 3485 146481 3519
rect 148241 3485 148275 3519
rect 155233 3485 155267 3519
rect 155877 3485 155911 3519
rect 158545 3485 158579 3519
rect 159419 3485 159453 3519
rect 160845 3485 160879 3519
rect 204913 3485 204947 3519
rect 212641 3485 212675 3519
rect 213377 3485 213411 3519
rect 213494 3485 213528 3519
rect 213653 3485 213687 3519
rect 215401 3485 215435 3519
rect 216413 3485 216447 3519
rect 217517 3485 217551 3519
rect 222761 3485 222795 3519
rect 225705 3485 225739 3519
rect 226441 3485 226475 3519
rect 226717 3485 226751 3519
rect 230673 3485 230707 3519
rect 252109 3485 252143 3519
rect 258089 3485 258123 3519
rect 259009 3485 259043 3519
rect 265541 3485 265575 3519
rect 266185 3485 266219 3519
rect 267381 3485 267415 3519
rect 268025 3485 268059 3519
rect 268669 3485 268703 3519
rect 269129 3485 269163 3519
rect 269865 3485 269899 3519
rect 270601 3485 270635 3519
rect 37197 3417 37231 3451
rect 40233 3417 40267 3451
rect 40877 3417 40911 3451
rect 41521 3417 41555 3451
rect 41613 3417 41647 3451
rect 41981 3417 42015 3451
rect 42349 3417 42383 3451
rect 46673 3417 46707 3451
rect 46949 3417 46983 3451
rect 47041 3417 47075 3451
rect 47409 3417 47443 3451
rect 83657 3417 83691 3451
rect 85313 3417 85347 3451
rect 91937 3417 91971 3451
rect 93593 3417 93627 3451
rect 94237 3417 94271 3451
rect 99665 3417 99699 3451
rect 102149 3417 102183 3451
rect 104817 3417 104851 3451
rect 109325 3417 109359 3451
rect 139133 3417 139167 3451
rect 140789 3417 140823 3451
rect 148425 3417 148459 3451
rect 150081 3417 150115 3451
rect 161029 3417 161063 3451
rect 162685 3417 162719 3451
rect 205097 3417 205131 3451
rect 206753 3417 206787 3451
rect 207397 3417 207431 3451
rect 212365 3417 212399 3451
rect 217701 3417 217735 3451
rect 256433 3417 256467 3451
rect 258457 3417 258491 3451
rect 259929 3417 259963 3451
rect 260297 3417 260331 3451
rect 25329 3349 25363 3383
rect 25973 3349 26007 3383
rect 26709 3349 26743 3383
rect 27445 3349 27479 3383
rect 35909 3349 35943 3383
rect 36461 3349 36495 3383
rect 37565 3349 37599 3383
rect 40325 3349 40359 3383
rect 41245 3349 41279 3383
rect 46121 3349 46155 3383
rect 47777 3349 47811 3383
rect 85681 3349 85715 3383
rect 89085 3349 89119 3383
rect 98469 3349 98503 3383
rect 98745 3349 98779 3383
rect 122849 3349 122883 3383
rect 138673 3349 138707 3383
rect 155417 3349 155451 3383
rect 160569 3349 160603 3383
rect 203901 3349 203935 3383
rect 204269 3349 204303 3383
rect 214297 3349 214331 3383
rect 214665 3349 214699 3383
rect 217425 3349 217459 3383
rect 227729 3349 227763 3383
rect 230857 3349 230891 3383
rect 252385 3349 252419 3383
rect 258733 3349 258767 3383
rect 259653 3349 259687 3383
rect 267841 3349 267875 3383
rect 83289 3145 83323 3179
rect 84025 3145 84059 3179
rect 98745 3145 98779 3179
rect 101505 3145 101539 3179
rect 139593 3145 139627 3179
rect 144653 3145 144687 3179
rect 147505 3145 147539 3179
rect 211905 3145 211939 3179
rect 214481 3145 214515 3179
rect 214849 3145 214883 3179
rect 217241 3145 217275 3179
rect 218713 3145 218747 3179
rect 223865 3145 223899 3179
rect 268577 3145 268611 3179
rect 37841 3077 37875 3111
rect 38117 3077 38151 3111
rect 38209 3077 38243 3111
rect 38577 3077 38611 3111
rect 38945 3077 38979 3111
rect 39865 3077 39899 3111
rect 40141 3077 40175 3111
rect 40601 3077 40635 3111
rect 40969 3077 41003 3111
rect 86141 3077 86175 3111
rect 96629 3077 96663 3111
rect 110429 3077 110463 3111
rect 120641 3077 120675 3111
rect 121009 3077 121043 3111
rect 123217 3077 123251 3111
rect 123493 3077 123527 3111
rect 140697 3077 140731 3111
rect 157809 3077 157843 3111
rect 159741 3077 159775 3111
rect 225981 3077 226015 3111
rect 226073 3077 226107 3111
rect 259837 3077 259871 3111
rect 24317 3009 24351 3043
rect 25421 3009 25455 3043
rect 26249 3009 26283 3043
rect 27537 3009 27571 3043
rect 27997 3009 28031 3043
rect 40233 3009 40267 3043
rect 82369 3009 82403 3043
rect 86601 3009 86635 3043
rect 89177 3009 89211 3043
rect 91937 3009 91971 3043
rect 92305 3009 92339 3043
rect 94237 3009 94271 3043
rect 96077 3009 96111 3043
rect 96905 3009 96939 3043
rect 97089 3009 97123 3043
rect 98101 3009 98135 3043
rect 99665 3009 99699 3043
rect 101689 3009 101723 3043
rect 102627 3009 102661 3043
rect 102885 3009 102919 3043
rect 107117 3009 107151 3043
rect 110245 3009 110279 3043
rect 112085 3009 112119 3043
rect 116501 3009 116535 3043
rect 121377 3009 121411 3043
rect 137753 3009 137787 3043
rect 138673 3009 138707 3043
rect 142997 3009 143031 3043
rect 143733 3009 143767 3043
rect 145849 3009 145883 3043
rect 146585 3009 146619 3043
rect 146861 3009 146895 3043
rect 147965 3009 147999 3043
rect 148885 3009 148919 3043
rect 149161 3009 149195 3043
rect 155969 3009 156003 3043
rect 156889 3009 156923 3043
rect 157006 3009 157040 3043
rect 158821 3009 158855 3043
rect 158938 3009 158972 3043
rect 160201 3009 160235 3043
rect 160569 3009 160603 3043
rect 161213 3009 161247 3043
rect 162961 3009 162995 3043
rect 206017 3009 206051 3043
rect 207765 3009 207799 3043
rect 208685 3009 208719 3043
rect 210985 3009 211019 3043
rect 211102 3009 211136 3043
rect 212641 3009 212675 3043
rect 213561 3009 213595 3043
rect 213699 3009 213733 3043
rect 215585 3009 215619 3043
rect 216321 3009 216355 3043
rect 216597 3009 216631 3043
rect 217977 3009 218011 3043
rect 221565 3009 221599 3043
rect 222209 3009 222243 3043
rect 222945 3009 222979 3043
rect 223221 3009 223255 3043
rect 224049 3009 224083 3043
rect 227085 3009 227119 3043
rect 228097 3009 228131 3043
rect 257629 3009 257663 3043
rect 259009 3009 259043 3043
rect 266185 3009 266219 3043
rect 266829 3009 266863 3043
rect 267473 3009 267507 3043
rect 268117 3009 268151 3043
rect 268761 3009 268795 3043
rect 269865 3009 269899 3043
rect 270969 3009 271003 3043
rect 24961 2941 24995 2975
rect 25237 2941 25271 2975
rect 26065 2941 26099 2975
rect 27353 2941 27387 2975
rect 82093 2941 82127 2975
rect 84301 2941 84335 2975
rect 84485 2941 84519 2975
rect 86785 2941 86819 2975
rect 88441 2941 88475 2975
rect 90097 2941 90131 2975
rect 90281 2941 90315 2975
rect 94421 2941 94455 2975
rect 97825 2941 97859 2975
rect 97963 2941 97997 2975
rect 99849 2941 99883 2975
rect 100585 2941 100619 2975
rect 100702 2941 100736 2975
rect 100861 2941 100895 2975
rect 101873 2941 101907 2975
rect 102333 2941 102367 2975
rect 102747 2941 102781 2975
rect 103529 2941 103563 2975
rect 104449 2941 104483 2975
rect 104633 2941 104667 2975
rect 106289 2941 106323 2975
rect 107301 2941 107335 2975
rect 107669 2941 107703 2975
rect 116685 2941 116719 2975
rect 116961 2941 116995 2975
rect 121561 2941 121595 2975
rect 137937 2941 137971 2975
rect 138790 2941 138824 2975
rect 138949 2941 138983 2975
rect 140513 2941 140547 2975
rect 140973 2941 141007 2975
rect 142813 2941 142847 2975
rect 143457 2941 143491 2975
rect 143871 2941 143905 2975
rect 144009 2941 144043 2975
rect 145665 2941 145699 2975
rect 146723 2941 146757 2975
rect 148149 2941 148183 2975
rect 148609 2941 148643 2975
rect 149002 2941 149036 2975
rect 149805 2941 149839 2975
rect 150817 2941 150851 2975
rect 151001 2941 151035 2975
rect 151277 2941 151311 2975
rect 156153 2941 156187 2975
rect 157165 2941 157199 2975
rect 157901 2941 157935 2975
rect 158085 2941 158119 2975
rect 159097 2941 159131 2975
rect 161581 2941 161615 2975
rect 167745 2941 167779 2975
rect 202337 2941 202371 2975
rect 204177 2941 204211 2975
rect 204361 2941 204395 2975
rect 207949 2941 207983 2975
rect 208409 2941 208443 2975
rect 208823 2941 208857 2975
rect 208961 2941 208995 2975
rect 210065 2941 210099 2975
rect 210249 2941 210283 2975
rect 211261 2941 211295 2975
rect 212825 2941 212859 2975
rect 213837 2941 213871 2975
rect 215401 2941 215435 2975
rect 216045 2941 216079 2975
rect 216459 2941 216493 2975
rect 217793 2941 217827 2975
rect 218897 2941 218931 2975
rect 219081 2941 219115 2975
rect 221749 2941 221783 2975
rect 226625 2941 226659 2975
rect 235825 2941 235859 2975
rect 24501 2873 24535 2907
rect 28181 2873 28215 2907
rect 39129 2873 39163 2907
rect 41153 2873 41187 2907
rect 88993 2873 89027 2907
rect 97549 2873 97583 2907
rect 100309 2873 100343 2907
rect 115765 2873 115799 2907
rect 116133 2873 116167 2907
rect 138397 2873 138431 2907
rect 146309 2873 146343 2907
rect 156613 2873 156647 2907
rect 158545 2873 158579 2907
rect 203809 2873 203843 2907
rect 210709 2873 210743 2907
rect 213285 2873 213319 2907
rect 260113 2873 260147 2907
rect 267289 2873 267323 2907
rect 267933 2873 267967 2907
rect 270785 2873 270819 2907
rect 25605 2805 25639 2839
rect 26433 2805 26467 2839
rect 27261 2805 27295 2839
rect 27721 2805 27755 2839
rect 89361 2805 89395 2839
rect 89729 2805 89763 2839
rect 103897 2805 103931 2839
rect 106565 2805 106599 2839
rect 118709 2805 118743 2839
rect 139869 2805 139903 2839
rect 142629 2805 142663 2839
rect 163145 2805 163179 2839
rect 209605 2805 209639 2839
rect 218161 2805 218195 2839
rect 219449 2805 219483 2839
rect 227269 2805 227303 2839
rect 228281 2805 228315 2839
rect 257813 2805 257847 2839
rect 259193 2805 259227 2839
rect 265541 2805 265575 2839
rect 266645 2805 266679 2839
rect 270049 2805 270083 2839
rect 23949 2601 23983 2635
rect 25237 2601 25271 2635
rect 26249 2601 26283 2635
rect 27077 2601 27111 2635
rect 28089 2601 28123 2635
rect 58633 2601 58667 2635
rect 60841 2601 60875 2635
rect 85773 2601 85807 2635
rect 98561 2601 98595 2635
rect 105277 2601 105311 2635
rect 157901 2601 157935 2635
rect 160569 2601 160603 2635
rect 161305 2601 161339 2635
rect 190561 2601 190595 2635
rect 192033 2601 192067 2635
rect 202981 2601 203015 2635
rect 211905 2601 211939 2635
rect 224141 2601 224175 2635
rect 224509 2601 224543 2635
rect 225889 2601 225923 2635
rect 227177 2601 227211 2635
rect 236009 2601 236043 2635
rect 267105 2601 267139 2635
rect 97365 2533 97399 2567
rect 104081 2533 104115 2567
rect 143733 2533 143767 2567
rect 144929 2533 144963 2567
rect 148885 2533 148919 2567
rect 155049 2533 155083 2567
rect 210709 2533 210743 2567
rect 243691 2533 243725 2567
rect 1869 2465 1903 2499
rect 53757 2465 53791 2499
rect 78229 2465 78263 2499
rect 88073 2465 88107 2499
rect 90189 2465 90223 2499
rect 90557 2465 90591 2499
rect 96721 2465 96755 2499
rect 97758 2465 97792 2499
rect 99389 2465 99423 2499
rect 99573 2465 99607 2499
rect 103437 2465 103471 2499
rect 104357 2465 104391 2499
rect 104495 2465 104529 2499
rect 108497 2465 108531 2499
rect 109049 2465 109083 2499
rect 139133 2465 139167 2499
rect 143089 2465 143123 2499
rect 144009 2465 144043 2499
rect 148241 2465 148275 2499
rect 149161 2465 149195 2499
rect 149299 2465 149333 2499
rect 150725 2465 150759 2499
rect 152381 2465 152415 2499
rect 179889 2465 179923 2499
rect 187249 2465 187283 2499
rect 201969 2465 202003 2499
rect 204913 2465 204947 2499
rect 205097 2465 205131 2499
rect 205373 2465 205407 2499
rect 210065 2465 210099 2499
rect 210985 2465 211019 2499
rect 216229 2465 216263 2499
rect 218621 2465 218655 2499
rect 219541 2465 219575 2499
rect 221013 2465 221047 2499
rect 221933 2465 221967 2499
rect 222117 2465 222151 2499
rect 223221 2465 223255 2499
rect 246681 2465 246715 2499
rect 258917 2465 258951 2499
rect 1593 2397 1627 2431
rect 23765 2397 23799 2431
rect 24961 2397 24995 2431
rect 25053 2397 25087 2431
rect 25605 2397 25639 2431
rect 25881 2397 25915 2431
rect 26065 2397 26099 2431
rect 26801 2397 26835 2431
rect 26893 2397 26927 2431
rect 27445 2397 27479 2431
rect 27813 2397 27847 2431
rect 27905 2397 27939 2431
rect 28549 2397 28583 2431
rect 32229 2397 32263 2431
rect 32413 2397 32447 2431
rect 53941 2397 53975 2431
rect 54677 2397 54711 2431
rect 55505 2397 55539 2431
rect 57621 2397 57655 2431
rect 59185 2397 59219 2431
rect 60657 2397 60691 2431
rect 62773 2397 62807 2431
rect 65809 2397 65843 2431
rect 71329 2397 71363 2431
rect 71605 2397 71639 2431
rect 73537 2397 73571 2431
rect 73813 2397 73847 2431
rect 76481 2397 76515 2431
rect 76757 2397 76791 2431
rect 77953 2397 77987 2431
rect 79425 2397 79459 2431
rect 79701 2397 79735 2431
rect 82093 2397 82127 2431
rect 82369 2397 82403 2431
rect 83565 2397 83599 2431
rect 87429 2397 87463 2431
rect 88349 2397 88383 2431
rect 90649 2397 90683 2431
rect 91569 2397 91603 2431
rect 92857 2397 92891 2431
rect 93685 2397 93719 2431
rect 94421 2397 94455 2431
rect 95157 2397 95191 2431
rect 95893 2397 95927 2431
rect 96905 2397 96939 2431
rect 97641 2397 97675 2431
rect 97917 2397 97951 2431
rect 103621 2397 103655 2431
rect 104633 2397 104667 2431
rect 122481 2397 122515 2431
rect 124597 2397 124631 2431
rect 126161 2397 126195 2431
rect 127633 2397 127667 2431
rect 128369 2397 128403 2431
rect 129841 2397 129875 2431
rect 131405 2397 131439 2431
rect 132785 2397 132819 2431
rect 133521 2397 133555 2431
rect 134257 2397 134291 2431
rect 138949 2397 138983 2431
rect 143273 2397 143307 2431
rect 144147 2397 144181 2431
rect 144285 2397 144319 2431
rect 148425 2397 148459 2431
rect 149437 2397 149471 2431
rect 150081 2397 150115 2431
rect 150541 2397 150575 2431
rect 155233 2397 155267 2431
rect 156567 2397 156601 2431
rect 157349 2397 157383 2431
rect 157717 2397 157751 2431
rect 158637 2397 158671 2431
rect 159925 2397 159959 2431
rect 160109 2397 160143 2431
rect 160385 2397 160419 2431
rect 160753 2397 160787 2431
rect 161581 2397 161615 2431
rect 163697 2397 163731 2431
rect 164433 2397 164467 2431
rect 165169 2397 165203 2431
rect 165905 2397 165939 2431
rect 166641 2397 166675 2431
rect 167745 2397 167779 2431
rect 167837 2397 167871 2431
rect 176669 2397 176703 2431
rect 176945 2397 176979 2431
rect 179613 2397 179647 2431
rect 186973 2397 187007 2431
rect 190377 2397 190411 2431
rect 191113 2397 191147 2431
rect 191849 2397 191883 2431
rect 194885 2397 194919 2431
rect 196265 2397 196299 2431
rect 197185 2397 197219 2431
rect 197277 2397 197311 2431
rect 198381 2397 198415 2431
rect 199761 2397 199795 2431
rect 201233 2397 201267 2431
rect 202153 2397 202187 2431
rect 202337 2397 202371 2431
rect 202797 2397 202831 2431
rect 210249 2397 210283 2431
rect 211102 2397 211136 2431
rect 211261 2397 211295 2431
rect 216045 2397 216079 2431
rect 217333 2397 217367 2431
rect 217517 2397 217551 2431
rect 218805 2397 218839 2431
rect 220829 2397 220863 2431
rect 222853 2397 222887 2431
rect 223037 2397 223071 2431
rect 225337 2397 225371 2431
rect 225705 2397 225739 2431
rect 226257 2397 226291 2431
rect 226993 2397 227027 2431
rect 227913 2397 227947 2431
rect 228189 2397 228223 2431
rect 228833 2397 228867 2431
rect 231133 2397 231167 2431
rect 231869 2397 231903 2431
rect 232605 2397 232639 2431
rect 235825 2397 235859 2431
rect 236561 2397 236595 2431
rect 243461 2397 243495 2431
rect 246405 2397 246439 2431
rect 256709 2397 256743 2431
rect 256985 2397 257019 2431
rect 259101 2397 259135 2431
rect 259285 2397 259319 2431
rect 259745 2397 259779 2431
rect 261585 2397 261619 2431
rect 263977 2397 264011 2431
rect 264161 2397 264195 2431
rect 264345 2397 264379 2431
rect 264805 2397 264839 2431
rect 267289 2397 267323 2431
rect 267933 2397 267967 2431
rect 268577 2397 268611 2431
rect 269129 2397 269163 2431
rect 269221 2397 269255 2431
rect 269865 2397 269899 2431
rect 270601 2397 270635 2431
rect 24777 2329 24811 2363
rect 37197 2329 37231 2363
rect 37289 2329 37323 2363
rect 37657 2329 37691 2363
rect 83749 2329 83783 2363
rect 85405 2329 85439 2363
rect 88533 2329 88567 2363
rect 101229 2329 101263 2363
rect 108681 2329 108715 2363
rect 140789 2329 140823 2363
rect 156981 2329 157015 2363
rect 159097 2329 159131 2363
rect 160293 2329 160327 2363
rect 216965 2329 216999 2363
rect 218253 2329 218287 2363
rect 219265 2329 219299 2363
rect 258089 2329 258123 2363
rect 28733 2261 28767 2295
rect 32597 2261 32631 2295
rect 33057 2261 33091 2295
rect 36921 2261 36955 2295
rect 38025 2261 38059 2295
rect 38209 2261 38243 2295
rect 54125 2261 54159 2295
rect 54861 2261 54895 2295
rect 55689 2261 55723 2295
rect 57805 2261 57839 2295
rect 59369 2261 59403 2295
rect 62957 2261 62991 2295
rect 65993 2261 66027 2295
rect 66637 2261 66671 2295
rect 83289 2261 83323 2295
rect 87613 2261 87647 2295
rect 90833 2261 90867 2295
rect 91753 2261 91787 2295
rect 93041 2261 93075 2295
rect 93869 2261 93903 2295
rect 94605 2261 94639 2295
rect 95341 2261 95375 2295
rect 96077 2261 96111 2295
rect 99021 2261 99055 2295
rect 122665 2261 122699 2295
rect 124781 2261 124815 2295
rect 126345 2261 126379 2295
rect 127817 2261 127851 2295
rect 128553 2261 128587 2295
rect 130025 2261 130059 2295
rect 131589 2261 131623 2295
rect 132969 2261 133003 2295
rect 133705 2261 133739 2295
rect 134441 2261 134475 2295
rect 134993 2261 135027 2295
rect 138673 2261 138707 2295
rect 141157 2261 141191 2295
rect 157533 2261 157567 2295
rect 160937 2261 160971 2295
rect 161765 2261 161799 2295
rect 163881 2261 163915 2295
rect 164617 2261 164651 2295
rect 165353 2261 165387 2295
rect 166089 2261 166123 2295
rect 166825 2261 166859 2295
rect 168021 2261 168055 2295
rect 191297 2261 191331 2295
rect 195069 2261 195103 2295
rect 196449 2261 196483 2295
rect 197461 2261 197495 2295
rect 198565 2261 198599 2295
rect 199945 2261 199979 2295
rect 201417 2261 201451 2295
rect 204269 2261 204303 2295
rect 207029 2261 207063 2295
rect 216689 2261 216723 2295
rect 217977 2261 218011 2295
rect 220461 2261 220495 2295
rect 221473 2261 221507 2295
rect 222577 2261 222611 2295
rect 223681 2261 223715 2295
rect 224969 2261 225003 2295
rect 225521 2261 225555 2295
rect 226441 2261 226475 2295
rect 229017 2261 229051 2295
rect 231317 2261 231351 2295
rect 232053 2261 232087 2295
rect 232789 2261 232823 2295
rect 236745 2261 236779 2295
rect 258181 2261 258215 2295
rect 259929 2261 259963 2295
rect 261769 2261 261803 2295
rect 264989 2261 265023 2295
rect 266001 2261 266035 2295
rect 267749 2261 267783 2295
rect 268393 2261 268427 2295
rect 269405 2261 269439 2295
rect 270049 2261 270083 2295
rect 270785 2261 270819 2295
rect 6929 2057 6963 2091
rect 23857 2057 23891 2091
rect 26341 2057 26375 2091
rect 57529 2057 57563 2091
rect 58541 2057 58575 2091
rect 59277 2057 59311 2091
rect 62681 2057 62715 2091
rect 65257 2057 65291 2091
rect 91109 2057 91143 2091
rect 92765 2057 92799 2091
rect 94513 2057 94547 2091
rect 95433 2057 95467 2091
rect 96261 2057 96295 2091
rect 102057 2057 102091 2091
rect 112085 2057 112119 2091
rect 117237 2057 117271 2091
rect 122021 2057 122055 2091
rect 124505 2057 124539 2091
rect 126253 2057 126287 2091
rect 127909 2057 127943 2091
rect 129657 2057 129691 2091
rect 131681 2057 131715 2091
rect 149897 2057 149931 2091
rect 155325 2057 155359 2091
rect 162317 2057 162351 2091
rect 163973 2057 164007 2091
rect 165629 2057 165663 2091
rect 166641 2057 166675 2091
rect 167469 2057 167503 2091
rect 191113 2057 191147 2091
rect 192401 2057 192435 2091
rect 195713 2057 195747 2091
rect 197553 2057 197587 2091
rect 199209 2057 199243 2091
rect 200865 2057 200899 2091
rect 211537 2057 211571 2091
rect 216137 2057 216171 2091
rect 217149 2057 217183 2091
rect 221657 2057 221691 2091
rect 225337 2057 225371 2091
rect 226165 2057 226199 2091
rect 226993 2057 227027 2091
rect 228465 2057 228499 2091
rect 236101 2057 236135 2091
rect 245071 2057 245105 2091
rect 251465 2057 251499 2091
rect 257997 2057 258031 2091
rect 259377 2057 259411 2091
rect 261861 2057 261895 2091
rect 269681 2057 269715 2091
rect 270509 2057 270543 2091
rect 9229 1989 9263 2023
rect 17141 1989 17175 2023
rect 25237 1989 25271 2023
rect 26249 1989 26283 2023
rect 27261 1989 27295 2023
rect 35541 1989 35575 2023
rect 35817 1989 35851 2023
rect 36277 1989 36311 2023
rect 36645 1989 36679 2023
rect 39037 1989 39071 2023
rect 39313 1989 39347 2023
rect 39773 1989 39807 2023
rect 40141 1989 40175 2023
rect 54217 1989 54251 2023
rect 55045 1989 55079 2023
rect 99481 1989 99515 2023
rect 133613 1989 133647 2023
rect 139961 1989 139995 2023
rect 216689 1989 216723 2023
rect 218437 1989 218471 2023
rect 231777 1989 231811 2023
rect 232605 1989 232639 2023
rect 2605 1921 2639 1955
rect 4813 1921 4847 1955
rect 6837 1921 6871 1955
rect 7573 1921 7607 1955
rect 9045 1921 9079 1955
rect 14381 1921 14415 1955
rect 15669 1921 15703 1955
rect 15853 1921 15887 1955
rect 16957 1921 16991 1955
rect 23581 1921 23615 1955
rect 23673 1921 23707 1955
rect 24317 1921 24351 1955
rect 24501 1921 24535 1955
rect 28641 1921 28675 1955
rect 28825 1921 28859 1955
rect 29561 1921 29595 1955
rect 29653 1921 29687 1955
rect 30389 1921 30423 1955
rect 30573 1921 30607 1955
rect 31401 1921 31435 1955
rect 31585 1921 31619 1955
rect 32413 1921 32447 1955
rect 32505 1921 32539 1955
rect 32689 1921 32723 1955
rect 33149 1921 33183 1955
rect 35909 1921 35943 1955
rect 38117 1921 38151 1955
rect 39405 1921 39439 1955
rect 45477 1921 45511 1955
rect 50629 1921 50663 1955
rect 52929 1921 52963 1955
rect 54033 1921 54067 1955
rect 54861 1921 54895 1955
rect 55505 1921 55539 1955
rect 55689 1921 55723 1955
rect 56333 1921 56367 1955
rect 56517 1921 56551 1955
rect 57161 1921 57195 1955
rect 57345 1921 57379 1955
rect 58081 1921 58115 1955
rect 59093 1921 59127 1955
rect 59829 1921 59863 1955
rect 60013 1921 60047 1955
rect 60657 1921 60691 1955
rect 60841 1921 60875 1955
rect 61577 1921 61611 1955
rect 61669 1921 61703 1955
rect 62405 1921 62439 1955
rect 62497 1921 62531 1955
rect 63233 1921 63267 1955
rect 63417 1921 63451 1955
rect 64061 1921 64095 1955
rect 64245 1921 64279 1955
rect 65073 1921 65107 1955
rect 65717 1921 65751 1955
rect 65901 1921 65935 1955
rect 66637 1921 66671 1955
rect 66729 1921 66763 1955
rect 66913 1921 66947 1955
rect 67373 1921 67407 1955
rect 70869 1921 70903 1955
rect 72341 1921 72375 1955
rect 76021 1921 76055 1955
rect 77493 1921 77527 1955
rect 80161 1921 80195 1955
rect 82461 1921 82495 1955
rect 86417 1921 86451 1955
rect 87797 1921 87831 1955
rect 88073 1921 88107 1955
rect 88257 1921 88291 1955
rect 88441 1921 88475 1955
rect 89269 1921 89303 1955
rect 89453 1921 89487 1955
rect 90005 1921 90039 1955
rect 90097 1921 90131 1955
rect 90741 1921 90775 1955
rect 90925 1921 90959 1955
rect 91753 1921 91787 1955
rect 92397 1921 92431 1955
rect 92581 1921 92615 1955
rect 93317 1921 93351 1955
rect 93409 1921 93443 1955
rect 94145 1921 94179 1955
rect 94329 1921 94363 1955
rect 95157 1921 95191 1955
rect 95249 1921 95283 1955
rect 96077 1921 96111 1955
rect 96905 1921 96939 1955
rect 97733 1921 97767 1955
rect 98561 1921 98595 1955
rect 100493 1921 100527 1955
rect 100677 1921 100711 1955
rect 101137 1921 101171 1955
rect 101873 1921 101907 1955
rect 107117 1921 107151 1955
rect 112269 1921 112303 1955
rect 117421 1921 117455 1955
rect 120917 1921 120951 1955
rect 121009 1921 121043 1955
rect 121837 1921 121871 1955
rect 122665 1921 122699 1955
rect 123493 1921 123527 1955
rect 124137 1921 124171 1955
rect 124321 1921 124355 1955
rect 125057 1921 125091 1955
rect 125241 1921 125275 1955
rect 125977 1921 126011 1955
rect 126069 1921 126103 1955
rect 126713 1921 126747 1955
rect 126897 1921 126931 1955
rect 127633 1921 127667 1955
rect 127725 1921 127759 1955
rect 128553 1921 128587 1955
rect 128645 1921 128679 1955
rect 129381 1921 129415 1955
rect 129473 1921 129507 1955
rect 130577 1921 130611 1955
rect 130669 1921 130703 1955
rect 131313 1921 131347 1955
rect 131497 1921 131531 1955
rect 132233 1921 132267 1955
rect 132417 1921 132451 1955
rect 133245 1921 133279 1955
rect 133429 1921 133463 1955
rect 134165 1921 134199 1955
rect 134257 1921 134291 1955
rect 134441 1921 134475 1955
rect 135361 1921 135395 1955
rect 138121 1921 138155 1955
rect 139041 1921 139075 1955
rect 139179 1921 139213 1955
rect 140513 1921 140547 1955
rect 141433 1921 141467 1955
rect 141709 1921 141743 1955
rect 142997 1921 143031 1955
rect 144929 1921 144963 1955
rect 150081 1921 150115 1955
rect 155141 1921 155175 1955
rect 155969 1921 156003 1955
rect 156797 1921 156831 1955
rect 157993 1921 158027 1955
rect 159281 1921 159315 1955
rect 159925 1921 159959 1955
rect 160109 1921 160143 1955
rect 161213 1921 161247 1955
rect 161305 1921 161339 1955
rect 161949 1921 161983 1955
rect 162133 1921 162167 1955
rect 162777 1921 162811 1955
rect 162961 1921 162995 1955
rect 163697 1921 163731 1955
rect 163789 1921 163823 1955
rect 164433 1921 164467 1955
rect 164617 1921 164651 1955
rect 165261 1921 165295 1955
rect 165445 1921 165479 1955
rect 166273 1921 166307 1955
rect 166457 1921 166491 1955
rect 167101 1921 167135 1955
rect 167285 1921 167319 1955
rect 167929 1921 167963 1955
rect 168113 1921 168147 1955
rect 168297 1921 168331 1955
rect 168757 1921 168791 1955
rect 173265 1921 173299 1955
rect 174737 1921 174771 1955
rect 176853 1921 176887 1955
rect 179429 1921 179463 1955
rect 181913 1921 181947 1955
rect 183569 1921 183603 1955
rect 185041 1921 185075 1955
rect 187157 1921 187191 1955
rect 189733 1921 189767 1955
rect 190837 1921 190871 1955
rect 190929 1921 190963 1955
rect 192125 1921 192159 1955
rect 192217 1921 192251 1955
rect 192953 1921 192987 1955
rect 193045 1921 193079 1955
rect 193689 1921 193723 1955
rect 193873 1921 193907 1955
rect 194609 1921 194643 1955
rect 194701 1921 194735 1955
rect 195437 1921 195471 1955
rect 195529 1921 195563 1955
rect 196173 1921 196207 1955
rect 196357 1921 196391 1955
rect 197185 1921 197219 1955
rect 197369 1921 197403 1955
rect 198013 1921 198047 1955
rect 198197 1921 198231 1955
rect 198841 1921 198875 1955
rect 199025 1921 199059 1955
rect 199669 1921 199703 1955
rect 199853 1921 199887 1955
rect 200497 1921 200531 1955
rect 200681 1921 200715 1955
rect 201325 1921 201359 1955
rect 201509 1921 201543 1955
rect 202337 1921 202371 1955
rect 202521 1921 202555 1955
rect 202705 1921 202739 1955
rect 203165 1921 203199 1955
rect 211721 1921 211755 1955
rect 216321 1921 216355 1955
rect 216413 1921 216447 1955
rect 217793 1921 217827 1955
rect 218713 1921 218747 1955
rect 218897 1921 218931 1955
rect 219817 1921 219851 1955
rect 220093 1921 220127 1955
rect 220737 1921 220771 1955
rect 221841 1921 221875 1955
rect 222945 1921 222979 1955
rect 223221 1921 223255 1955
rect 223865 1921 223899 1955
rect 224969 1921 225003 1955
rect 225153 1921 225187 1955
rect 225889 1921 225923 1955
rect 225981 1921 226015 1955
rect 226717 1921 226751 1955
rect 226812 1921 226846 1955
rect 228097 1921 228131 1955
rect 228281 1921 228315 1955
rect 228925 1921 228959 1955
rect 229109 1921 229143 1955
rect 229753 1921 229787 1955
rect 229957 1921 229991 1955
rect 230581 1921 230615 1955
rect 230765 1921 230799 1955
rect 231501 1921 231535 1955
rect 231593 1921 231627 1955
rect 232237 1921 232271 1955
rect 232421 1921 232455 1955
rect 233341 1921 233375 1955
rect 233433 1921 233467 1955
rect 234261 1921 234295 1955
rect 234905 1921 234939 1955
rect 235089 1921 235123 1955
rect 235917 1921 235951 1955
rect 236745 1921 236779 1955
rect 236929 1921 236963 1955
rect 237389 1921 237423 1955
rect 241529 1921 241563 1955
rect 250269 1921 250303 1955
rect 251373 1921 251407 1955
rect 252569 1921 252603 1955
rect 255421 1921 255455 1955
rect 256709 1921 256743 1955
rect 257905 1921 257939 1955
rect 259009 1921 259043 1955
rect 259193 1921 259227 1955
rect 259929 1921 259963 1955
rect 260021 1921 260055 1955
rect 260665 1921 260699 1955
rect 260849 1921 260883 1955
rect 261493 1921 261527 1955
rect 261677 1921 261711 1955
rect 262321 1921 262355 1955
rect 262505 1921 262539 1955
rect 263149 1921 263183 1955
rect 263333 1921 263367 1955
rect 264345 1921 264379 1955
rect 265173 1921 265207 1955
rect 266001 1921 266035 1955
rect 266829 1921 266863 1955
rect 267657 1921 267691 1955
rect 268485 1921 268519 1955
rect 269497 1921 269531 1955
rect 270233 1921 270267 1955
rect 270325 1921 270359 1955
rect 2329 1853 2363 1887
rect 4537 1853 4571 1887
rect 14105 1853 14139 1887
rect 53849 1853 53883 1887
rect 54677 1853 54711 1887
rect 57897 1853 57931 1887
rect 58909 1853 58943 1887
rect 64889 1853 64923 1887
rect 70593 1853 70627 1887
rect 72065 1853 72099 1887
rect 74273 1853 74307 1887
rect 74549 1853 74583 1887
rect 75745 1853 75779 1887
rect 77217 1853 77251 1887
rect 79885 1853 79919 1887
rect 81173 1853 81207 1887
rect 81449 1853 81483 1887
rect 82737 1853 82771 1887
rect 83841 1853 83875 1887
rect 84025 1853 84059 1887
rect 85681 1853 85715 1887
rect 86141 1853 86175 1887
rect 89085 1853 89119 1887
rect 91569 1853 91603 1887
rect 95893 1853 95927 1887
rect 96721 1853 96755 1887
rect 97549 1853 97583 1887
rect 98377 1853 98411 1887
rect 99757 1853 99791 1887
rect 100309 1853 100343 1887
rect 121653 1853 121687 1887
rect 122481 1853 122515 1887
rect 123309 1853 123343 1887
rect 138305 1853 138339 1887
rect 138765 1853 138799 1887
rect 139317 1853 139351 1887
rect 140697 1853 140731 1887
rect 141550 1853 141584 1887
rect 157073 1853 157107 1887
rect 158269 1853 158303 1887
rect 159097 1853 159131 1887
rect 172989 1853 173023 1887
rect 174461 1853 174495 1887
rect 176577 1853 176611 1887
rect 177865 1853 177899 1887
rect 178141 1853 178175 1887
rect 179153 1853 179187 1887
rect 183293 1853 183327 1887
rect 184765 1853 184799 1887
rect 186881 1853 186915 1887
rect 188169 1853 188203 1887
rect 188445 1853 188479 1887
rect 189457 1853 189491 1887
rect 217977 1853 218011 1887
rect 219173 1853 219207 1887
rect 221013 1853 221047 1887
rect 224141 1853 224175 1887
rect 234077 1853 234111 1887
rect 235733 1853 235767 1887
rect 236561 1853 236595 1887
rect 241253 1853 241287 1887
rect 243553 1853 243587 1887
rect 243829 1853 243863 1887
rect 244841 1853 244875 1887
rect 246129 1853 246163 1887
rect 246405 1853 246439 1887
rect 248705 1853 248739 1887
rect 248981 1853 249015 1887
rect 249993 1853 250027 1887
rect 252293 1853 252327 1887
rect 253857 1853 253891 1887
rect 254133 1853 254167 1887
rect 255145 1853 255179 1887
rect 256433 1853 256467 1887
rect 264161 1853 264195 1887
rect 264989 1853 265023 1887
rect 265817 1853 265851 1887
rect 266645 1853 266679 1887
rect 267473 1853 267507 1887
rect 268301 1853 268335 1887
rect 269313 1853 269347 1887
rect 7757 1785 7791 1819
rect 25421 1785 25455 1819
rect 37933 1785 37967 1819
rect 40325 1785 40359 1819
rect 45293 1785 45327 1819
rect 50445 1785 50479 1819
rect 53113 1785 53147 1819
rect 98745 1785 98779 1819
rect 106933 1785 106967 1819
rect 141157 1785 141191 1819
rect 142813 1785 142847 1819
rect 144745 1785 144779 1819
rect 24685 1717 24719 1751
rect 27353 1717 27387 1751
rect 29009 1717 29043 1751
rect 29837 1717 29871 1751
rect 30757 1717 30791 1751
rect 31769 1717 31803 1751
rect 33333 1717 33367 1751
rect 36829 1717 36863 1751
rect 53481 1717 53515 1751
rect 55873 1717 55907 1751
rect 56701 1717 56735 1751
rect 58265 1717 58299 1751
rect 60197 1717 60231 1751
rect 61025 1717 61059 1751
rect 61853 1717 61887 1751
rect 63601 1717 63635 1751
rect 64429 1717 64463 1751
rect 66085 1717 66119 1751
rect 67557 1717 67591 1751
rect 86049 1717 86083 1751
rect 90281 1717 90315 1751
rect 91937 1717 91971 1751
rect 93593 1717 93627 1751
rect 97089 1717 97123 1751
rect 97917 1717 97951 1751
rect 101321 1717 101355 1751
rect 121193 1717 121227 1751
rect 122849 1717 122883 1751
rect 123677 1717 123711 1751
rect 125425 1717 125459 1751
rect 127081 1717 127115 1751
rect 128829 1717 128863 1751
rect 130853 1717 130887 1751
rect 132601 1717 132635 1751
rect 135545 1717 135579 1751
rect 142353 1717 142387 1751
rect 156153 1717 156187 1751
rect 159465 1717 159499 1751
rect 160293 1717 160327 1751
rect 161489 1717 161523 1751
rect 163145 1717 163179 1751
rect 164801 1717 164835 1751
rect 168941 1717 168975 1751
rect 182005 1717 182039 1751
rect 193229 1717 193263 1751
rect 194057 1717 194091 1751
rect 194885 1717 194919 1751
rect 196541 1717 196575 1751
rect 198381 1717 198415 1751
rect 200037 1717 200071 1751
rect 201693 1717 201727 1751
rect 203349 1717 203383 1751
rect 229293 1717 229327 1751
rect 230121 1717 230155 1751
rect 230949 1717 230983 1751
rect 233617 1717 233651 1751
rect 234445 1717 234479 1751
rect 235273 1717 235307 1751
rect 237573 1717 237607 1751
rect 260205 1717 260239 1751
rect 261033 1717 261067 1751
rect 262689 1717 262723 1751
rect 263517 1717 263551 1751
rect 264529 1717 264563 1751
rect 265357 1717 265391 1751
rect 266185 1717 266219 1751
rect 267013 1717 267047 1751
rect 267841 1717 267875 1751
rect 268669 1717 268703 1751
rect 25973 1513 26007 1547
rect 28365 1513 28399 1547
rect 35449 1513 35483 1547
rect 60013 1513 60047 1547
rect 95157 1513 95191 1547
rect 113373 1513 113407 1547
rect 156797 1513 156831 1547
rect 157625 1513 157659 1547
rect 180625 1513 180659 1547
rect 221657 1513 221691 1547
rect 225889 1513 225923 1547
rect 228465 1513 228499 1547
rect 232513 1513 232547 1547
rect 236193 1513 236227 1547
rect 36737 1445 36771 1479
rect 38669 1445 38703 1479
rect 44465 1445 44499 1479
rect 133337 1445 133371 1479
rect 134349 1445 134383 1479
rect 138121 1445 138155 1479
rect 139225 1445 139259 1479
rect 140513 1445 140547 1479
rect 191389 1445 191423 1479
rect 213285 1445 213319 1479
rect 1777 1377 1811 1411
rect 24961 1377 24995 1411
rect 27169 1377 27203 1411
rect 27997 1377 28031 1411
rect 34345 1377 34379 1411
rect 53941 1377 53975 1411
rect 69121 1377 69155 1411
rect 88073 1377 88107 1411
rect 98377 1377 98411 1411
rect 99941 1377 99975 1411
rect 103253 1377 103287 1411
rect 157257 1377 157291 1411
rect 158545 1377 158579 1411
rect 159373 1377 159407 1411
rect 163697 1377 163731 1411
rect 167009 1377 167043 1411
rect 171701 1377 171735 1411
rect 201233 1377 201267 1411
rect 202337 1377 202371 1411
rect 205833 1377 205867 1411
rect 225521 1377 225555 1411
rect 226533 1377 226567 1411
rect 228097 1377 228131 1411
rect 232145 1377 232179 1411
rect 235825 1377 235859 1411
rect 239965 1377 239999 1411
rect 257721 1377 257755 1411
rect 269313 1377 269347 1411
rect 2605 1309 2639 1343
rect 2881 1309 2915 1343
rect 5181 1309 5215 1343
rect 5457 1309 5491 1343
rect 6561 1309 6595 1343
rect 6837 1309 6871 1343
rect 9505 1309 9539 1343
rect 11161 1309 11195 1343
rect 12173 1309 12207 1343
rect 14841 1309 14875 1343
rect 15117 1309 15151 1343
rect 23765 1309 23799 1343
rect 24685 1309 24719 1343
rect 25145 1309 25179 1343
rect 27353 1309 27387 1343
rect 27537 1309 27571 1343
rect 28181 1309 28215 1343
rect 28917 1309 28951 1343
rect 29745 1309 29779 1343
rect 30573 1309 30607 1343
rect 31401 1309 31435 1343
rect 32321 1309 32355 1343
rect 35633 1309 35667 1343
rect 36277 1309 36311 1343
rect 36921 1309 36955 1343
rect 38209 1309 38243 1343
rect 38853 1309 38887 1343
rect 39497 1309 39531 1343
rect 40785 1309 40819 1343
rect 41429 1309 41463 1343
rect 42073 1309 42107 1343
rect 43269 1309 43303 1343
rect 44005 1309 44039 1343
rect 44649 1309 44683 1343
rect 45937 1309 45971 1343
rect 46581 1309 46615 1343
rect 47225 1309 47259 1343
rect 48421 1309 48455 1343
rect 49157 1309 49191 1343
rect 49801 1309 49835 1343
rect 51089 1309 51123 1343
rect 51733 1309 51767 1343
rect 52377 1309 52411 1343
rect 53205 1309 53239 1343
rect 54125 1309 54159 1343
rect 56057 1309 56091 1343
rect 56885 1309 56919 1343
rect 58449 1309 58483 1343
rect 59369 1309 59403 1343
rect 59737 1309 59771 1343
rect 59829 1309 59863 1343
rect 60657 1309 60691 1343
rect 61393 1309 61427 1343
rect 62129 1309 62163 1343
rect 63601 1309 63635 1343
rect 64337 1309 64371 1343
rect 65993 1309 66027 1343
rect 69581 1309 69615 1343
rect 69857 1309 69891 1343
rect 72157 1309 72191 1343
rect 72433 1309 72467 1343
rect 74733 1309 74767 1343
rect 75009 1309 75043 1343
rect 77309 1309 77343 1343
rect 77585 1309 77619 1343
rect 79885 1309 79919 1343
rect 80161 1309 80195 1343
rect 82461 1309 82495 1343
rect 82737 1309 82771 1343
rect 85037 1309 85071 1343
rect 85313 1309 85347 1343
rect 86785 1309 86819 1343
rect 87061 1309 87095 1343
rect 88257 1309 88291 1343
rect 88441 1309 88475 1343
rect 89085 1309 89119 1343
rect 89177 1309 89211 1343
rect 89361 1309 89395 1343
rect 90465 1309 90499 1343
rect 92029 1309 92063 1343
rect 93317 1309 93351 1343
rect 94881 1309 94915 1343
rect 94973 1309 95007 1343
rect 95893 1309 95927 1343
rect 96905 1309 96939 1343
rect 97641 1309 97675 1343
rect 98561 1309 98595 1343
rect 98745 1309 98779 1343
rect 99297 1309 99331 1343
rect 100125 1309 100159 1343
rect 100309 1309 100343 1343
rect 100769 1309 100803 1343
rect 103897 1309 103931 1343
rect 104909 1309 104943 1343
rect 105645 1309 105679 1343
rect 106381 1309 106415 1343
rect 107761 1309 107795 1343
rect 108405 1309 108439 1343
rect 109049 1309 109083 1343
rect 110061 1309 110095 1343
rect 110797 1309 110831 1343
rect 111533 1309 111567 1343
rect 112913 1309 112947 1343
rect 113557 1309 113591 1343
rect 114201 1309 114235 1343
rect 115213 1309 115247 1343
rect 115949 1309 115983 1343
rect 116685 1309 116719 1343
rect 118065 1309 118099 1343
rect 118709 1309 118743 1343
rect 119353 1309 119387 1343
rect 120365 1309 120399 1343
rect 121101 1309 121135 1343
rect 121653 1309 121687 1343
rect 122941 1309 122975 1343
rect 123769 1309 123803 1343
rect 125425 1309 125459 1343
rect 126805 1309 126839 1343
rect 128277 1309 128311 1343
rect 128461 1309 128495 1343
rect 128645 1309 128679 1343
rect 129105 1309 129139 1343
rect 130669 1309 130703 1343
rect 131957 1309 131991 1343
rect 132969 1309 133003 1343
rect 133153 1309 133187 1343
rect 133981 1309 134015 1343
rect 134165 1309 134199 1343
rect 138765 1309 138799 1343
rect 139409 1309 139443 1343
rect 140697 1309 140731 1343
rect 141341 1309 141375 1343
rect 141985 1309 142019 1343
rect 143273 1309 143307 1343
rect 143917 1309 143951 1343
rect 144561 1309 144595 1343
rect 145849 1309 145883 1343
rect 146493 1309 146527 1343
rect 147137 1309 147171 1343
rect 148425 1309 148459 1343
rect 149069 1309 149103 1343
rect 149713 1309 149747 1343
rect 151001 1309 151035 1343
rect 151645 1309 151679 1343
rect 152289 1309 152323 1343
rect 153577 1309 153611 1343
rect 154221 1309 154255 1343
rect 154865 1309 154899 1343
rect 156429 1309 156463 1343
rect 156613 1309 156647 1343
rect 157441 1309 157475 1343
rect 158729 1309 158763 1343
rect 159557 1309 159591 1343
rect 159741 1309 159775 1343
rect 160201 1309 160235 1343
rect 161121 1309 161155 1343
rect 162317 1309 162351 1343
rect 163881 1309 163915 1343
rect 164065 1309 164099 1343
rect 164525 1309 164559 1343
rect 167193 1309 167227 1343
rect 167377 1309 167411 1343
rect 167837 1309 167871 1343
rect 168849 1309 168883 1343
rect 172253 1309 172287 1343
rect 172529 1309 172563 1343
rect 174001 1309 174035 1343
rect 174277 1309 174311 1343
rect 176577 1309 176611 1343
rect 176853 1309 176887 1343
rect 179153 1309 179187 1343
rect 179429 1309 179463 1343
rect 182557 1309 182591 1343
rect 182833 1309 182867 1343
rect 184305 1309 184339 1343
rect 184581 1309 184615 1343
rect 186881 1309 186915 1343
rect 187157 1309 187191 1343
rect 189457 1309 189491 1343
rect 189733 1309 189767 1343
rect 191113 1309 191147 1343
rect 191205 1309 191239 1343
rect 192493 1309 192527 1343
rect 193321 1309 193355 1343
rect 194609 1309 194643 1343
rect 195621 1309 195655 1343
rect 197185 1309 197219 1343
rect 197921 1309 197955 1343
rect 199761 1309 199795 1343
rect 200497 1309 200531 1343
rect 201417 1309 201451 1343
rect 202521 1309 202555 1343
rect 202705 1309 202739 1343
rect 203165 1309 203199 1343
rect 206569 1309 206603 1343
rect 207673 1309 207707 1343
rect 208317 1309 208351 1343
rect 208961 1309 208995 1343
rect 210249 1309 210283 1343
rect 210893 1309 210927 1343
rect 211537 1309 211571 1343
rect 212825 1309 212859 1343
rect 213469 1309 213503 1343
rect 214113 1309 214147 1343
rect 215401 1309 215435 1343
rect 216045 1309 216079 1343
rect 216689 1309 216723 1343
rect 217793 1309 217827 1343
rect 218713 1309 218747 1343
rect 219817 1309 219851 1343
rect 220553 1309 220587 1343
rect 221197 1309 221231 1343
rect 221841 1309 221875 1343
rect 223129 1309 223163 1343
rect 223773 1309 223807 1343
rect 224877 1309 224911 1343
rect 225705 1309 225739 1343
rect 226717 1309 226751 1343
rect 226901 1309 226935 1343
rect 228281 1309 228315 1343
rect 228925 1309 228959 1343
rect 229661 1309 229695 1343
rect 230673 1309 230707 1343
rect 232329 1309 232363 1343
rect 233249 1309 233283 1343
rect 233985 1309 234019 1343
rect 234721 1309 234755 1343
rect 236009 1309 236043 1343
rect 240977 1309 241011 1343
rect 241253 1309 241287 1343
rect 243553 1309 243587 1343
rect 243829 1309 243863 1343
rect 246129 1309 246163 1343
rect 246405 1309 246439 1343
rect 248705 1309 248739 1343
rect 248981 1309 249015 1343
rect 251557 1309 251591 1343
rect 251833 1309 251867 1343
rect 253857 1309 253891 1343
rect 254133 1309 254167 1343
rect 256433 1309 256467 1343
rect 256709 1309 256743 1343
rect 257905 1309 257939 1343
rect 258089 1309 258123 1343
rect 259009 1309 259043 1343
rect 259285 1309 259319 1343
rect 260297 1309 260331 1343
rect 261585 1309 261619 1343
rect 262321 1309 262355 1343
rect 263057 1309 263091 1343
rect 264161 1309 264195 1343
rect 265173 1309 265207 1343
rect 265909 1309 265943 1343
rect 266737 1309 266771 1343
rect 267473 1309 267507 1343
rect 268209 1309 268243 1343
rect 269497 1309 269531 1343
rect 269681 1309 269715 1343
rect 270141 1309 270175 1343
rect 4077 1241 4111 1275
rect 8309 1241 8343 1275
rect 9689 1241 9723 1275
rect 10241 1241 10275 1275
rect 10425 1241 10459 1275
rect 10977 1241 11011 1275
rect 11989 1241 12023 1275
rect 12725 1241 12759 1275
rect 13461 1241 13495 1275
rect 17141 1241 17175 1275
rect 17877 1241 17911 1275
rect 18613 1241 18647 1275
rect 25329 1241 25363 1275
rect 25881 1241 25915 1275
rect 54309 1241 54343 1275
rect 180533 1241 180567 1275
rect 181821 1241 181855 1275
rect 218069 1241 218103 1275
rect 218989 1241 219023 1275
rect 224049 1241 224083 1275
rect 247969 1241 248003 1275
rect 250177 1241 250211 1275
rect 4169 1173 4203 1207
rect 8401 1173 8435 1207
rect 12817 1173 12851 1207
rect 13553 1173 13587 1207
rect 17233 1173 17267 1207
rect 17969 1173 18003 1207
rect 18705 1173 18739 1207
rect 23949 1173 23983 1207
rect 29101 1173 29135 1207
rect 29929 1173 29963 1207
rect 30757 1173 30791 1207
rect 31585 1173 31619 1207
rect 32505 1173 32539 1207
rect 36093 1173 36127 1207
rect 38025 1173 38059 1207
rect 39313 1173 39347 1207
rect 40601 1173 40635 1207
rect 41245 1173 41279 1207
rect 41889 1173 41923 1207
rect 43085 1173 43119 1207
rect 43821 1173 43855 1207
rect 45753 1173 45787 1207
rect 46397 1173 46431 1207
rect 47041 1173 47075 1207
rect 48237 1173 48271 1207
rect 48973 1173 49007 1207
rect 49617 1173 49651 1207
rect 50905 1173 50939 1207
rect 51549 1173 51583 1207
rect 52193 1173 52227 1207
rect 53389 1173 53423 1207
rect 56241 1173 56275 1207
rect 57069 1173 57103 1207
rect 58633 1173 58667 1207
rect 60841 1173 60875 1207
rect 61577 1173 61611 1207
rect 62313 1173 62347 1207
rect 63785 1173 63819 1207
rect 64521 1173 64555 1207
rect 66177 1173 66211 1207
rect 90649 1173 90683 1207
rect 92213 1173 92247 1207
rect 93501 1173 93535 1207
rect 96077 1173 96111 1207
rect 97089 1173 97123 1207
rect 97825 1173 97859 1207
rect 100953 1173 100987 1207
rect 103713 1173 103747 1207
rect 104725 1173 104759 1207
rect 105461 1173 105495 1207
rect 106197 1173 106231 1207
rect 107577 1173 107611 1207
rect 108221 1173 108255 1207
rect 108865 1173 108899 1207
rect 109877 1173 109911 1207
rect 110613 1173 110647 1207
rect 111349 1173 111383 1207
rect 112729 1173 112763 1207
rect 114017 1173 114051 1207
rect 115029 1173 115063 1207
rect 115765 1173 115799 1207
rect 116501 1173 116535 1207
rect 117881 1173 117915 1207
rect 118525 1173 118559 1207
rect 119169 1173 119203 1207
rect 120181 1173 120215 1207
rect 120917 1173 120951 1207
rect 121837 1173 121871 1207
rect 123125 1173 123159 1207
rect 123953 1173 123987 1207
rect 125609 1173 125643 1207
rect 126989 1173 127023 1207
rect 129289 1173 129323 1207
rect 130853 1173 130887 1207
rect 132141 1173 132175 1207
rect 138581 1173 138615 1207
rect 141157 1173 141191 1207
rect 141801 1173 141835 1207
rect 143089 1173 143123 1207
rect 143733 1173 143767 1207
rect 144377 1173 144411 1207
rect 145665 1173 145699 1207
rect 146309 1173 146343 1207
rect 146953 1173 146987 1207
rect 148241 1173 148275 1207
rect 148885 1173 148919 1207
rect 149529 1173 149563 1207
rect 150817 1173 150851 1207
rect 151461 1173 151495 1207
rect 152105 1173 152139 1207
rect 153393 1173 153427 1207
rect 154037 1173 154071 1207
rect 154681 1173 154715 1207
rect 158913 1173 158947 1207
rect 160385 1173 160419 1207
rect 161305 1173 161339 1207
rect 162501 1173 162535 1207
rect 164709 1173 164743 1207
rect 168021 1173 168055 1207
rect 169033 1173 169067 1207
rect 181913 1173 181947 1207
rect 192677 1173 192711 1207
rect 193505 1173 193539 1207
rect 194793 1173 194827 1207
rect 195805 1173 195839 1207
rect 197369 1173 197403 1207
rect 198105 1173 198139 1207
rect 199945 1173 199979 1207
rect 200681 1173 200715 1207
rect 201601 1173 201635 1207
rect 203349 1173 203383 1207
rect 206385 1173 206419 1207
rect 207489 1173 207523 1207
rect 208133 1173 208167 1207
rect 208777 1173 208811 1207
rect 210065 1173 210099 1207
rect 210709 1173 210743 1207
rect 211353 1173 211387 1207
rect 212641 1173 212675 1207
rect 213929 1173 213963 1207
rect 215217 1173 215251 1207
rect 215861 1173 215895 1207
rect 216505 1173 216539 1207
rect 219633 1173 219667 1207
rect 220369 1173 220403 1207
rect 221013 1173 221047 1207
rect 222945 1173 222979 1207
rect 224693 1173 224727 1207
rect 229109 1173 229143 1207
rect 229845 1173 229879 1207
rect 230857 1173 230891 1207
rect 233433 1173 233467 1207
rect 234169 1173 234203 1207
rect 234905 1173 234939 1207
rect 248061 1173 248095 1207
rect 250269 1173 250303 1207
rect 260481 1173 260515 1207
rect 261769 1173 261803 1207
rect 262505 1173 262539 1207
rect 263241 1173 263275 1207
rect 264345 1173 264379 1207
rect 265357 1173 265391 1207
rect 266093 1173 266127 1207
rect 266921 1173 266955 1207
rect 267657 1173 267691 1207
rect 268393 1173 268427 1207
rect 270325 1173 270359 1207
<< metal1 >>
rect 97626 10860 97632 10872
rect 90744 10832 97632 10860
rect 90744 10792 90772 10832
rect 97626 10820 97632 10832
rect 97684 10820 97690 10872
rect 98454 10820 98460 10872
rect 98512 10860 98518 10872
rect 98512 10832 109034 10860
rect 98512 10820 98518 10832
rect 64846 10764 90772 10792
rect 28442 10684 28448 10736
rect 28500 10724 28506 10736
rect 33778 10724 33784 10736
rect 28500 10696 33784 10724
rect 28500 10684 28506 10696
rect 33778 10684 33784 10696
rect 33836 10684 33842 10736
rect 29914 10616 29920 10668
rect 29972 10656 29978 10668
rect 63218 10656 63224 10668
rect 29972 10628 30328 10656
rect 29972 10616 29978 10628
rect 23934 10548 23940 10600
rect 23992 10588 23998 10600
rect 30300 10588 30328 10628
rect 38626 10628 63224 10656
rect 38626 10588 38654 10628
rect 63218 10616 63224 10628
rect 63276 10656 63282 10668
rect 64846 10656 64874 10764
rect 90818 10752 90824 10804
rect 90876 10792 90882 10804
rect 95050 10792 95056 10804
rect 90876 10764 95056 10792
rect 90876 10752 90882 10764
rect 95050 10752 95056 10764
rect 95108 10792 95114 10804
rect 96982 10792 96988 10804
rect 95108 10764 96988 10792
rect 95108 10752 95114 10764
rect 96982 10752 96988 10764
rect 97040 10752 97046 10804
rect 109006 10792 109034 10832
rect 152366 10820 152372 10872
rect 152424 10860 152430 10872
rect 163958 10860 163964 10872
rect 152424 10832 163964 10860
rect 152424 10820 152430 10832
rect 163958 10820 163964 10832
rect 164016 10820 164022 10872
rect 214282 10820 214288 10872
rect 214340 10860 214346 10872
rect 227438 10860 227444 10872
rect 214340 10832 227444 10860
rect 214340 10820 214346 10832
rect 227438 10820 227444 10832
rect 227496 10820 227502 10872
rect 229094 10820 229100 10872
rect 229152 10860 229158 10872
rect 233602 10860 233608 10872
rect 229152 10832 233608 10860
rect 229152 10820 229158 10832
rect 233602 10820 233608 10832
rect 233660 10820 233666 10872
rect 233694 10820 233700 10872
rect 233752 10860 233758 10872
rect 246758 10860 246764 10872
rect 233752 10832 246764 10860
rect 233752 10820 233758 10832
rect 246758 10820 246764 10832
rect 246816 10820 246822 10872
rect 258534 10820 258540 10872
rect 258592 10860 258598 10872
rect 267826 10860 267832 10872
rect 258592 10832 267832 10860
rect 258592 10820 258598 10832
rect 267826 10820 267832 10832
rect 267884 10820 267890 10872
rect 132862 10792 132868 10804
rect 109006 10764 132868 10792
rect 132862 10752 132868 10764
rect 132920 10792 132926 10804
rect 133690 10792 133696 10804
rect 132920 10764 133696 10792
rect 132920 10752 132926 10764
rect 133690 10752 133696 10764
rect 133748 10752 133754 10804
rect 152458 10752 152464 10804
rect 152516 10792 152522 10804
rect 164142 10792 164148 10804
rect 152516 10764 164148 10792
rect 152516 10752 152522 10764
rect 164142 10752 164148 10764
rect 164200 10752 164206 10804
rect 164326 10752 164332 10804
rect 164384 10792 164390 10804
rect 239398 10792 239404 10804
rect 164384 10764 239404 10792
rect 164384 10752 164390 10764
rect 239398 10752 239404 10764
rect 239456 10752 239462 10804
rect 255682 10752 255688 10804
rect 255740 10792 255746 10804
rect 267734 10792 267740 10804
rect 255740 10764 267740 10792
rect 255740 10752 255746 10764
rect 267734 10752 267740 10764
rect 267792 10752 267798 10804
rect 65978 10684 65984 10736
rect 66036 10724 66042 10736
rect 99374 10724 99380 10736
rect 66036 10696 99380 10724
rect 66036 10684 66042 10696
rect 99374 10684 99380 10696
rect 99432 10724 99438 10736
rect 104342 10724 104348 10736
rect 99432 10696 104348 10724
rect 99432 10684 99438 10696
rect 104342 10684 104348 10696
rect 104400 10684 104406 10736
rect 130562 10684 130568 10736
rect 130620 10724 130626 10736
rect 164602 10724 164608 10736
rect 130620 10696 164608 10724
rect 130620 10684 130626 10696
rect 164602 10684 164608 10696
rect 164660 10684 164666 10736
rect 164786 10684 164792 10736
rect 164844 10724 164850 10736
rect 264790 10724 264796 10736
rect 164844 10696 264796 10724
rect 164844 10684 164850 10696
rect 264790 10684 264796 10696
rect 264848 10684 264854 10736
rect 63276 10628 64874 10656
rect 63276 10616 63282 10628
rect 74994 10616 75000 10668
rect 75052 10656 75058 10668
rect 104802 10656 104808 10668
rect 75052 10628 104808 10656
rect 75052 10616 75058 10628
rect 104802 10616 104808 10628
rect 104860 10616 104866 10668
rect 165338 10656 165344 10668
rect 132466 10628 165344 10656
rect 23992 10560 30236 10588
rect 30300 10560 38654 10588
rect 23992 10548 23998 10560
rect 23750 10480 23756 10532
rect 23808 10520 23814 10532
rect 30006 10520 30012 10532
rect 23808 10492 30012 10520
rect 23808 10480 23814 10492
rect 30006 10480 30012 10492
rect 30064 10480 30070 10532
rect 25774 10412 25780 10464
rect 25832 10452 25838 10464
rect 25832 10424 29316 10452
rect 25832 10412 25838 10424
rect 20714 10344 20720 10396
rect 20772 10384 20778 10396
rect 25958 10384 25964 10396
rect 20772 10356 25964 10384
rect 20772 10344 20778 10356
rect 25958 10344 25964 10356
rect 26016 10344 26022 10396
rect 22830 10276 22836 10328
rect 22888 10316 22894 10328
rect 24946 10316 24952 10328
rect 22888 10288 24952 10316
rect 22888 10276 22894 10288
rect 24946 10276 24952 10288
rect 25004 10316 25010 10328
rect 25004 10288 29224 10316
rect 25004 10276 25010 10288
rect 26050 10208 26056 10260
rect 26108 10248 26114 10260
rect 29086 10248 29092 10260
rect 26108 10220 29092 10248
rect 26108 10208 26114 10220
rect 29086 10208 29092 10220
rect 29144 10208 29150 10260
rect 27614 10180 27620 10192
rect 26804 10152 27620 10180
rect 7650 10072 7656 10124
rect 7708 10112 7714 10124
rect 26694 10112 26700 10124
rect 7708 10084 26700 10112
rect 7708 10072 7714 10084
rect 26694 10072 26700 10084
rect 26752 10072 26758 10124
rect 5902 10004 5908 10056
rect 5960 10044 5966 10056
rect 23658 10044 23664 10056
rect 5960 10016 23664 10044
rect 5960 10004 5966 10016
rect 23658 10004 23664 10016
rect 23716 10004 23722 10056
rect 17310 9936 17316 9988
rect 17368 9976 17374 9988
rect 26804 9976 26832 10152
rect 27614 10140 27620 10152
rect 27672 10140 27678 10192
rect 29196 10112 29224 10288
rect 29288 10248 29316 10424
rect 30208 10316 30236 10560
rect 60366 10548 60372 10600
rect 60424 10588 60430 10600
rect 94958 10588 94964 10600
rect 60424 10560 94964 10588
rect 60424 10548 60430 10560
rect 94958 10548 94964 10560
rect 95016 10548 95022 10600
rect 96982 10548 96988 10600
rect 97040 10588 97046 10600
rect 129458 10588 129464 10600
rect 97040 10560 129464 10588
rect 97040 10548 97046 10560
rect 129458 10548 129464 10560
rect 129516 10548 129522 10600
rect 60090 10480 60096 10532
rect 60148 10520 60154 10532
rect 90818 10520 90824 10532
rect 60148 10492 90824 10520
rect 60148 10480 60154 10492
rect 90818 10480 90824 10492
rect 90876 10480 90882 10532
rect 91002 10480 91008 10532
rect 91060 10520 91066 10532
rect 91060 10492 92520 10520
rect 91060 10480 91066 10492
rect 57146 10412 57152 10464
rect 57204 10452 57210 10464
rect 92382 10452 92388 10464
rect 57204 10424 92388 10452
rect 57204 10412 57210 10424
rect 92382 10412 92388 10424
rect 92440 10412 92446 10464
rect 92492 10452 92520 10492
rect 94038 10480 94044 10532
rect 94096 10520 94102 10532
rect 96706 10520 96712 10532
rect 94096 10492 96712 10520
rect 94096 10480 94102 10492
rect 96706 10480 96712 10492
rect 96764 10520 96770 10532
rect 131114 10520 131120 10532
rect 96764 10492 131120 10520
rect 96764 10480 96770 10492
rect 131114 10480 131120 10492
rect 131172 10520 131178 10532
rect 132466 10520 132494 10628
rect 165338 10616 165344 10628
rect 165396 10616 165402 10668
rect 225322 10616 225328 10668
rect 225380 10656 225386 10668
rect 226426 10656 226432 10668
rect 225380 10628 226432 10656
rect 225380 10616 225386 10628
rect 226426 10616 226432 10628
rect 226484 10656 226490 10668
rect 226484 10628 233556 10656
rect 226484 10616 226490 10628
rect 133690 10548 133696 10600
rect 133748 10588 133754 10600
rect 167086 10588 167092 10600
rect 133748 10560 167092 10588
rect 133748 10548 133754 10560
rect 167086 10548 167092 10560
rect 167144 10548 167150 10600
rect 196710 10548 196716 10600
rect 196768 10588 196774 10600
rect 227530 10588 227536 10600
rect 196768 10560 227536 10588
rect 196768 10548 196774 10560
rect 227530 10548 227536 10560
rect 227588 10548 227594 10600
rect 233418 10588 233424 10600
rect 227640 10560 233424 10588
rect 131172 10492 132494 10520
rect 131172 10480 131178 10492
rect 133782 10480 133788 10532
rect 133840 10520 133846 10532
rect 167730 10520 167736 10532
rect 133840 10492 167736 10520
rect 133840 10480 133846 10492
rect 167730 10480 167736 10492
rect 167788 10480 167794 10532
rect 192478 10480 192484 10532
rect 192536 10520 192542 10532
rect 224586 10520 224592 10532
rect 192536 10492 224592 10520
rect 192536 10480 192542 10492
rect 224586 10480 224592 10492
rect 224644 10520 224650 10532
rect 225414 10520 225420 10532
rect 224644 10492 225420 10520
rect 224644 10480 224650 10492
rect 225414 10480 225420 10492
rect 225472 10520 225478 10532
rect 227640 10520 227668 10560
rect 233418 10548 233424 10560
rect 233476 10548 233482 10600
rect 225472 10492 227668 10520
rect 225472 10480 225478 10492
rect 227714 10480 227720 10532
rect 227772 10520 227778 10532
rect 230842 10520 230848 10532
rect 227772 10492 230848 10520
rect 227772 10480 227778 10492
rect 230842 10480 230848 10492
rect 230900 10480 230906 10532
rect 233528 10520 233556 10628
rect 233786 10616 233792 10668
rect 233844 10656 233850 10668
rect 233844 10628 258672 10656
rect 233844 10616 233850 10628
rect 233602 10548 233608 10600
rect 233660 10588 233666 10600
rect 258350 10588 258356 10600
rect 233660 10560 258356 10588
rect 233660 10548 233666 10560
rect 258350 10548 258356 10560
rect 258408 10548 258414 10600
rect 258644 10588 258672 10628
rect 258718 10616 258724 10668
rect 258776 10656 258782 10668
rect 266814 10656 266820 10668
rect 258776 10628 266820 10656
rect 258776 10616 258782 10628
rect 266814 10616 266820 10628
rect 266872 10616 266878 10668
rect 260190 10588 260196 10600
rect 258644 10560 260196 10588
rect 260190 10548 260196 10560
rect 260248 10548 260254 10600
rect 260282 10548 260288 10600
rect 260340 10588 260346 10600
rect 263134 10588 263140 10600
rect 260340 10560 263140 10588
rect 260340 10548 260346 10560
rect 263134 10548 263140 10560
rect 263192 10548 263198 10600
rect 258442 10520 258448 10532
rect 233528 10492 258448 10520
rect 258442 10480 258448 10492
rect 258500 10480 258506 10532
rect 258810 10480 258816 10532
rect 258868 10520 258874 10532
rect 268194 10520 268200 10532
rect 258868 10492 268200 10520
rect 258868 10480 258874 10492
rect 268194 10480 268200 10492
rect 268252 10480 268258 10532
rect 125042 10452 125048 10464
rect 92492 10424 125048 10452
rect 125042 10412 125048 10424
rect 125100 10412 125106 10464
rect 162302 10412 162308 10464
rect 162360 10452 162366 10464
rect 263594 10452 263600 10464
rect 162360 10424 263600 10452
rect 162360 10412 162366 10424
rect 263594 10412 263600 10424
rect 263652 10412 263658 10464
rect 33778 10344 33784 10396
rect 33836 10384 33842 10396
rect 62390 10384 62396 10396
rect 33836 10356 62396 10384
rect 33836 10344 33842 10356
rect 62390 10344 62396 10356
rect 62448 10384 62454 10396
rect 94038 10384 94044 10396
rect 62448 10356 94044 10384
rect 62448 10344 62454 10356
rect 94038 10344 94044 10356
rect 94096 10344 94102 10396
rect 96430 10384 96436 10396
rect 94148 10356 96436 10384
rect 57146 10316 57152 10328
rect 30208 10288 57152 10316
rect 57146 10276 57152 10288
rect 57204 10276 57210 10328
rect 61470 10276 61476 10328
rect 61528 10316 61534 10328
rect 94148 10316 94176 10356
rect 96430 10344 96436 10356
rect 96488 10344 96494 10396
rect 98362 10384 98368 10396
rect 96586 10356 98368 10384
rect 61528 10288 94176 10316
rect 61528 10276 61534 10288
rect 59630 10248 59636 10260
rect 29288 10220 59636 10248
rect 59630 10208 59636 10220
rect 59688 10208 59694 10260
rect 66070 10208 66076 10260
rect 66128 10248 66134 10260
rect 96586 10248 96614 10356
rect 98362 10344 98368 10356
rect 98420 10384 98426 10396
rect 99282 10384 99288 10396
rect 98420 10356 99288 10384
rect 98420 10344 98426 10356
rect 99282 10344 99288 10356
rect 99340 10384 99346 10396
rect 103514 10384 103520 10396
rect 99340 10356 103520 10384
rect 99340 10344 99346 10356
rect 103514 10344 103520 10356
rect 103572 10344 103578 10396
rect 104342 10344 104348 10396
rect 104400 10384 104406 10396
rect 133966 10384 133972 10396
rect 104400 10356 133972 10384
rect 104400 10344 104406 10356
rect 133966 10344 133972 10356
rect 134024 10344 134030 10396
rect 151722 10344 151728 10396
rect 151780 10384 151786 10396
rect 181990 10384 181996 10396
rect 151780 10356 181996 10384
rect 151780 10344 151786 10356
rect 181990 10344 181996 10356
rect 182048 10344 182054 10396
rect 202782 10344 202788 10396
rect 202840 10384 202846 10396
rect 235718 10384 235724 10396
rect 202840 10356 235724 10384
rect 202840 10344 202846 10356
rect 235718 10344 235724 10356
rect 235776 10344 235782 10396
rect 255866 10344 255872 10396
rect 255924 10384 255930 10396
rect 268010 10384 268016 10396
rect 255924 10356 268016 10384
rect 255924 10344 255930 10356
rect 268010 10344 268016 10356
rect 268068 10344 268074 10396
rect 103330 10316 103336 10328
rect 66128 10220 96614 10248
rect 96816 10288 103336 10316
rect 66128 10208 66134 10220
rect 30374 10140 30380 10192
rect 30432 10180 30438 10192
rect 64046 10180 64052 10192
rect 30432 10152 64052 10180
rect 30432 10140 30438 10152
rect 64046 10140 64052 10152
rect 64104 10140 64110 10192
rect 77478 10140 77484 10192
rect 77536 10180 77542 10192
rect 96816 10180 96844 10288
rect 103330 10276 103336 10288
rect 103388 10276 103394 10328
rect 131850 10316 131856 10328
rect 103440 10288 131856 10316
rect 97626 10208 97632 10260
rect 97684 10248 97690 10260
rect 103440 10248 103468 10288
rect 131850 10276 131856 10288
rect 131908 10316 131914 10328
rect 131908 10288 138014 10316
rect 131908 10276 131914 10288
rect 97684 10220 103468 10248
rect 97684 10208 97690 10220
rect 103514 10208 103520 10260
rect 103572 10248 103578 10260
rect 132954 10248 132960 10260
rect 103572 10220 132960 10248
rect 103572 10208 103578 10220
rect 132954 10208 132960 10220
rect 133012 10248 133018 10260
rect 133782 10248 133788 10260
rect 133012 10220 133788 10248
rect 133012 10208 133018 10220
rect 133782 10208 133788 10220
rect 133840 10208 133846 10260
rect 137986 10248 138014 10288
rect 149054 10276 149060 10328
rect 149112 10316 149118 10328
rect 172514 10316 172520 10328
rect 149112 10288 172520 10316
rect 149112 10276 149118 10288
rect 172514 10276 172520 10288
rect 172572 10276 172578 10328
rect 193214 10276 193220 10328
rect 193272 10316 193278 10328
rect 225322 10316 225328 10328
rect 193272 10288 225328 10316
rect 193272 10276 193278 10288
rect 225322 10276 225328 10288
rect 225380 10276 225386 10328
rect 225506 10276 225512 10328
rect 225564 10316 225570 10328
rect 227714 10316 227720 10328
rect 225564 10288 227720 10316
rect 225564 10276 225570 10288
rect 227714 10276 227720 10288
rect 227772 10276 227778 10328
rect 228082 10276 228088 10328
rect 228140 10316 228146 10328
rect 228140 10288 230796 10316
rect 228140 10276 228146 10288
rect 166258 10248 166264 10260
rect 137986 10220 166264 10248
rect 166258 10208 166264 10220
rect 166316 10208 166322 10260
rect 170306 10208 170312 10260
rect 170364 10248 170370 10260
rect 208394 10248 208400 10260
rect 170364 10220 208400 10248
rect 170364 10208 170370 10220
rect 208394 10208 208400 10220
rect 208452 10208 208458 10260
rect 215266 10220 218284 10248
rect 77536 10152 96844 10180
rect 77536 10140 77542 10152
rect 97534 10140 97540 10192
rect 97592 10180 97598 10192
rect 103698 10180 103704 10192
rect 97592 10152 103704 10180
rect 97592 10140 97598 10152
rect 103698 10140 103704 10152
rect 103756 10140 103762 10192
rect 122742 10140 122748 10192
rect 122800 10180 122806 10192
rect 156506 10180 156512 10192
rect 122800 10152 156512 10180
rect 122800 10140 122806 10152
rect 156506 10140 156512 10152
rect 156564 10140 156570 10192
rect 162210 10140 162216 10192
rect 162268 10180 162274 10192
rect 215266 10180 215294 10220
rect 162268 10152 215294 10180
rect 218256 10180 218284 10220
rect 218330 10208 218336 10260
rect 218388 10248 218394 10260
rect 230658 10248 230664 10260
rect 218388 10220 230664 10248
rect 218388 10208 218394 10220
rect 230658 10208 230664 10220
rect 230716 10208 230722 10260
rect 230768 10248 230796 10288
rect 230842 10276 230848 10328
rect 230900 10316 230906 10328
rect 258166 10316 258172 10328
rect 230900 10288 258172 10316
rect 230900 10276 230906 10288
rect 258166 10276 258172 10288
rect 258224 10276 258230 10328
rect 258626 10276 258632 10328
rect 258684 10316 258690 10328
rect 266630 10316 266636 10328
rect 258684 10288 266636 10316
rect 258684 10276 258690 10288
rect 266630 10276 266636 10288
rect 266688 10276 266694 10328
rect 258350 10248 258356 10260
rect 230768 10220 258356 10248
rect 258350 10208 258356 10220
rect 258408 10208 258414 10260
rect 258902 10208 258908 10260
rect 258960 10248 258966 10260
rect 266998 10248 267004 10260
rect 258960 10220 267004 10248
rect 258960 10208 258966 10220
rect 266998 10208 267004 10220
rect 267056 10208 267062 10260
rect 262858 10180 262864 10192
rect 218256 10152 262864 10180
rect 162268 10140 162274 10152
rect 262858 10140 262864 10152
rect 262916 10140 262922 10192
rect 270402 10180 270408 10192
rect 262968 10152 270408 10180
rect 17368 9948 26832 9976
rect 26896 10084 27108 10112
rect 29196 10084 41414 10112
rect 17368 9936 17374 9948
rect 8478 9868 8484 9920
rect 8536 9908 8542 9920
rect 26896 9908 26924 10084
rect 27080 10044 27108 10084
rect 33042 10044 33048 10056
rect 27080 10016 33048 10044
rect 33042 10004 33048 10016
rect 33100 10004 33106 10056
rect 41386 10044 41414 10084
rect 56410 10072 56416 10124
rect 56468 10112 56474 10124
rect 91002 10112 91008 10124
rect 56468 10084 91008 10112
rect 56468 10072 56474 10084
rect 91002 10072 91008 10084
rect 91060 10072 91066 10124
rect 93210 10072 93216 10124
rect 93268 10112 93274 10124
rect 126698 10112 126704 10124
rect 93268 10084 126704 10112
rect 93268 10072 93274 10084
rect 126698 10072 126704 10084
rect 126756 10112 126762 10124
rect 126756 10084 128354 10112
rect 126756 10072 126762 10084
rect 55398 10044 55404 10056
rect 41386 10016 55404 10044
rect 55398 10004 55404 10016
rect 55456 10004 55462 10056
rect 92382 10004 92388 10056
rect 92440 10044 92446 10056
rect 102410 10044 102416 10056
rect 92440 10016 102416 10044
rect 92440 10004 92446 10016
rect 102410 10004 102416 10016
rect 102468 10004 102474 10056
rect 122742 10044 122748 10056
rect 102520 10016 122748 10044
rect 27062 9936 27068 9988
rect 27120 9976 27126 9988
rect 28994 9976 29000 9988
rect 27120 9948 29000 9976
rect 27120 9936 27126 9948
rect 28994 9936 29000 9948
rect 29052 9936 29058 9988
rect 31202 9936 31208 9988
rect 31260 9976 31266 9988
rect 64966 9976 64972 9988
rect 31260 9948 64972 9976
rect 31260 9936 31266 9948
rect 64966 9936 64972 9948
rect 65024 9976 65030 9988
rect 66070 9976 66076 9988
rect 65024 9948 66076 9976
rect 65024 9936 65030 9948
rect 66070 9936 66076 9948
rect 66128 9936 66134 9988
rect 76742 9936 76748 9988
rect 76800 9976 76806 9988
rect 101674 9976 101680 9988
rect 76800 9948 101680 9976
rect 76800 9936 76806 9948
rect 101674 9936 101680 9948
rect 101732 9936 101738 9988
rect 102520 9976 102548 10016
rect 122742 10004 122748 10016
rect 122800 10004 122806 10056
rect 128326 10044 128354 10084
rect 158622 10072 158628 10124
rect 158680 10112 158686 10124
rect 182450 10112 182456 10124
rect 158680 10084 182456 10112
rect 158680 10072 158686 10084
rect 182450 10072 182456 10084
rect 182508 10072 182514 10124
rect 198642 10072 198648 10124
rect 198700 10112 198706 10124
rect 218146 10112 218152 10124
rect 198700 10084 218152 10112
rect 198700 10072 198706 10084
rect 218146 10072 218152 10084
rect 218204 10072 218210 10124
rect 218238 10072 218244 10124
rect 218296 10112 218302 10124
rect 225506 10112 225512 10124
rect 218296 10084 225512 10112
rect 218296 10072 218302 10084
rect 225506 10072 225512 10084
rect 225564 10072 225570 10124
rect 225598 10072 225604 10124
rect 225656 10112 225662 10124
rect 233694 10112 233700 10124
rect 225656 10084 233700 10112
rect 225656 10072 225662 10084
rect 233694 10072 233700 10084
rect 233752 10112 233758 10124
rect 258626 10112 258632 10124
rect 233752 10084 258632 10112
rect 233752 10072 233758 10084
rect 258626 10072 258632 10084
rect 258684 10072 258690 10124
rect 262398 10072 262404 10124
rect 262456 10112 262462 10124
rect 262968 10112 262996 10152
rect 270402 10140 270408 10152
rect 270460 10140 270466 10192
rect 262456 10084 262996 10112
rect 262456 10072 262462 10084
rect 263318 10072 263324 10124
rect 263376 10112 263382 10124
rect 268930 10112 268936 10124
rect 263376 10084 268936 10112
rect 263376 10072 263382 10084
rect 268930 10072 268936 10084
rect 268988 10072 268994 10124
rect 160922 10044 160928 10056
rect 128326 10016 160928 10044
rect 160922 10004 160928 10016
rect 160980 10004 160986 10056
rect 163682 10004 163688 10056
rect 163740 10044 163746 10056
rect 243078 10044 243084 10056
rect 163740 10016 243084 10044
rect 163740 10004 163746 10016
rect 243078 10004 243084 10016
rect 243136 10004 243142 10056
rect 257982 10004 257988 10056
rect 258040 10044 258046 10056
rect 265894 10044 265900 10056
rect 258040 10016 265900 10044
rect 258040 10004 258046 10016
rect 265894 10004 265900 10016
rect 265952 10004 265958 10056
rect 266262 10004 266268 10056
rect 266320 10044 266326 10056
rect 269022 10044 269028 10056
rect 266320 10016 269028 10044
rect 266320 10004 266326 10016
rect 269022 10004 269028 10016
rect 269080 10004 269086 10056
rect 102336 9948 102548 9976
rect 8536 9880 26924 9908
rect 8536 9868 8542 9880
rect 26970 9868 26976 9920
rect 27028 9908 27034 9920
rect 31846 9908 31852 9920
rect 27028 9880 31852 9908
rect 27028 9868 27034 9880
rect 31846 9868 31852 9880
rect 31904 9868 31910 9920
rect 58894 9868 58900 9920
rect 58952 9908 58958 9920
rect 92842 9908 92848 9920
rect 58952 9880 92848 9908
rect 58952 9868 58958 9880
rect 92842 9868 92848 9880
rect 92900 9868 92906 9920
rect 92934 9868 92940 9920
rect 92992 9908 92998 9920
rect 102336 9908 102364 9948
rect 124122 9936 124128 9988
rect 124180 9976 124186 9988
rect 158714 9976 158720 9988
rect 124180 9948 158720 9976
rect 124180 9936 124186 9948
rect 158714 9936 158720 9948
rect 158772 9936 158778 9988
rect 162578 9976 162584 9988
rect 161400 9948 162584 9976
rect 161400 9920 161428 9948
rect 162578 9936 162584 9948
rect 162636 9936 162642 9988
rect 165246 9936 165252 9988
rect 165304 9976 165310 9988
rect 258718 9976 258724 9988
rect 165304 9948 258724 9976
rect 165304 9936 165310 9948
rect 258718 9936 258724 9948
rect 258776 9936 258782 9988
rect 261018 9936 261024 9988
rect 261076 9976 261082 9988
rect 267918 9976 267924 9988
rect 261076 9948 267924 9976
rect 261076 9936 261082 9948
rect 267918 9936 267924 9948
rect 267976 9936 267982 9988
rect 92992 9880 102364 9908
rect 92992 9868 92998 9880
rect 102410 9868 102416 9920
rect 102468 9908 102474 9920
rect 113818 9908 113824 9920
rect 102468 9880 113824 9908
rect 102468 9868 102474 9880
rect 113818 9868 113824 9880
rect 113876 9868 113882 9920
rect 121270 9868 121276 9920
rect 121328 9908 121334 9920
rect 127618 9908 127624 9920
rect 121328 9880 127624 9908
rect 121328 9868 121334 9880
rect 127618 9868 127624 9880
rect 127676 9908 127682 9920
rect 161382 9908 161388 9920
rect 127676 9880 161388 9908
rect 127676 9868 127682 9880
rect 161382 9868 161388 9880
rect 161440 9868 161446 9920
rect 163590 9868 163596 9920
rect 163648 9908 163654 9920
rect 187050 9908 187056 9920
rect 163648 9880 187056 9908
rect 163648 9868 163654 9880
rect 187050 9868 187056 9880
rect 187108 9868 187114 9920
rect 199654 9868 199660 9920
rect 199712 9908 199718 9920
rect 229186 9908 229192 9920
rect 199712 9880 229192 9908
rect 199712 9868 199718 9880
rect 229186 9868 229192 9880
rect 229244 9868 229250 9920
rect 229462 9868 229468 9920
rect 229520 9908 229526 9920
rect 263962 9908 263968 9920
rect 229520 9880 263968 9908
rect 229520 9868 229526 9880
rect 263962 9868 263968 9880
rect 264020 9868 264026 9920
rect 264974 9868 264980 9920
rect 265032 9908 265038 9920
rect 268470 9908 268476 9920
rect 265032 9880 268476 9908
rect 265032 9868 265038 9880
rect 268470 9868 268476 9880
rect 268528 9868 268534 9920
rect 1104 9818 271651 9840
rect 1104 9766 68546 9818
rect 68598 9766 68610 9818
rect 68662 9766 68674 9818
rect 68726 9766 68738 9818
rect 68790 9766 68802 9818
rect 68854 9766 136143 9818
rect 136195 9766 136207 9818
rect 136259 9766 136271 9818
rect 136323 9766 136335 9818
rect 136387 9766 136399 9818
rect 136451 9766 203740 9818
rect 203792 9766 203804 9818
rect 203856 9766 203868 9818
rect 203920 9766 203932 9818
rect 203984 9766 203996 9818
rect 204048 9766 271337 9818
rect 271389 9766 271401 9818
rect 271453 9766 271465 9818
rect 271517 9766 271529 9818
rect 271581 9766 271593 9818
rect 271645 9766 271651 9818
rect 1104 9744 271651 9766
rect 5902 9664 5908 9716
rect 5960 9664 5966 9716
rect 7650 9664 7656 9716
rect 7708 9664 7714 9716
rect 8478 9664 8484 9716
rect 8536 9664 8542 9716
rect 16209 9707 16267 9713
rect 16209 9673 16221 9707
rect 16255 9704 16267 9707
rect 51074 9704 51080 9716
rect 16255 9676 51080 9704
rect 16255 9673 16267 9676
rect 16209 9667 16267 9673
rect 51074 9664 51080 9676
rect 51132 9664 51138 9716
rect 54662 9664 54668 9716
rect 54720 9664 54726 9716
rect 57790 9664 57796 9716
rect 57848 9704 57854 9716
rect 58253 9707 58311 9713
rect 58253 9704 58265 9707
rect 57848 9676 58265 9704
rect 57848 9664 57854 9676
rect 58253 9673 58265 9676
rect 58299 9673 58311 9707
rect 58253 9667 58311 9673
rect 59262 9664 59268 9716
rect 59320 9664 59326 9716
rect 59998 9664 60004 9716
rect 60056 9664 60062 9716
rect 60826 9664 60832 9716
rect 60884 9664 60890 9716
rect 63402 9664 63408 9716
rect 63460 9664 63466 9716
rect 66162 9664 66168 9716
rect 66220 9664 66226 9716
rect 66898 9664 66904 9716
rect 66956 9664 66962 9716
rect 69799 9707 69857 9713
rect 69799 9673 69811 9707
rect 69845 9704 69857 9707
rect 90266 9704 90272 9716
rect 69845 9676 90272 9704
rect 69845 9673 69857 9676
rect 69799 9667 69857 9673
rect 90266 9664 90272 9676
rect 90324 9664 90330 9716
rect 90358 9664 90364 9716
rect 90416 9664 90422 9716
rect 93486 9664 93492 9716
rect 93544 9664 93550 9716
rect 95970 9664 95976 9716
rect 96028 9664 96034 9716
rect 96338 9664 96344 9716
rect 96396 9704 96402 9716
rect 96893 9707 96951 9713
rect 96893 9704 96905 9707
rect 96396 9676 96905 9704
rect 96396 9664 96402 9676
rect 96893 9673 96905 9676
rect 96939 9673 96951 9707
rect 96893 9667 96951 9673
rect 97994 9664 98000 9716
rect 98052 9704 98058 9716
rect 98181 9707 98239 9713
rect 98181 9704 98193 9707
rect 98052 9676 98193 9704
rect 98052 9664 98058 9676
rect 98181 9673 98193 9676
rect 98227 9673 98239 9707
rect 98181 9667 98239 9673
rect 98270 9664 98276 9716
rect 98328 9704 98334 9716
rect 98328 9676 100616 9704
rect 98328 9664 98334 9676
rect 1670 9596 1676 9648
rect 1728 9596 1734 9648
rect 2406 9596 2412 9648
rect 2464 9596 2470 9648
rect 3234 9596 3240 9648
rect 3292 9596 3298 9648
rect 4338 9596 4344 9648
rect 4396 9596 4402 9648
rect 5074 9596 5080 9648
rect 5132 9596 5138 9648
rect 5810 9596 5816 9648
rect 5868 9596 5874 9648
rect 6822 9596 6828 9648
rect 6880 9596 6886 9648
rect 7558 9596 7564 9648
rect 7616 9596 7622 9648
rect 8386 9596 8392 9648
rect 8444 9596 8450 9648
rect 11974 9596 11980 9648
rect 12032 9596 12038 9648
rect 12710 9596 12716 9648
rect 12768 9596 12774 9648
rect 13541 9639 13599 9645
rect 13541 9605 13553 9639
rect 13587 9636 13599 9639
rect 13722 9636 13728 9648
rect 13587 9608 13728 9636
rect 13587 9605 13599 9608
rect 13541 9599 13599 9605
rect 13722 9596 13728 9608
rect 13780 9596 13786 9648
rect 14642 9596 14648 9648
rect 14700 9596 14706 9648
rect 15378 9596 15384 9648
rect 15436 9596 15442 9648
rect 16114 9596 16120 9648
rect 16172 9596 16178 9648
rect 17126 9596 17132 9648
rect 17184 9596 17190 9648
rect 17310 9596 17316 9648
rect 17368 9596 17374 9648
rect 17862 9596 17868 9648
rect 17920 9596 17926 9648
rect 18598 9596 18604 9648
rect 18656 9596 18662 9648
rect 18785 9639 18843 9645
rect 18785 9605 18797 9639
rect 18831 9636 18843 9639
rect 18831 9608 22324 9636
rect 18831 9605 18843 9608
rect 18785 9599 18843 9605
rect 4525 9571 4583 9577
rect 4525 9537 4537 9571
rect 4571 9568 4583 9571
rect 4571 9540 6914 9568
rect 4571 9537 4583 9540
rect 4525 9531 4583 9537
rect 6886 9500 6914 9540
rect 9674 9528 9680 9580
rect 9732 9528 9738 9580
rect 9876 9558 22140 9568
rect 22296 9558 22324 9608
rect 22370 9596 22376 9648
rect 22428 9636 22434 9648
rect 25501 9639 25559 9645
rect 25501 9636 25513 9639
rect 22428 9608 25513 9636
rect 22428 9596 22434 9608
rect 25501 9605 25513 9608
rect 25547 9605 25559 9639
rect 25501 9599 25559 9605
rect 26605 9639 26663 9645
rect 26605 9605 26617 9639
rect 26651 9636 26663 9639
rect 28902 9636 28908 9648
rect 26651 9608 28908 9636
rect 26651 9605 26663 9608
rect 26605 9599 26663 9605
rect 28902 9596 28908 9608
rect 28960 9596 28966 9648
rect 28994 9596 29000 9648
rect 29052 9636 29058 9648
rect 46198 9636 46204 9648
rect 29052 9608 46204 9636
rect 29052 9596 29058 9608
rect 46198 9596 46204 9608
rect 46256 9596 46262 9648
rect 60090 9636 60096 9648
rect 46400 9608 60096 9636
rect 9876 9540 22232 9558
rect 9876 9500 9904 9540
rect 22112 9530 22232 9540
rect 22296 9530 22416 9558
rect 6886 9472 9904 9500
rect 9950 9460 9956 9512
rect 10008 9460 10014 9512
rect 12161 9503 12219 9509
rect 12161 9469 12173 9503
rect 12207 9500 12219 9503
rect 14734 9500 14740 9512
rect 12207 9472 14740 9500
rect 12207 9469 12219 9472
rect 12161 9463 12219 9469
rect 14734 9460 14740 9472
rect 14792 9460 14798 9512
rect 14829 9503 14887 9509
rect 14829 9469 14841 9503
rect 14875 9500 14887 9503
rect 22204 9500 22232 9530
rect 22388 9500 22416 9530
rect 23566 9528 23572 9580
rect 23624 9568 23630 9580
rect 23750 9568 23756 9580
rect 23624 9540 23756 9568
rect 23624 9528 23630 9540
rect 23750 9528 23756 9540
rect 23808 9528 23814 9580
rect 23842 9528 23848 9580
rect 23900 9528 23906 9580
rect 25130 9528 25136 9580
rect 25188 9528 25194 9580
rect 26421 9571 26479 9577
rect 26421 9537 26433 9571
rect 26467 9568 26479 9571
rect 27522 9568 27528 9580
rect 26467 9540 27528 9568
rect 26467 9537 26479 9540
rect 26421 9531 26479 9537
rect 27522 9528 27528 9540
rect 27580 9568 27586 9580
rect 27985 9571 28043 9577
rect 27985 9568 27997 9571
rect 27580 9540 27997 9568
rect 27580 9528 27586 9540
rect 27985 9537 27997 9540
rect 28031 9537 28043 9571
rect 27985 9531 28043 9537
rect 28629 9571 28687 9577
rect 28629 9537 28641 9571
rect 28675 9568 28687 9571
rect 28718 9568 28724 9580
rect 28675 9540 28724 9568
rect 28675 9537 28687 9540
rect 28629 9531 28687 9537
rect 14875 9472 22094 9500
rect 22204 9472 22324 9500
rect 22388 9472 24624 9500
rect 14875 9469 14887 9472
rect 14829 9463 14887 9469
rect 3418 9392 3424 9444
rect 3476 9392 3482 9444
rect 5261 9435 5319 9441
rect 5261 9401 5273 9435
rect 5307 9432 5319 9435
rect 5307 9404 13676 9432
rect 5307 9401 5319 9404
rect 5261 9395 5319 9401
rect 1765 9367 1823 9373
rect 1765 9333 1777 9367
rect 1811 9364 1823 9367
rect 2406 9364 2412 9376
rect 1811 9336 2412 9364
rect 1811 9333 1823 9336
rect 1765 9327 1823 9333
rect 2406 9324 2412 9336
rect 2464 9324 2470 9376
rect 2498 9324 2504 9376
rect 2556 9324 2562 9376
rect 6914 9324 6920 9376
rect 6972 9324 6978 9376
rect 12802 9324 12808 9376
rect 12860 9324 12866 9376
rect 13648 9364 13676 9404
rect 13722 9392 13728 9444
rect 13780 9392 13786 9444
rect 15562 9392 15568 9444
rect 15620 9392 15626 9444
rect 18049 9435 18107 9441
rect 18049 9401 18061 9435
rect 18095 9432 18107 9435
rect 20346 9432 20352 9444
rect 18095 9404 20352 9432
rect 18095 9401 18107 9404
rect 18049 9395 18107 9401
rect 20346 9392 20352 9404
rect 20404 9392 20410 9444
rect 15286 9364 15292 9376
rect 13648 9336 15292 9364
rect 15286 9324 15292 9336
rect 15344 9324 15350 9376
rect 22066 9364 22094 9472
rect 22296 9432 22324 9472
rect 24394 9432 24400 9444
rect 22296 9404 24400 9432
rect 24394 9392 24400 9404
rect 24452 9392 24458 9444
rect 23382 9364 23388 9376
rect 22066 9336 23388 9364
rect 23382 9324 23388 9336
rect 23440 9324 23446 9376
rect 23750 9324 23756 9376
rect 23808 9364 23814 9376
rect 23934 9364 23940 9376
rect 23808 9336 23940 9364
rect 23808 9324 23814 9336
rect 23934 9324 23940 9336
rect 23992 9324 23998 9376
rect 24029 9367 24087 9373
rect 24029 9333 24041 9367
rect 24075 9364 24087 9367
rect 24486 9364 24492 9376
rect 24075 9336 24492 9364
rect 24075 9333 24087 9336
rect 24029 9327 24087 9333
rect 24486 9324 24492 9336
rect 24544 9324 24550 9376
rect 24596 9364 24624 9472
rect 26050 9460 26056 9512
rect 26108 9500 26114 9512
rect 26237 9503 26295 9509
rect 26237 9500 26249 9503
rect 26108 9472 26249 9500
rect 26108 9460 26114 9472
rect 26237 9469 26249 9472
rect 26283 9469 26295 9503
rect 26237 9463 26295 9469
rect 27706 9460 27712 9512
rect 27764 9500 27770 9512
rect 27801 9503 27859 9509
rect 27801 9500 27813 9503
rect 27764 9472 27813 9500
rect 27764 9460 27770 9472
rect 27801 9469 27813 9472
rect 27847 9469 27859 9503
rect 28000 9500 28028 9531
rect 28718 9528 28724 9540
rect 28776 9528 28782 9580
rect 29730 9528 29736 9580
rect 29788 9528 29794 9580
rect 32401 9571 32459 9577
rect 32401 9537 32413 9571
rect 32447 9568 32459 9571
rect 32674 9568 32680 9580
rect 32447 9540 32680 9568
rect 32447 9537 32459 9540
rect 32401 9531 32459 9537
rect 32674 9528 32680 9540
rect 32732 9528 32738 9580
rect 35618 9528 35624 9580
rect 35676 9528 35682 9580
rect 36262 9528 36268 9580
rect 36320 9528 36326 9580
rect 36906 9528 36912 9580
rect 36964 9528 36970 9580
rect 38102 9528 38108 9580
rect 38160 9528 38166 9580
rect 38838 9528 38844 9580
rect 38896 9528 38902 9580
rect 39482 9528 39488 9580
rect 39540 9528 39546 9580
rect 40770 9528 40776 9580
rect 40828 9528 40834 9580
rect 41414 9528 41420 9580
rect 41472 9528 41478 9580
rect 42058 9528 42064 9580
rect 42116 9528 42122 9580
rect 43254 9528 43260 9580
rect 43312 9528 43318 9580
rect 43990 9528 43996 9580
rect 44048 9528 44054 9580
rect 44634 9528 44640 9580
rect 44692 9528 44698 9580
rect 45922 9528 45928 9580
rect 45980 9528 45986 9580
rect 46400 9568 46428 9608
rect 60090 9596 60096 9608
rect 60148 9596 60154 9648
rect 94130 9636 94136 9648
rect 74506 9608 94136 9636
rect 46216 9540 46428 9568
rect 28994 9500 29000 9512
rect 28000 9472 29000 9500
rect 27801 9463 27859 9469
rect 28994 9460 29000 9472
rect 29052 9460 29058 9512
rect 29086 9460 29092 9512
rect 29144 9500 29150 9512
rect 46216 9500 46244 9540
rect 46566 9528 46572 9580
rect 46624 9528 46630 9580
rect 47210 9528 47216 9580
rect 47268 9528 47274 9580
rect 48222 9528 48228 9580
rect 48280 9568 48286 9580
rect 48409 9571 48467 9577
rect 48409 9568 48421 9571
rect 48280 9540 48421 9568
rect 48280 9528 48286 9540
rect 48409 9537 48421 9540
rect 48455 9537 48467 9571
rect 48409 9531 48467 9537
rect 49142 9528 49148 9580
rect 49200 9528 49206 9580
rect 49786 9528 49792 9580
rect 49844 9528 49850 9580
rect 50614 9528 50620 9580
rect 50672 9528 50678 9580
rect 51350 9528 51356 9580
rect 51408 9528 51414 9580
rect 52086 9528 52092 9580
rect 52144 9528 52150 9580
rect 53006 9528 53012 9580
rect 53064 9528 53070 9580
rect 53837 9571 53895 9577
rect 53837 9537 53849 9571
rect 53883 9568 53895 9571
rect 54018 9568 54024 9580
rect 53883 9540 54024 9568
rect 53883 9537 53895 9540
rect 53837 9531 53895 9537
rect 54018 9528 54024 9540
rect 54076 9528 54082 9580
rect 54110 9528 54116 9580
rect 54168 9568 54174 9580
rect 54481 9571 54539 9577
rect 54481 9568 54493 9571
rect 54168 9540 54493 9568
rect 54168 9528 54174 9540
rect 54481 9537 54493 9540
rect 54527 9537 54539 9571
rect 54481 9531 54539 9537
rect 57514 9528 57520 9580
rect 57572 9568 57578 9580
rect 58069 9571 58127 9577
rect 58069 9568 58081 9571
rect 57572 9540 58081 9568
rect 57572 9528 57578 9540
rect 58069 9537 58081 9540
rect 58115 9537 58127 9571
rect 58069 9531 58127 9537
rect 59081 9571 59139 9577
rect 59081 9537 59093 9571
rect 59127 9568 59139 9571
rect 59170 9568 59176 9580
rect 59127 9540 59176 9568
rect 59127 9537 59139 9540
rect 59081 9531 59139 9537
rect 59170 9528 59176 9540
rect 59228 9528 59234 9580
rect 59817 9571 59875 9577
rect 59817 9537 59829 9571
rect 59863 9568 59875 9571
rect 59998 9568 60004 9580
rect 59863 9540 60004 9568
rect 59863 9537 59875 9540
rect 59817 9531 59875 9537
rect 59998 9528 60004 9540
rect 60056 9528 60062 9580
rect 60645 9571 60703 9577
rect 60645 9537 60657 9571
rect 60691 9568 60703 9571
rect 60734 9568 60740 9580
rect 60691 9540 60740 9568
rect 60691 9537 60703 9540
rect 60645 9531 60703 9537
rect 60734 9528 60740 9540
rect 60792 9528 60798 9580
rect 62758 9528 62764 9580
rect 62816 9568 62822 9580
rect 63221 9571 63279 9577
rect 63221 9568 63233 9571
rect 62816 9540 63233 9568
rect 62816 9528 62822 9540
rect 63221 9537 63233 9540
rect 63267 9537 63279 9571
rect 63221 9531 63279 9537
rect 65981 9571 66039 9577
rect 65981 9537 65993 9571
rect 66027 9568 66039 9571
rect 66346 9568 66352 9580
rect 66027 9540 66352 9568
rect 66027 9537 66039 9540
rect 65981 9531 66039 9537
rect 66346 9528 66352 9540
rect 66404 9528 66410 9580
rect 66717 9571 66775 9577
rect 66717 9537 66729 9571
rect 66763 9568 66775 9571
rect 66990 9568 66996 9580
rect 66763 9540 66996 9568
rect 66763 9537 66775 9540
rect 66717 9531 66775 9537
rect 66990 9528 66996 9540
rect 67048 9528 67054 9580
rect 69106 9528 69112 9580
rect 69164 9528 69170 9580
rect 69569 9571 69627 9577
rect 69569 9537 69581 9571
rect 69615 9568 69627 9571
rect 70302 9568 70308 9580
rect 69615 9540 70308 9568
rect 69615 9537 69627 9540
rect 69569 9531 69627 9537
rect 70302 9528 70308 9540
rect 70360 9528 70366 9580
rect 72142 9528 72148 9580
rect 72200 9528 72206 9580
rect 72421 9571 72479 9577
rect 72421 9537 72433 9571
rect 72467 9568 72479 9571
rect 74506 9568 74534 9608
rect 94130 9596 94136 9608
rect 94188 9596 94194 9648
rect 100588 9636 100616 9676
rect 100662 9664 100668 9716
rect 100720 9664 100726 9716
rect 103698 9664 103704 9716
rect 103756 9664 103762 9716
rect 104710 9664 104716 9716
rect 104768 9664 104774 9716
rect 105446 9664 105452 9716
rect 105504 9664 105510 9716
rect 105906 9664 105912 9716
rect 105964 9704 105970 9716
rect 108853 9707 108911 9713
rect 108853 9704 108865 9707
rect 105964 9676 108865 9704
rect 105964 9664 105970 9676
rect 108853 9673 108865 9676
rect 108899 9673 108911 9707
rect 108853 9667 108911 9673
rect 108942 9664 108948 9716
rect 109000 9704 109006 9716
rect 111337 9707 111395 9713
rect 111337 9704 111349 9707
rect 109000 9676 111349 9704
rect 109000 9664 109006 9676
rect 111337 9673 111349 9676
rect 111383 9673 111395 9707
rect 111337 9667 111395 9673
rect 113818 9664 113824 9716
rect 113876 9704 113882 9716
rect 113876 9676 122604 9704
rect 113876 9664 113882 9676
rect 94240 9608 100156 9636
rect 100588 9608 122420 9636
rect 72467 9540 74534 9568
rect 72467 9537 72479 9540
rect 72421 9531 72479 9537
rect 74718 9528 74724 9580
rect 74776 9528 74782 9580
rect 77294 9528 77300 9580
rect 77352 9528 77358 9580
rect 79873 9571 79931 9577
rect 79873 9537 79885 9571
rect 79919 9568 79931 9571
rect 79962 9568 79968 9580
rect 79919 9540 79968 9568
rect 79919 9537 79931 9540
rect 79873 9531 79931 9537
rect 79962 9528 79968 9540
rect 80020 9528 80026 9580
rect 82449 9571 82507 9577
rect 82449 9537 82461 9571
rect 82495 9568 82507 9571
rect 82630 9568 82636 9580
rect 82495 9540 82636 9568
rect 82495 9537 82507 9540
rect 82449 9531 82507 9537
rect 82630 9528 82636 9540
rect 82688 9528 82694 9580
rect 84562 9528 84568 9580
rect 84620 9528 84626 9580
rect 86770 9528 86776 9580
rect 86828 9528 86834 9580
rect 89162 9528 89168 9580
rect 89220 9568 89226 9580
rect 89257 9571 89315 9577
rect 89257 9568 89269 9571
rect 89220 9540 89269 9568
rect 89220 9528 89226 9540
rect 89257 9537 89269 9540
rect 89303 9537 89315 9571
rect 89257 9531 89315 9537
rect 90174 9528 90180 9580
rect 90232 9528 90238 9580
rect 93305 9571 93363 9577
rect 93305 9537 93317 9571
rect 93351 9568 93363 9571
rect 93670 9568 93676 9580
rect 93351 9540 93676 9568
rect 93351 9537 93363 9540
rect 93305 9531 93363 9537
rect 93670 9528 93676 9540
rect 93728 9528 93734 9580
rect 29144 9472 46244 9500
rect 29144 9460 29150 9472
rect 46290 9460 46296 9512
rect 46348 9500 46354 9512
rect 53377 9503 53435 9509
rect 53377 9500 53389 9503
rect 46348 9472 53389 9500
rect 46348 9460 46354 9472
rect 53377 9469 53389 9472
rect 53423 9500 53435 9503
rect 53653 9503 53711 9509
rect 53653 9500 53665 9503
rect 53423 9472 53665 9500
rect 53423 9469 53435 9472
rect 53377 9463 53435 9469
rect 53653 9469 53665 9472
rect 53699 9469 53711 9503
rect 53653 9463 53711 9469
rect 25866 9392 25872 9444
rect 25924 9432 25930 9444
rect 25924 9404 28304 9432
rect 25924 9392 25930 9404
rect 26878 9364 26884 9376
rect 24596 9336 26884 9364
rect 26878 9324 26884 9336
rect 26936 9324 26942 9376
rect 28166 9324 28172 9376
rect 28224 9324 28230 9376
rect 28276 9364 28304 9404
rect 28810 9392 28816 9444
rect 28868 9392 28874 9444
rect 32582 9392 32588 9444
rect 32640 9392 32646 9444
rect 46198 9432 46204 9444
rect 32784 9404 46204 9432
rect 29917 9367 29975 9373
rect 29917 9364 29929 9367
rect 28276 9336 29929 9364
rect 29917 9333 29929 9336
rect 29963 9333 29975 9367
rect 29917 9327 29975 9333
rect 30006 9324 30012 9376
rect 30064 9364 30070 9376
rect 32784 9364 32812 9404
rect 46198 9392 46204 9404
rect 46256 9392 46262 9444
rect 47762 9392 47768 9444
rect 47820 9432 47826 9444
rect 48961 9435 49019 9441
rect 48961 9432 48973 9435
rect 47820 9404 48973 9432
rect 47820 9392 47826 9404
rect 48961 9401 48973 9404
rect 49007 9401 49019 9435
rect 53668 9432 53696 9463
rect 55858 9460 55864 9512
rect 55916 9500 55922 9512
rect 61470 9500 61476 9512
rect 55916 9472 61476 9500
rect 55916 9460 55922 9472
rect 61470 9460 61476 9472
rect 61528 9460 61534 9512
rect 74997 9503 75055 9509
rect 74997 9469 75009 9503
rect 75043 9500 75055 9503
rect 75822 9500 75828 9512
rect 75043 9472 75828 9500
rect 75043 9469 75055 9472
rect 74997 9463 75055 9469
rect 75822 9460 75828 9472
rect 75880 9460 75886 9512
rect 77570 9460 77576 9512
rect 77628 9460 77634 9512
rect 80149 9503 80207 9509
rect 80149 9469 80161 9503
rect 80195 9500 80207 9503
rect 81342 9500 81348 9512
rect 80195 9472 81348 9500
rect 80195 9469 80207 9472
rect 80149 9463 80207 9469
rect 81342 9460 81348 9472
rect 81400 9460 81406 9512
rect 82722 9460 82728 9512
rect 82780 9460 82786 9512
rect 84838 9460 84844 9512
rect 84896 9460 84902 9512
rect 87046 9460 87052 9512
rect 87104 9460 87110 9512
rect 87782 9460 87788 9512
rect 87840 9500 87846 9512
rect 89073 9503 89131 9509
rect 89073 9500 89085 9503
rect 87840 9472 89085 9500
rect 87840 9460 87846 9472
rect 89073 9469 89085 9472
rect 89119 9500 89131 9503
rect 89809 9503 89867 9509
rect 89809 9500 89821 9503
rect 89119 9472 89821 9500
rect 89119 9469 89131 9472
rect 89073 9463 89131 9469
rect 89809 9469 89821 9472
rect 89855 9500 89867 9503
rect 89855 9472 91508 9500
rect 89855 9469 89867 9472
rect 89809 9463 89867 9469
rect 53742 9432 53748 9444
rect 53668 9404 53748 9432
rect 48961 9395 49019 9401
rect 53742 9392 53748 9404
rect 53800 9432 53806 9444
rect 53800 9404 74534 9432
rect 53800 9392 53806 9404
rect 30064 9336 32812 9364
rect 35437 9367 35495 9373
rect 30064 9324 30070 9336
rect 35437 9333 35449 9367
rect 35483 9364 35495 9367
rect 35802 9364 35808 9376
rect 35483 9336 35808 9364
rect 35483 9333 35495 9336
rect 35437 9327 35495 9333
rect 35802 9324 35808 9336
rect 35860 9324 35866 9376
rect 36081 9367 36139 9373
rect 36081 9333 36093 9367
rect 36127 9364 36139 9367
rect 36630 9364 36636 9376
rect 36127 9336 36636 9364
rect 36127 9333 36139 9336
rect 36081 9327 36139 9333
rect 36630 9324 36636 9336
rect 36688 9324 36694 9376
rect 36725 9367 36783 9373
rect 36725 9333 36737 9367
rect 36771 9364 36783 9367
rect 37090 9364 37096 9376
rect 36771 9336 37096 9364
rect 36771 9333 36783 9336
rect 36725 9327 36783 9333
rect 37090 9324 37096 9336
rect 37148 9324 37154 9376
rect 37918 9324 37924 9376
rect 37976 9324 37982 9376
rect 38102 9324 38108 9376
rect 38160 9364 38166 9376
rect 38657 9367 38715 9373
rect 38657 9364 38669 9367
rect 38160 9336 38669 9364
rect 38160 9324 38166 9336
rect 38657 9333 38669 9336
rect 38703 9333 38715 9367
rect 38657 9327 38715 9333
rect 39298 9324 39304 9376
rect 39356 9324 39362 9376
rect 40589 9367 40647 9373
rect 40589 9333 40601 9367
rect 40635 9364 40647 9367
rect 40862 9364 40868 9376
rect 40635 9336 40868 9364
rect 40635 9333 40647 9336
rect 40589 9327 40647 9333
rect 40862 9324 40868 9336
rect 40920 9324 40926 9376
rect 41233 9367 41291 9373
rect 41233 9333 41245 9367
rect 41279 9364 41291 9367
rect 41690 9364 41696 9376
rect 41279 9336 41696 9364
rect 41279 9333 41291 9336
rect 41233 9327 41291 9333
rect 41690 9324 41696 9336
rect 41748 9324 41754 9376
rect 41874 9324 41880 9376
rect 41932 9324 41938 9376
rect 43073 9367 43131 9373
rect 43073 9333 43085 9367
rect 43119 9364 43131 9367
rect 43254 9364 43260 9376
rect 43119 9336 43260 9364
rect 43119 9333 43131 9336
rect 43073 9327 43131 9333
rect 43254 9324 43260 9336
rect 43312 9324 43318 9376
rect 43346 9324 43352 9376
rect 43404 9364 43410 9376
rect 43809 9367 43867 9373
rect 43809 9364 43821 9367
rect 43404 9336 43821 9364
rect 43404 9324 43410 9336
rect 43809 9333 43821 9336
rect 43855 9333 43867 9367
rect 43809 9327 43867 9333
rect 43898 9324 43904 9376
rect 43956 9364 43962 9376
rect 44453 9367 44511 9373
rect 44453 9364 44465 9367
rect 43956 9336 44465 9364
rect 43956 9324 43962 9336
rect 44453 9333 44465 9336
rect 44499 9333 44511 9367
rect 44453 9327 44511 9333
rect 45554 9324 45560 9376
rect 45612 9364 45618 9376
rect 45741 9367 45799 9373
rect 45741 9364 45753 9367
rect 45612 9336 45753 9364
rect 45612 9324 45618 9336
rect 45741 9333 45753 9336
rect 45787 9333 45799 9367
rect 45741 9327 45799 9333
rect 46106 9324 46112 9376
rect 46164 9364 46170 9376
rect 46385 9367 46443 9373
rect 46385 9364 46397 9367
rect 46164 9336 46397 9364
rect 46164 9324 46170 9336
rect 46385 9333 46397 9336
rect 46431 9333 46443 9367
rect 46385 9327 46443 9333
rect 46842 9324 46848 9376
rect 46900 9364 46906 9376
rect 47029 9367 47087 9373
rect 47029 9364 47041 9367
rect 46900 9336 47041 9364
rect 46900 9324 46906 9336
rect 47029 9333 47041 9336
rect 47075 9333 47087 9367
rect 47029 9327 47087 9333
rect 47118 9324 47124 9376
rect 47176 9364 47182 9376
rect 48225 9367 48283 9373
rect 48225 9364 48237 9367
rect 47176 9336 48237 9364
rect 47176 9324 47182 9336
rect 48225 9333 48237 9336
rect 48271 9333 48283 9367
rect 48225 9327 48283 9333
rect 49234 9324 49240 9376
rect 49292 9364 49298 9376
rect 49605 9367 49663 9373
rect 49605 9364 49617 9367
rect 49292 9336 49617 9364
rect 49292 9324 49298 9336
rect 49605 9333 49617 9336
rect 49651 9333 49663 9367
rect 49605 9327 49663 9333
rect 50430 9324 50436 9376
rect 50488 9324 50494 9376
rect 51166 9324 51172 9376
rect 51224 9324 51230 9376
rect 51258 9324 51264 9376
rect 51316 9364 51322 9376
rect 51905 9367 51963 9373
rect 51905 9364 51917 9367
rect 51316 9336 51917 9364
rect 51316 9324 51322 9336
rect 51905 9333 51917 9336
rect 51951 9333 51963 9367
rect 51905 9327 51963 9333
rect 52270 9324 52276 9376
rect 52328 9364 52334 9376
rect 52825 9367 52883 9373
rect 52825 9364 52837 9367
rect 52328 9336 52837 9364
rect 52328 9324 52334 9336
rect 52825 9333 52837 9336
rect 52871 9333 52883 9367
rect 52825 9327 52883 9333
rect 53374 9324 53380 9376
rect 53432 9364 53438 9376
rect 54021 9367 54079 9373
rect 54021 9364 54033 9367
rect 53432 9336 54033 9364
rect 53432 9324 53438 9336
rect 54021 9333 54033 9336
rect 54067 9333 54079 9367
rect 54021 9327 54079 9333
rect 59630 9324 59636 9376
rect 59688 9364 59694 9376
rect 72418 9364 72424 9376
rect 59688 9336 72424 9364
rect 59688 9324 59694 9336
rect 72418 9324 72424 9336
rect 72476 9324 72482 9376
rect 74506 9364 74534 9404
rect 88242 9392 88248 9444
rect 88300 9432 88306 9444
rect 91480 9432 91508 9472
rect 92842 9460 92848 9512
rect 92900 9500 92906 9512
rect 93394 9500 93400 9512
rect 92900 9472 93400 9500
rect 92900 9460 92906 9472
rect 93394 9460 93400 9472
rect 93452 9500 93458 9512
rect 94240 9500 94268 9608
rect 94777 9571 94835 9577
rect 94777 9537 94789 9571
rect 94823 9537 94835 9571
rect 94777 9531 94835 9537
rect 95789 9571 95847 9577
rect 95789 9537 95801 9571
rect 95835 9568 95847 9571
rect 96154 9568 96160 9580
rect 95835 9540 96160 9568
rect 95835 9537 95847 9540
rect 95789 9531 95847 9537
rect 93452 9472 94268 9500
rect 94792 9500 94820 9531
rect 96154 9528 96160 9540
rect 96212 9528 96218 9580
rect 96709 9571 96767 9577
rect 96709 9537 96721 9571
rect 96755 9568 96767 9571
rect 96798 9568 96804 9580
rect 96755 9540 96804 9568
rect 96755 9537 96767 9540
rect 96709 9531 96767 9537
rect 96798 9528 96804 9540
rect 96856 9528 96862 9580
rect 97994 9528 98000 9580
rect 98052 9528 98058 9580
rect 99282 9528 99288 9580
rect 99340 9528 99346 9580
rect 99466 9528 99472 9580
rect 99524 9528 99530 9580
rect 98086 9500 98092 9512
rect 94792 9472 98092 9500
rect 93452 9460 93458 9472
rect 98086 9460 98092 9472
rect 98144 9460 98150 9512
rect 100128 9500 100156 9608
rect 100202 9528 100208 9580
rect 100260 9568 100266 9580
rect 100481 9571 100539 9577
rect 100481 9568 100493 9571
rect 100260 9540 100493 9568
rect 100260 9528 100266 9540
rect 100481 9537 100493 9540
rect 100527 9537 100539 9571
rect 100481 9531 100539 9537
rect 103238 9528 103244 9580
rect 103296 9528 103302 9580
rect 103882 9528 103888 9580
rect 103940 9528 103946 9580
rect 104894 9528 104900 9580
rect 104952 9528 104958 9580
rect 105630 9528 105636 9580
rect 105688 9528 105694 9580
rect 106274 9528 106280 9580
rect 106332 9568 106338 9580
rect 106369 9571 106427 9577
rect 106369 9568 106381 9571
rect 106332 9540 106381 9568
rect 106332 9528 106338 9540
rect 106369 9537 106381 9540
rect 106415 9537 106427 9571
rect 106369 9531 106427 9537
rect 107746 9528 107752 9580
rect 107804 9528 107810 9580
rect 108390 9528 108396 9580
rect 108448 9528 108454 9580
rect 109034 9528 109040 9580
rect 109092 9528 109098 9580
rect 110046 9528 110052 9580
rect 110104 9528 110110 9580
rect 110782 9528 110788 9580
rect 110840 9528 110846 9580
rect 111518 9528 111524 9580
rect 111576 9528 111582 9580
rect 112898 9528 112904 9580
rect 112956 9528 112962 9580
rect 113542 9528 113548 9580
rect 113600 9528 113606 9580
rect 114186 9528 114192 9580
rect 114244 9528 114250 9580
rect 115198 9528 115204 9580
rect 115256 9528 115262 9580
rect 115934 9528 115940 9580
rect 115992 9528 115998 9580
rect 116670 9528 116676 9580
rect 116728 9528 116734 9580
rect 118050 9528 118056 9580
rect 118108 9528 118114 9580
rect 118694 9528 118700 9580
rect 118752 9528 118758 9580
rect 119338 9528 119344 9580
rect 119396 9528 119402 9580
rect 120350 9528 120356 9580
rect 120408 9528 120414 9580
rect 121086 9528 121092 9580
rect 121144 9528 121150 9580
rect 121733 9571 121791 9577
rect 121733 9537 121745 9571
rect 121779 9537 121791 9571
rect 121733 9531 121791 9537
rect 121270 9500 121276 9512
rect 100128 9472 121276 9500
rect 121270 9460 121276 9472
rect 121328 9460 121334 9512
rect 121454 9460 121460 9512
rect 121512 9500 121518 9512
rect 121748 9500 121776 9531
rect 121512 9472 121960 9500
rect 121512 9460 121518 9472
rect 111702 9432 111708 9444
rect 88300 9404 89714 9432
rect 91480 9404 111708 9432
rect 88300 9392 88306 9404
rect 87782 9364 87788 9376
rect 74506 9336 87788 9364
rect 87782 9324 87788 9336
rect 87840 9324 87846 9376
rect 88794 9324 88800 9376
rect 88852 9364 88858 9376
rect 89441 9367 89499 9373
rect 89441 9364 89453 9367
rect 88852 9336 89453 9364
rect 88852 9324 88858 9336
rect 89441 9333 89453 9336
rect 89487 9333 89499 9367
rect 89686 9364 89714 9404
rect 111702 9392 111708 9404
rect 111760 9392 111766 9444
rect 111886 9392 111892 9444
rect 111944 9432 111950 9444
rect 114005 9435 114063 9441
rect 114005 9432 114017 9435
rect 111944 9404 114017 9432
rect 111944 9392 111950 9404
rect 114005 9401 114017 9404
rect 114051 9401 114063 9435
rect 114005 9395 114063 9401
rect 114278 9392 114284 9444
rect 114336 9432 114342 9444
rect 114336 9404 115152 9432
rect 114336 9392 114342 9404
rect 92198 9364 92204 9376
rect 89686 9336 92204 9364
rect 89441 9327 89499 9333
rect 92198 9324 92204 9336
rect 92256 9364 92262 9376
rect 93210 9364 93216 9376
rect 92256 9336 93216 9364
rect 92256 9324 92262 9336
rect 93210 9324 93216 9336
rect 93268 9324 93274 9376
rect 94314 9324 94320 9376
rect 94372 9364 94378 9376
rect 94869 9367 94927 9373
rect 94869 9364 94881 9367
rect 94372 9336 94881 9364
rect 94372 9324 94378 9336
rect 94869 9333 94881 9336
rect 94915 9333 94927 9367
rect 94869 9327 94927 9333
rect 94958 9324 94964 9376
rect 95016 9364 95022 9376
rect 98270 9364 98276 9376
rect 95016 9336 98276 9364
rect 95016 9324 95022 9336
rect 98270 9324 98276 9336
rect 98328 9324 98334 9376
rect 99374 9324 99380 9376
rect 99432 9364 99438 9376
rect 99653 9367 99711 9373
rect 99653 9364 99665 9367
rect 99432 9336 99665 9364
rect 99432 9324 99438 9336
rect 99653 9333 99665 9336
rect 99699 9333 99711 9367
rect 99653 9327 99711 9333
rect 100386 9324 100392 9376
rect 100444 9364 100450 9376
rect 106185 9367 106243 9373
rect 106185 9364 106197 9367
rect 100444 9336 106197 9364
rect 100444 9324 100450 9336
rect 106185 9333 106197 9336
rect 106231 9333 106243 9367
rect 106185 9327 106243 9333
rect 107562 9324 107568 9376
rect 107620 9324 107626 9376
rect 108206 9324 108212 9376
rect 108264 9324 108270 9376
rect 109862 9324 109868 9376
rect 109920 9324 109926 9376
rect 110598 9324 110604 9376
rect 110656 9324 110662 9376
rect 112714 9324 112720 9376
rect 112772 9324 112778 9376
rect 113358 9324 113364 9376
rect 113416 9324 113422 9376
rect 115014 9324 115020 9376
rect 115072 9324 115078 9376
rect 115124 9364 115152 9404
rect 115658 9392 115664 9444
rect 115716 9432 115722 9444
rect 117869 9435 117927 9441
rect 117869 9432 117881 9435
rect 115716 9404 117881 9432
rect 115716 9392 115722 9404
rect 117869 9401 117881 9404
rect 117915 9401 117927 9435
rect 117869 9395 117927 9401
rect 115753 9367 115811 9373
rect 115753 9364 115765 9367
rect 115124 9336 115765 9364
rect 115753 9333 115765 9336
rect 115799 9333 115811 9367
rect 115753 9327 115811 9333
rect 115842 9324 115848 9376
rect 115900 9364 115906 9376
rect 116489 9367 116547 9373
rect 116489 9364 116501 9367
rect 115900 9336 116501 9364
rect 115900 9324 115906 9336
rect 116489 9333 116501 9336
rect 116535 9333 116547 9367
rect 116489 9327 116547 9333
rect 118326 9324 118332 9376
rect 118384 9364 118390 9376
rect 118513 9367 118571 9373
rect 118513 9364 118525 9367
rect 118384 9336 118525 9364
rect 118384 9324 118390 9336
rect 118513 9333 118525 9336
rect 118559 9333 118571 9367
rect 118513 9327 118571 9333
rect 119154 9324 119160 9376
rect 119212 9324 119218 9376
rect 120166 9324 120172 9376
rect 120224 9324 120230 9376
rect 120905 9367 120963 9373
rect 120905 9333 120917 9367
rect 120951 9364 120963 9367
rect 120994 9364 121000 9376
rect 120951 9336 121000 9364
rect 120951 9333 120963 9336
rect 120905 9327 120963 9333
rect 120994 9324 121000 9336
rect 121052 9324 121058 9376
rect 121730 9324 121736 9376
rect 121788 9364 121794 9376
rect 121825 9367 121883 9373
rect 121825 9364 121837 9367
rect 121788 9336 121837 9364
rect 121788 9324 121794 9336
rect 121825 9333 121837 9336
rect 121871 9333 121883 9367
rect 121932 9364 121960 9472
rect 122392 9432 122420 9608
rect 122466 9528 122472 9580
rect 122524 9528 122530 9580
rect 122576 9500 122604 9676
rect 122650 9664 122656 9716
rect 122708 9664 122714 9716
rect 125226 9664 125232 9716
rect 125284 9664 125290 9716
rect 127894 9664 127900 9716
rect 127952 9664 127958 9716
rect 128814 9664 128820 9716
rect 128872 9664 128878 9716
rect 129553 9707 129611 9713
rect 129553 9673 129565 9707
rect 129599 9704 129611 9707
rect 129642 9704 129648 9716
rect 129599 9676 129648 9704
rect 129599 9673 129611 9676
rect 129553 9667 129611 9673
rect 129642 9664 129648 9676
rect 129700 9664 129706 9716
rect 131482 9664 131488 9716
rect 131540 9664 131546 9716
rect 133506 9664 133512 9716
rect 133564 9664 133570 9716
rect 134242 9664 134248 9716
rect 134300 9664 134306 9716
rect 137278 9664 137284 9716
rect 137336 9704 137342 9716
rect 152458 9704 152464 9716
rect 137336 9676 152464 9704
rect 137336 9664 137342 9676
rect 152458 9664 152464 9676
rect 152516 9664 152522 9716
rect 153381 9707 153439 9713
rect 153381 9673 153393 9707
rect 153427 9704 153439 9707
rect 155862 9704 155868 9716
rect 153427 9676 155868 9704
rect 153427 9673 153439 9676
rect 153381 9667 153439 9673
rect 155862 9664 155868 9676
rect 155920 9664 155926 9716
rect 155954 9664 155960 9716
rect 156012 9704 156018 9716
rect 156141 9707 156199 9713
rect 156141 9704 156153 9707
rect 156012 9676 156153 9704
rect 156012 9664 156018 9676
rect 156141 9673 156153 9676
rect 156187 9673 156199 9707
rect 156141 9667 156199 9673
rect 156874 9664 156880 9716
rect 156932 9664 156938 9716
rect 157242 9664 157248 9716
rect 157300 9704 157306 9716
rect 157613 9707 157671 9713
rect 157613 9704 157625 9707
rect 157300 9676 157625 9704
rect 157300 9664 157306 9676
rect 157613 9673 157625 9676
rect 157659 9673 157671 9707
rect 157613 9667 157671 9673
rect 157978 9664 157984 9716
rect 158036 9704 158042 9716
rect 158717 9707 158775 9713
rect 158717 9704 158729 9707
rect 158036 9676 158729 9704
rect 158036 9664 158042 9676
rect 158717 9673 158729 9676
rect 158763 9673 158775 9707
rect 158717 9667 158775 9673
rect 159450 9664 159456 9716
rect 159508 9704 159514 9716
rect 160189 9707 160247 9713
rect 160189 9704 160201 9707
rect 159508 9676 160201 9704
rect 159508 9664 159514 9676
rect 160189 9673 160201 9676
rect 160235 9673 160247 9707
rect 160189 9667 160247 9673
rect 161937 9707 161995 9713
rect 161937 9673 161949 9707
rect 161983 9704 161995 9707
rect 162302 9704 162308 9716
rect 161983 9676 162308 9704
rect 161983 9673 161995 9676
rect 161937 9667 161995 9673
rect 162302 9664 162308 9676
rect 162360 9664 162366 9716
rect 163866 9664 163872 9716
rect 163924 9704 163930 9716
rect 165617 9707 165675 9713
rect 165617 9704 165629 9707
rect 163924 9676 165629 9704
rect 163924 9664 163930 9676
rect 165617 9673 165629 9676
rect 165663 9673 165675 9707
rect 165617 9667 165675 9673
rect 165724 9676 179460 9704
rect 130565 9639 130623 9645
rect 130565 9636 130577 9639
rect 129384 9608 130577 9636
rect 124582 9528 124588 9580
rect 124640 9568 124646 9580
rect 125045 9571 125103 9577
rect 125045 9568 125057 9571
rect 124640 9540 125057 9568
rect 124640 9528 124646 9540
rect 125045 9537 125057 9540
rect 125091 9537 125103 9571
rect 125045 9531 125103 9537
rect 127713 9571 127771 9577
rect 127713 9537 127725 9571
rect 127759 9568 127771 9571
rect 127986 9568 127992 9580
rect 127759 9540 127992 9568
rect 127759 9537 127771 9540
rect 127713 9531 127771 9537
rect 127986 9528 127992 9540
rect 128044 9528 128050 9580
rect 128630 9528 128636 9580
rect 128688 9528 128694 9580
rect 129384 9577 129412 9608
rect 130565 9605 130577 9608
rect 130611 9605 130623 9639
rect 130565 9599 130623 9605
rect 146386 9596 146392 9648
rect 146444 9636 146450 9648
rect 146444 9608 162072 9636
rect 146444 9596 146450 9608
rect 129369 9571 129427 9577
rect 129369 9537 129381 9571
rect 129415 9537 129427 9571
rect 129369 9531 129427 9537
rect 129458 9528 129464 9580
rect 129516 9568 129522 9580
rect 130197 9571 130255 9577
rect 130197 9568 130209 9571
rect 129516 9540 130209 9568
rect 129516 9528 129522 9540
rect 130197 9537 130209 9540
rect 130243 9537 130255 9571
rect 130197 9531 130255 9537
rect 125870 9500 125876 9512
rect 122576 9472 125876 9500
rect 125870 9460 125876 9472
rect 125928 9460 125934 9512
rect 130212 9500 130240 9531
rect 130378 9528 130384 9580
rect 130436 9528 130442 9580
rect 131301 9571 131359 9577
rect 131301 9537 131313 9571
rect 131347 9568 131359 9571
rect 131390 9568 131396 9580
rect 131347 9540 131396 9568
rect 131347 9537 131359 9540
rect 131301 9531 131359 9537
rect 131390 9528 131396 9540
rect 131448 9528 131454 9580
rect 133325 9571 133383 9577
rect 133325 9537 133337 9571
rect 133371 9568 133383 9571
rect 133414 9568 133420 9580
rect 133371 9540 133420 9568
rect 133371 9537 133383 9540
rect 133325 9531 133383 9537
rect 133414 9528 133420 9540
rect 133472 9528 133478 9580
rect 134061 9571 134119 9577
rect 134061 9537 134073 9571
rect 134107 9568 134119 9571
rect 134242 9568 134248 9580
rect 134107 9540 134248 9568
rect 134107 9537 134119 9540
rect 134061 9531 134119 9537
rect 134242 9528 134248 9540
rect 134300 9528 134306 9580
rect 137370 9528 137376 9580
rect 137428 9568 137434 9580
rect 138109 9571 138167 9577
rect 138109 9568 138121 9571
rect 137428 9540 138121 9568
rect 137428 9528 137434 9540
rect 138109 9537 138121 9540
rect 138155 9537 138167 9571
rect 138109 9531 138167 9537
rect 138750 9528 138756 9580
rect 138808 9528 138814 9580
rect 138842 9528 138848 9580
rect 138900 9568 138906 9580
rect 139397 9571 139455 9577
rect 139397 9568 139409 9571
rect 138900 9540 139409 9568
rect 138900 9528 138906 9540
rect 139397 9537 139409 9540
rect 139443 9537 139455 9571
rect 139397 9531 139455 9537
rect 140682 9528 140688 9580
rect 140740 9528 140746 9580
rect 141326 9528 141332 9580
rect 141384 9528 141390 9580
rect 141970 9528 141976 9580
rect 142028 9528 142034 9580
rect 143258 9528 143264 9580
rect 143316 9528 143322 9580
rect 143350 9528 143356 9580
rect 143408 9568 143414 9580
rect 143905 9571 143963 9577
rect 143905 9568 143917 9571
rect 143408 9540 143917 9568
rect 143408 9528 143414 9540
rect 143905 9537 143917 9540
rect 143951 9537 143963 9571
rect 143905 9531 143963 9537
rect 144546 9528 144552 9580
rect 144604 9528 144610 9580
rect 145834 9528 145840 9580
rect 145892 9528 145898 9580
rect 146202 9528 146208 9580
rect 146260 9568 146266 9580
rect 146481 9571 146539 9577
rect 146481 9568 146493 9571
rect 146260 9540 146493 9568
rect 146260 9528 146266 9540
rect 146481 9537 146493 9540
rect 146527 9537 146539 9571
rect 146481 9531 146539 9537
rect 147122 9528 147128 9580
rect 147180 9528 147186 9580
rect 148410 9528 148416 9580
rect 148468 9528 148474 9580
rect 148502 9528 148508 9580
rect 148560 9568 148566 9580
rect 149057 9571 149115 9577
rect 149057 9568 149069 9571
rect 148560 9540 149069 9568
rect 148560 9528 148566 9540
rect 149057 9537 149069 9540
rect 149103 9537 149115 9571
rect 149057 9531 149115 9537
rect 149698 9528 149704 9580
rect 149756 9528 149762 9580
rect 150986 9528 150992 9580
rect 151044 9528 151050 9580
rect 151630 9528 151636 9580
rect 151688 9528 151694 9580
rect 152274 9528 152280 9580
rect 152332 9528 152338 9580
rect 153194 9528 153200 9580
rect 153252 9568 153258 9580
rect 153565 9571 153623 9577
rect 153565 9568 153577 9571
rect 153252 9540 153577 9568
rect 153252 9528 153258 9540
rect 153565 9537 153577 9540
rect 153611 9537 153623 9571
rect 153565 9531 153623 9537
rect 154206 9528 154212 9580
rect 154264 9528 154270 9580
rect 154574 9528 154580 9580
rect 154632 9568 154638 9580
rect 154853 9571 154911 9577
rect 154853 9568 154865 9571
rect 154632 9540 154865 9568
rect 154632 9528 154638 9540
rect 154853 9537 154865 9540
rect 154899 9537 154911 9571
rect 154853 9531 154911 9537
rect 155512 9540 155724 9568
rect 152366 9500 152372 9512
rect 130212 9472 152372 9500
rect 152366 9460 152372 9472
rect 152424 9460 152430 9512
rect 155512 9500 155540 9540
rect 154040 9472 155540 9500
rect 129090 9432 129096 9444
rect 122392 9404 129096 9432
rect 129090 9392 129096 9404
rect 129148 9432 129154 9444
rect 138569 9435 138627 9441
rect 138569 9432 138581 9435
rect 129148 9404 132494 9432
rect 129148 9392 129154 9404
rect 129274 9364 129280 9376
rect 121932 9336 129280 9364
rect 121825 9327 121883 9333
rect 129274 9324 129280 9336
rect 129332 9324 129338 9376
rect 132466 9364 132494 9404
rect 137986 9404 138581 9432
rect 137278 9364 137284 9376
rect 132466 9336 137284 9364
rect 137278 9324 137284 9336
rect 137336 9324 137342 9376
rect 137738 9324 137744 9376
rect 137796 9364 137802 9376
rect 137986 9364 138014 9404
rect 138569 9401 138581 9404
rect 138615 9401 138627 9435
rect 138569 9395 138627 9401
rect 141145 9435 141203 9441
rect 141145 9401 141157 9435
rect 141191 9432 141203 9435
rect 142706 9432 142712 9444
rect 141191 9404 142712 9432
rect 141191 9401 141203 9404
rect 141145 9395 141203 9401
rect 142706 9392 142712 9404
rect 142764 9392 142770 9444
rect 143721 9435 143779 9441
rect 143721 9401 143733 9435
rect 143767 9432 143779 9435
rect 145374 9432 145380 9444
rect 143767 9404 145380 9432
rect 143767 9401 143779 9404
rect 143721 9395 143779 9401
rect 145374 9392 145380 9404
rect 145432 9392 145438 9444
rect 145834 9392 145840 9444
rect 145892 9432 145898 9444
rect 146941 9435 146999 9441
rect 146941 9432 146953 9435
rect 145892 9404 146953 9432
rect 145892 9392 145898 9404
rect 146941 9401 146953 9404
rect 146987 9401 146999 9435
rect 146941 9395 146999 9401
rect 148873 9435 148931 9441
rect 148873 9401 148885 9435
rect 148919 9432 148931 9435
rect 150526 9432 150532 9444
rect 148919 9404 150532 9432
rect 148919 9401 148931 9404
rect 148873 9395 148931 9401
rect 150526 9392 150532 9404
rect 150584 9392 150590 9444
rect 154040 9441 154068 9472
rect 154025 9435 154083 9441
rect 154025 9401 154037 9435
rect 154071 9401 154083 9435
rect 154025 9395 154083 9401
rect 137796 9336 138014 9364
rect 137796 9324 137802 9336
rect 138106 9324 138112 9376
rect 138164 9364 138170 9376
rect 139213 9367 139271 9373
rect 139213 9364 139225 9367
rect 138164 9336 139225 9364
rect 138164 9324 138170 9336
rect 139213 9333 139225 9336
rect 139259 9333 139271 9367
rect 139213 9327 139271 9333
rect 140498 9324 140504 9376
rect 140556 9324 140562 9376
rect 141789 9367 141847 9373
rect 141789 9333 141801 9367
rect 141835 9364 141847 9367
rect 142982 9364 142988 9376
rect 141835 9336 142988 9364
rect 141835 9333 141847 9336
rect 141789 9327 141847 9333
rect 142982 9324 142988 9336
rect 143040 9324 143046 9376
rect 143077 9367 143135 9373
rect 143077 9333 143089 9367
rect 143123 9364 143135 9367
rect 143258 9364 143264 9376
rect 143123 9336 143264 9364
rect 143123 9333 143135 9336
rect 143077 9327 143135 9333
rect 143258 9324 143264 9336
rect 143316 9324 143322 9376
rect 144365 9367 144423 9373
rect 144365 9333 144377 9367
rect 144411 9364 144423 9367
rect 145558 9364 145564 9376
rect 144411 9336 145564 9364
rect 144411 9333 144423 9336
rect 144365 9327 144423 9333
rect 145558 9324 145564 9336
rect 145616 9324 145622 9376
rect 145653 9367 145711 9373
rect 145653 9333 145665 9367
rect 145699 9364 145711 9367
rect 146202 9364 146208 9376
rect 145699 9336 146208 9364
rect 145699 9333 145711 9336
rect 145653 9327 145711 9333
rect 146202 9324 146208 9336
rect 146260 9324 146266 9376
rect 146294 9324 146300 9376
rect 146352 9324 146358 9376
rect 148226 9324 148232 9376
rect 148284 9324 148290 9376
rect 149517 9367 149575 9373
rect 149517 9333 149529 9367
rect 149563 9364 149575 9367
rect 150434 9364 150440 9376
rect 149563 9336 150440 9364
rect 149563 9333 149575 9336
rect 149517 9327 149575 9333
rect 150434 9324 150440 9336
rect 150492 9324 150498 9376
rect 150805 9367 150863 9373
rect 150805 9333 150817 9367
rect 150851 9364 150863 9367
rect 151262 9364 151268 9376
rect 150851 9336 151268 9364
rect 150851 9333 150863 9336
rect 150805 9327 150863 9333
rect 151262 9324 151268 9336
rect 151320 9324 151326 9376
rect 151449 9367 151507 9373
rect 151449 9333 151461 9367
rect 151495 9364 151507 9367
rect 151906 9364 151912 9376
rect 151495 9336 151912 9364
rect 151495 9333 151507 9336
rect 151449 9327 151507 9333
rect 151906 9324 151912 9336
rect 151964 9324 151970 9376
rect 152093 9367 152151 9373
rect 152093 9333 152105 9367
rect 152139 9364 152151 9367
rect 154574 9364 154580 9376
rect 152139 9336 154580 9364
rect 152139 9333 152151 9336
rect 152093 9327 152151 9333
rect 154574 9324 154580 9336
rect 154632 9324 154638 9376
rect 154669 9367 154727 9373
rect 154669 9333 154681 9367
rect 154715 9364 154727 9367
rect 155586 9364 155592 9376
rect 154715 9336 155592 9364
rect 154715 9333 154727 9336
rect 154669 9327 154727 9333
rect 155586 9324 155592 9336
rect 155644 9324 155650 9376
rect 155696 9364 155724 9540
rect 155770 9528 155776 9580
rect 155828 9528 155834 9580
rect 155957 9571 156015 9577
rect 155957 9537 155969 9571
rect 156003 9568 156015 9571
rect 156138 9568 156144 9580
rect 156003 9540 156144 9568
rect 156003 9537 156015 9540
rect 155957 9531 156015 9537
rect 156138 9528 156144 9540
rect 156196 9528 156202 9580
rect 156693 9571 156751 9577
rect 156693 9537 156705 9571
rect 156739 9568 156751 9571
rect 156966 9568 156972 9580
rect 156739 9540 156972 9568
rect 156739 9537 156751 9540
rect 156693 9531 156751 9537
rect 156966 9528 156972 9540
rect 157024 9528 157030 9580
rect 157426 9528 157432 9580
rect 157484 9528 157490 9580
rect 157794 9528 157800 9580
rect 157852 9568 157858 9580
rect 158533 9571 158591 9577
rect 158533 9568 158545 9571
rect 157852 9540 158545 9568
rect 157852 9528 157858 9540
rect 158533 9537 158545 9540
rect 158579 9537 158591 9571
rect 158533 9531 158591 9537
rect 159266 9528 159272 9580
rect 159324 9528 159330 9580
rect 159358 9528 159364 9580
rect 159416 9568 159422 9580
rect 160005 9571 160063 9577
rect 160005 9568 160017 9571
rect 159416 9540 160017 9568
rect 159416 9528 159422 9540
rect 160005 9537 160017 9540
rect 160051 9537 160063 9571
rect 160005 9531 160063 9537
rect 161293 9571 161351 9577
rect 161293 9537 161305 9571
rect 161339 9568 161351 9571
rect 161658 9568 161664 9580
rect 161339 9540 161664 9568
rect 161339 9537 161351 9540
rect 161293 9531 161351 9537
rect 161658 9528 161664 9540
rect 161716 9528 161722 9580
rect 155788 9500 155816 9528
rect 157978 9500 157984 9512
rect 155788 9472 157984 9500
rect 157978 9460 157984 9472
rect 158036 9460 158042 9512
rect 159376 9472 159588 9500
rect 155770 9392 155776 9444
rect 155828 9432 155834 9444
rect 159376 9432 159404 9472
rect 155828 9404 159404 9432
rect 155828 9392 155834 9404
rect 159450 9392 159456 9444
rect 159508 9392 159514 9444
rect 159560 9432 159588 9472
rect 160922 9460 160928 9512
rect 160980 9500 160986 9512
rect 161109 9503 161167 9509
rect 161109 9500 161121 9503
rect 160980 9472 161121 9500
rect 160980 9460 160986 9472
rect 161109 9469 161121 9472
rect 161155 9469 161167 9503
rect 161109 9463 161167 9469
rect 161750 9432 161756 9444
rect 159560 9404 161756 9432
rect 161750 9392 161756 9404
rect 161808 9392 161814 9444
rect 162044 9432 162072 9608
rect 162394 9596 162400 9648
rect 162452 9636 162458 9648
rect 165724 9636 165752 9676
rect 162452 9608 165752 9636
rect 162452 9596 162458 9608
rect 165798 9596 165804 9648
rect 165856 9636 165862 9648
rect 170582 9636 170588 9648
rect 165856 9608 170588 9636
rect 165856 9596 165862 9608
rect 170582 9596 170588 9608
rect 170640 9596 170646 9648
rect 172330 9596 172336 9648
rect 172388 9596 172394 9648
rect 172514 9596 172520 9648
rect 172572 9596 172578 9648
rect 173066 9596 173072 9648
rect 173124 9596 173130 9648
rect 175182 9596 175188 9648
rect 175240 9636 175246 9648
rect 175829 9639 175887 9645
rect 175829 9636 175841 9639
rect 175240 9608 175841 9636
rect 175240 9596 175246 9608
rect 175829 9605 175841 9608
rect 175875 9605 175887 9639
rect 175829 9599 175887 9605
rect 175918 9596 175924 9648
rect 175976 9636 175982 9648
rect 176657 9639 176715 9645
rect 176657 9636 176669 9639
rect 175976 9608 176669 9636
rect 175976 9596 175982 9608
rect 176657 9605 176669 9608
rect 176703 9605 176715 9639
rect 176657 9599 176715 9605
rect 162302 9528 162308 9580
rect 162360 9528 162366 9580
rect 163961 9571 164019 9577
rect 163961 9537 163973 9571
rect 164007 9568 164019 9571
rect 164326 9568 164332 9580
rect 164007 9540 164332 9568
rect 164007 9537 164019 9540
rect 163961 9531 164019 9537
rect 164326 9528 164332 9540
rect 164384 9528 164390 9580
rect 165154 9528 165160 9580
rect 165212 9568 165218 9580
rect 165433 9571 165491 9577
rect 165433 9568 165445 9571
rect 165212 9540 165445 9568
rect 165212 9528 165218 9540
rect 165433 9537 165445 9540
rect 165479 9537 165491 9571
rect 165433 9531 165491 9537
rect 165522 9528 165528 9580
rect 165580 9568 165586 9580
rect 166445 9571 166503 9577
rect 166445 9568 166457 9571
rect 165580 9540 166457 9568
rect 165580 9528 165586 9540
rect 166445 9537 166457 9540
rect 166491 9568 166503 9571
rect 167273 9571 167331 9577
rect 167273 9568 167285 9571
rect 166491 9540 167285 9568
rect 166491 9537 166503 9540
rect 166445 9531 166503 9537
rect 167273 9537 167285 9540
rect 167319 9568 167331 9571
rect 168098 9568 168104 9580
rect 167319 9540 168104 9568
rect 167319 9537 167331 9540
rect 167273 9531 167331 9537
rect 168098 9528 168104 9540
rect 168156 9568 168162 9580
rect 168156 9540 169248 9568
rect 168156 9528 168162 9540
rect 162762 9460 162768 9512
rect 162820 9460 162826 9512
rect 164602 9460 164608 9512
rect 164660 9460 164666 9512
rect 166258 9460 166264 9512
rect 166316 9460 166322 9512
rect 167086 9460 167092 9512
rect 167144 9460 167150 9512
rect 167546 9460 167552 9512
rect 167604 9500 167610 9512
rect 167914 9500 167920 9512
rect 167604 9472 167920 9500
rect 167604 9460 167610 9472
rect 167914 9460 167920 9472
rect 167972 9500 167978 9512
rect 168282 9500 168288 9512
rect 167972 9472 168288 9500
rect 167972 9460 167978 9472
rect 168282 9460 168288 9472
rect 168340 9460 168346 9512
rect 169110 9460 169116 9512
rect 169168 9460 169174 9512
rect 169220 9500 169248 9540
rect 169294 9528 169300 9580
rect 169352 9568 169358 9580
rect 169352 9540 171134 9568
rect 169352 9528 169358 9540
rect 169389 9503 169447 9509
rect 169389 9500 169401 9503
rect 169220 9472 169401 9500
rect 169389 9469 169401 9472
rect 169435 9500 169447 9503
rect 169754 9500 169760 9512
rect 169435 9472 169760 9500
rect 169435 9469 169447 9472
rect 169389 9463 169447 9469
rect 169754 9460 169760 9472
rect 169812 9460 169818 9512
rect 171106 9500 171134 9540
rect 171686 9528 171692 9580
rect 171744 9528 171750 9580
rect 174446 9528 174452 9580
rect 174504 9528 174510 9580
rect 177761 9571 177819 9577
rect 174648 9540 177712 9568
rect 174648 9500 174676 9540
rect 171106 9472 174676 9500
rect 174722 9460 174728 9512
rect 174780 9460 174786 9512
rect 176841 9435 176899 9441
rect 176841 9432 176853 9435
rect 162044 9404 176853 9432
rect 176841 9401 176853 9404
rect 176887 9401 176899 9435
rect 177684 9432 177712 9540
rect 177761 9537 177773 9571
rect 177807 9568 177819 9571
rect 177942 9568 177948 9580
rect 177807 9540 177948 9568
rect 177807 9537 177819 9540
rect 177761 9531 177819 9537
rect 177942 9528 177948 9540
rect 178000 9528 178006 9580
rect 179138 9528 179144 9580
rect 179196 9528 179202 9580
rect 179432 9577 179460 9676
rect 179966 9664 179972 9716
rect 180024 9704 180030 9716
rect 180024 9676 192524 9704
rect 180024 9664 180030 9676
rect 179417 9571 179475 9577
rect 179417 9537 179429 9571
rect 179463 9537 179475 9571
rect 179417 9531 179475 9537
rect 181714 9528 181720 9580
rect 181772 9528 181778 9580
rect 181990 9528 181996 9580
rect 182048 9528 182054 9580
rect 182542 9528 182548 9580
rect 182600 9568 182606 9580
rect 184293 9571 184351 9577
rect 184293 9568 184305 9571
rect 182600 9540 184305 9568
rect 182600 9528 182606 9540
rect 184293 9537 184305 9540
rect 184339 9537 184351 9571
rect 184293 9531 184351 9537
rect 185486 9528 185492 9580
rect 185544 9568 185550 9580
rect 186869 9571 186927 9577
rect 186869 9568 186881 9571
rect 185544 9540 186881 9568
rect 185544 9528 185550 9540
rect 186869 9537 186881 9540
rect 186915 9537 186927 9571
rect 186869 9531 186927 9537
rect 187694 9528 187700 9580
rect 187752 9568 187758 9580
rect 189445 9571 189503 9577
rect 189445 9568 189457 9571
rect 187752 9540 189457 9568
rect 187752 9528 187758 9540
rect 189445 9537 189457 9540
rect 189491 9537 189503 9571
rect 189445 9531 189503 9537
rect 189994 9528 190000 9580
rect 190052 9568 190058 9580
rect 190822 9568 190828 9580
rect 190052 9540 190828 9568
rect 190052 9528 190058 9540
rect 190822 9528 190828 9540
rect 190880 9528 190886 9580
rect 192386 9528 192392 9580
rect 192444 9528 192450 9580
rect 178034 9460 178040 9512
rect 178092 9460 178098 9512
rect 184566 9460 184572 9512
rect 184624 9460 184630 9512
rect 187145 9503 187203 9509
rect 187145 9469 187157 9503
rect 187191 9469 187203 9503
rect 187145 9463 187203 9469
rect 185946 9432 185952 9444
rect 177684 9404 185952 9432
rect 176841 9395 176899 9401
rect 185946 9392 185952 9404
rect 186004 9392 186010 9444
rect 157702 9364 157708 9376
rect 155696 9336 157708 9364
rect 157702 9324 157708 9336
rect 157760 9324 157766 9376
rect 161106 9324 161112 9376
rect 161164 9364 161170 9376
rect 161477 9367 161535 9373
rect 161477 9364 161489 9367
rect 161164 9336 161489 9364
rect 161164 9324 161170 9336
rect 161477 9333 161489 9336
rect 161523 9333 161535 9367
rect 161477 9327 161535 9333
rect 161842 9324 161848 9376
rect 161900 9364 161906 9376
rect 165798 9364 165804 9376
rect 161900 9336 165804 9364
rect 161900 9324 161906 9336
rect 165798 9324 165804 9336
rect 165856 9324 165862 9376
rect 166166 9324 166172 9376
rect 166224 9364 166230 9376
rect 166629 9367 166687 9373
rect 166629 9364 166641 9367
rect 166224 9336 166641 9364
rect 166224 9324 166230 9336
rect 166629 9333 166641 9336
rect 166675 9333 166687 9367
rect 166629 9327 166687 9333
rect 167454 9324 167460 9376
rect 167512 9324 167518 9376
rect 168285 9367 168343 9373
rect 168285 9333 168297 9367
rect 168331 9364 168343 9367
rect 168834 9364 168840 9376
rect 168331 9336 168840 9364
rect 168331 9333 168343 9336
rect 168285 9327 168343 9333
rect 168834 9324 168840 9336
rect 168892 9324 168898 9376
rect 173158 9324 173164 9376
rect 173216 9324 173222 9376
rect 175918 9324 175924 9376
rect 175976 9324 175982 9376
rect 177942 9324 177948 9376
rect 178000 9364 178006 9376
rect 187160 9364 187188 9463
rect 189718 9460 189724 9512
rect 189776 9460 189782 9512
rect 192496 9500 192524 9676
rect 192570 9664 192576 9716
rect 192628 9664 192634 9716
rect 192846 9664 192852 9716
rect 192904 9704 192910 9716
rect 193401 9707 193459 9713
rect 193401 9704 193413 9707
rect 192904 9676 193413 9704
rect 192904 9664 192910 9676
rect 193401 9673 193413 9676
rect 193447 9673 193459 9707
rect 193401 9667 193459 9673
rect 194318 9664 194324 9716
rect 194376 9704 194382 9716
rect 194873 9707 194931 9713
rect 194873 9704 194885 9707
rect 194376 9676 194885 9704
rect 194376 9664 194382 9676
rect 194873 9673 194885 9676
rect 194919 9673 194931 9707
rect 194873 9667 194931 9673
rect 195790 9664 195796 9716
rect 195848 9704 195854 9716
rect 196345 9707 196403 9713
rect 196345 9704 196357 9707
rect 195848 9676 196357 9704
rect 195848 9664 195854 9676
rect 196345 9673 196357 9676
rect 196391 9673 196403 9707
rect 196345 9667 196403 9673
rect 196526 9664 196532 9716
rect 196584 9704 196590 9716
rect 197357 9707 197415 9713
rect 197357 9704 197369 9707
rect 196584 9676 197369 9704
rect 196584 9664 196590 9676
rect 197357 9673 197369 9676
rect 197403 9673 197415 9707
rect 197357 9667 197415 9673
rect 197998 9664 198004 9716
rect 198056 9704 198062 9716
rect 198829 9707 198887 9713
rect 198829 9704 198841 9707
rect 198056 9676 198841 9704
rect 198056 9664 198062 9676
rect 198829 9673 198841 9676
rect 198875 9673 198887 9707
rect 198829 9667 198887 9673
rect 200022 9664 200028 9716
rect 200080 9664 200086 9716
rect 200114 9664 200120 9716
rect 200172 9704 200178 9716
rect 200172 9676 200896 9704
rect 200172 9664 200178 9676
rect 200868 9636 200896 9676
rect 202506 9664 202512 9716
rect 202564 9664 202570 9716
rect 202598 9664 202604 9716
rect 202656 9704 202662 9716
rect 203245 9707 203303 9713
rect 203245 9704 203257 9707
rect 202656 9676 203257 9704
rect 202656 9664 202662 9676
rect 203245 9673 203257 9676
rect 203291 9673 203303 9707
rect 203245 9667 203303 9673
rect 207477 9707 207535 9713
rect 207477 9673 207489 9707
rect 207523 9704 207535 9707
rect 209590 9704 209596 9716
rect 207523 9676 209596 9704
rect 207523 9673 207535 9676
rect 207477 9667 207535 9673
rect 209590 9664 209596 9676
rect 209648 9664 209654 9716
rect 212534 9704 212540 9716
rect 209746 9676 212540 9704
rect 209746 9636 209774 9676
rect 212534 9664 212540 9676
rect 212592 9664 212598 9716
rect 212629 9707 212687 9713
rect 212629 9673 212641 9707
rect 212675 9673 212687 9707
rect 212629 9667 212687 9673
rect 200868 9608 209774 9636
rect 210786 9596 210792 9648
rect 210844 9636 210850 9648
rect 212644 9636 212672 9667
rect 212718 9664 212724 9716
rect 212776 9704 212782 9716
rect 224310 9704 224316 9716
rect 212776 9676 224316 9704
rect 212776 9664 212782 9676
rect 224310 9664 224316 9676
rect 224368 9664 224374 9716
rect 225690 9664 225696 9716
rect 225748 9664 225754 9716
rect 227530 9664 227536 9716
rect 227588 9704 227594 9716
rect 229094 9704 229100 9716
rect 227588 9676 229100 9704
rect 227588 9664 227594 9676
rect 229094 9664 229100 9676
rect 229152 9664 229158 9716
rect 229186 9664 229192 9716
rect 229244 9704 229250 9716
rect 229244 9676 229784 9704
rect 229244 9664 229250 9676
rect 214926 9636 214932 9648
rect 210844 9608 211568 9636
rect 212644 9608 214932 9636
rect 210844 9596 210850 9608
rect 193217 9571 193275 9577
rect 193217 9537 193229 9571
rect 193263 9568 193275 9571
rect 193582 9568 193588 9580
rect 193263 9540 193588 9568
rect 193263 9537 193275 9540
rect 193217 9531 193275 9537
rect 193582 9528 193588 9540
rect 193640 9528 193646 9580
rect 194689 9571 194747 9577
rect 194689 9537 194701 9571
rect 194735 9568 194747 9571
rect 195790 9568 195796 9580
rect 194735 9540 195796 9568
rect 194735 9537 194747 9540
rect 194689 9531 194747 9537
rect 195790 9528 195796 9540
rect 195848 9528 195854 9580
rect 196161 9571 196219 9577
rect 196161 9537 196173 9571
rect 196207 9568 196219 9571
rect 196618 9568 196624 9580
rect 196207 9540 196624 9568
rect 196207 9537 196219 9540
rect 196161 9531 196219 9537
rect 196618 9528 196624 9540
rect 196676 9528 196682 9580
rect 197173 9571 197231 9577
rect 197173 9537 197185 9571
rect 197219 9568 197231 9571
rect 197538 9568 197544 9580
rect 197219 9540 197544 9568
rect 197219 9537 197231 9540
rect 197173 9531 197231 9537
rect 197538 9528 197544 9540
rect 197596 9528 197602 9580
rect 197906 9528 197912 9580
rect 197964 9528 197970 9580
rect 198645 9571 198703 9577
rect 198645 9537 198657 9571
rect 198691 9568 198703 9571
rect 198826 9568 198832 9580
rect 198691 9540 198832 9568
rect 198691 9537 198703 9540
rect 198645 9531 198703 9537
rect 198826 9528 198832 9540
rect 198884 9528 198890 9580
rect 199838 9528 199844 9580
rect 199896 9528 199902 9580
rect 202325 9571 202383 9577
rect 199948 9540 200620 9568
rect 194410 9500 194416 9512
rect 192496 9472 194416 9500
rect 194410 9460 194416 9472
rect 194468 9460 194474 9512
rect 194594 9460 194600 9512
rect 194652 9500 194658 9512
rect 199948 9500 199976 9540
rect 194652 9472 199976 9500
rect 200592 9500 200620 9540
rect 202325 9537 202337 9571
rect 202371 9568 202383 9571
rect 202690 9568 202696 9580
rect 202371 9540 202696 9568
rect 202371 9537 202383 9540
rect 202325 9531 202383 9537
rect 202690 9528 202696 9540
rect 202748 9528 202754 9580
rect 203061 9571 203119 9577
rect 203061 9537 203073 9571
rect 203107 9568 203119 9571
rect 203426 9568 203432 9580
rect 203107 9540 203432 9568
rect 203107 9537 203119 9540
rect 203061 9531 203119 9537
rect 203426 9528 203432 9540
rect 203484 9528 203490 9580
rect 205818 9528 205824 9580
rect 205876 9528 205882 9580
rect 206554 9528 206560 9580
rect 206612 9528 206618 9580
rect 207658 9528 207664 9580
rect 207716 9528 207722 9580
rect 208302 9528 208308 9580
rect 208360 9528 208366 9580
rect 208946 9528 208952 9580
rect 209004 9528 209010 9580
rect 209314 9528 209320 9580
rect 209372 9568 209378 9580
rect 210237 9571 210295 9577
rect 210237 9568 210249 9571
rect 209372 9540 210249 9568
rect 209372 9528 209378 9540
rect 210237 9537 210249 9540
rect 210283 9537 210295 9571
rect 210237 9531 210295 9537
rect 210878 9528 210884 9580
rect 210936 9528 210942 9580
rect 211540 9577 211568 9608
rect 214926 9596 214932 9608
rect 214984 9596 214990 9648
rect 229756 9636 229784 9676
rect 229830 9664 229836 9716
rect 229888 9664 229894 9716
rect 230658 9664 230664 9716
rect 230716 9704 230722 9716
rect 230716 9676 233004 9704
rect 230716 9664 230722 9676
rect 232866 9636 232872 9648
rect 215036 9608 229600 9636
rect 229756 9608 232872 9636
rect 211525 9571 211583 9577
rect 211525 9537 211537 9571
rect 211571 9537 211583 9571
rect 211525 9531 211583 9537
rect 212534 9528 212540 9580
rect 212592 9568 212598 9580
rect 212813 9571 212871 9577
rect 212813 9568 212825 9571
rect 212592 9540 212825 9568
rect 212592 9528 212598 9540
rect 212813 9537 212825 9540
rect 212859 9537 212871 9571
rect 212813 9531 212871 9537
rect 213454 9528 213460 9580
rect 213512 9528 213518 9580
rect 213914 9528 213920 9580
rect 213972 9568 213978 9580
rect 214101 9571 214159 9577
rect 214101 9568 214113 9571
rect 213972 9540 214113 9568
rect 213972 9528 213978 9540
rect 214101 9537 214113 9540
rect 214147 9537 214159 9571
rect 214101 9531 214159 9537
rect 214374 9528 214380 9580
rect 214432 9568 214438 9580
rect 215036 9568 215064 9608
rect 214432 9540 215064 9568
rect 214432 9528 214438 9540
rect 215294 9528 215300 9580
rect 215352 9568 215358 9580
rect 215389 9571 215447 9577
rect 215389 9568 215401 9571
rect 215352 9540 215401 9568
rect 215352 9528 215358 9540
rect 215389 9537 215401 9540
rect 215435 9537 215447 9571
rect 215389 9531 215447 9537
rect 215478 9528 215484 9580
rect 215536 9568 215542 9580
rect 216033 9571 216091 9577
rect 216033 9568 216045 9571
rect 215536 9540 216045 9568
rect 215536 9528 215542 9540
rect 216033 9537 216045 9540
rect 216079 9537 216091 9571
rect 216033 9531 216091 9537
rect 216674 9528 216680 9580
rect 216732 9528 216738 9580
rect 217962 9528 217968 9580
rect 218020 9528 218026 9580
rect 218606 9528 218612 9580
rect 218664 9528 218670 9580
rect 219250 9528 219256 9580
rect 219308 9528 219314 9580
rect 220538 9528 220544 9580
rect 220596 9528 220602 9580
rect 220814 9528 220820 9580
rect 220872 9568 220878 9580
rect 221185 9571 221243 9577
rect 221185 9568 221197 9571
rect 220872 9540 221197 9568
rect 220872 9528 220878 9540
rect 221185 9537 221197 9540
rect 221231 9537 221243 9571
rect 221185 9531 221243 9537
rect 221826 9528 221832 9580
rect 221884 9528 221890 9580
rect 223114 9528 223120 9580
rect 223172 9528 223178 9580
rect 223298 9528 223304 9580
rect 223356 9568 223362 9580
rect 223761 9571 223819 9577
rect 223761 9568 223773 9571
rect 223356 9540 223773 9568
rect 223356 9528 223362 9540
rect 223761 9537 223773 9540
rect 223807 9537 223819 9571
rect 223761 9531 223819 9537
rect 224310 9528 224316 9580
rect 224368 9568 224374 9580
rect 224368 9540 224540 9568
rect 224368 9528 224374 9540
rect 218238 9500 218244 9512
rect 200592 9472 218244 9500
rect 194652 9460 194658 9472
rect 218238 9460 218244 9472
rect 218296 9460 218302 9512
rect 224402 9500 224408 9512
rect 218348 9472 224408 9500
rect 197262 9392 197268 9444
rect 197320 9432 197326 9444
rect 198093 9435 198151 9441
rect 198093 9432 198105 9435
rect 197320 9404 198105 9432
rect 197320 9392 197326 9404
rect 198093 9401 198105 9404
rect 198139 9401 198151 9435
rect 198093 9395 198151 9401
rect 198182 9392 198188 9444
rect 198240 9432 198246 9444
rect 218348 9432 218376 9472
rect 224402 9460 224408 9472
rect 224460 9460 224466 9512
rect 224512 9500 224540 9540
rect 224586 9528 224592 9580
rect 224644 9528 224650 9580
rect 224770 9528 224776 9580
rect 224828 9528 224834 9580
rect 224957 9571 225015 9577
rect 224957 9537 224969 9571
rect 225003 9568 225015 9571
rect 225509 9571 225567 9577
rect 225509 9568 225521 9571
rect 225003 9540 225521 9568
rect 225003 9537 225015 9540
rect 224957 9531 225015 9537
rect 225509 9537 225521 9540
rect 225555 9537 225567 9571
rect 225509 9531 225567 9537
rect 228177 9571 228235 9577
rect 228177 9537 228189 9571
rect 228223 9568 228235 9571
rect 228358 9568 228364 9580
rect 228223 9540 228364 9568
rect 228223 9537 228235 9540
rect 228177 9531 228235 9537
rect 228358 9528 228364 9540
rect 228416 9528 228422 9580
rect 229462 9500 229468 9512
rect 224512 9472 229468 9500
rect 229462 9460 229468 9472
rect 229520 9460 229526 9512
rect 229572 9500 229600 9608
rect 232866 9596 232872 9608
rect 232924 9596 232930 9648
rect 232976 9636 233004 9676
rect 233510 9664 233516 9716
rect 233568 9664 233574 9716
rect 234338 9664 234344 9716
rect 234396 9664 234402 9716
rect 235074 9664 235080 9716
rect 235132 9664 235138 9716
rect 235810 9664 235816 9716
rect 235868 9704 235874 9716
rect 236546 9704 236552 9716
rect 235868 9676 236552 9704
rect 235868 9664 235874 9676
rect 236546 9664 236552 9676
rect 236604 9664 236610 9716
rect 239416 9676 253934 9704
rect 239416 9636 239444 9676
rect 232976 9608 239444 9636
rect 240226 9596 240232 9648
rect 240284 9596 240290 9648
rect 253906 9636 253934 9676
rect 255682 9664 255688 9716
rect 255740 9664 255746 9716
rect 258442 9664 258448 9716
rect 258500 9704 258506 9716
rect 259914 9704 259920 9716
rect 258500 9676 259920 9704
rect 258500 9664 258506 9676
rect 259914 9664 259920 9676
rect 259972 9664 259978 9716
rect 260006 9664 260012 9716
rect 260064 9664 260070 9716
rect 262122 9704 262128 9716
rect 260806 9676 262128 9704
rect 260806 9636 260834 9676
rect 262122 9664 262128 9676
rect 262180 9664 262186 9716
rect 262214 9664 262220 9716
rect 262272 9704 262278 9716
rect 262401 9707 262459 9713
rect 262401 9704 262413 9707
rect 262272 9676 262413 9704
rect 262272 9664 262278 9676
rect 262401 9673 262413 9676
rect 262447 9673 262459 9707
rect 262401 9667 262459 9673
rect 262858 9664 262864 9716
rect 262916 9664 262922 9716
rect 263134 9664 263140 9716
rect 263192 9704 263198 9716
rect 263321 9707 263379 9713
rect 263321 9704 263333 9707
rect 263192 9676 263333 9704
rect 263192 9664 263198 9676
rect 263321 9673 263333 9676
rect 263367 9673 263379 9707
rect 263321 9667 263379 9673
rect 267829 9707 267887 9713
rect 267829 9673 267841 9707
rect 267875 9704 267887 9707
rect 267875 9676 268240 9704
rect 267875 9673 267887 9676
rect 267829 9667 267887 9673
rect 253906 9608 260834 9636
rect 261021 9639 261079 9645
rect 261021 9605 261033 9639
rect 261067 9636 261079 9639
rect 261067 9608 262260 9636
rect 261067 9605 261079 9608
rect 261021 9599 261079 9605
rect 229649 9571 229707 9577
rect 229649 9537 229661 9571
rect 229695 9568 229707 9571
rect 230014 9568 230020 9580
rect 229695 9540 230020 9568
rect 229695 9537 229707 9540
rect 229649 9531 229707 9537
rect 230014 9528 230020 9540
rect 230072 9528 230078 9580
rect 230198 9528 230204 9580
rect 230256 9568 230262 9580
rect 230753 9571 230811 9577
rect 230753 9568 230765 9571
rect 230256 9540 230765 9568
rect 230256 9528 230262 9540
rect 230753 9537 230765 9540
rect 230799 9537 230811 9571
rect 230753 9531 230811 9537
rect 231026 9528 231032 9580
rect 231084 9568 231090 9580
rect 231397 9571 231455 9577
rect 231397 9568 231409 9571
rect 231084 9540 231409 9568
rect 231084 9528 231090 9540
rect 231397 9537 231409 9540
rect 231443 9537 231455 9571
rect 231397 9531 231455 9537
rect 233329 9571 233387 9577
rect 233329 9537 233341 9571
rect 233375 9568 233387 9571
rect 234062 9568 234068 9580
rect 233375 9540 234068 9568
rect 233375 9537 233387 9540
rect 233329 9531 233387 9537
rect 234062 9528 234068 9540
rect 234120 9528 234126 9580
rect 234154 9528 234160 9580
rect 234212 9528 234218 9580
rect 234890 9528 234896 9580
rect 234948 9528 234954 9580
rect 235810 9528 235816 9580
rect 235868 9528 235874 9580
rect 235902 9528 235908 9580
rect 235960 9568 235966 9580
rect 235997 9571 236055 9577
rect 235997 9568 236009 9571
rect 235960 9540 236009 9568
rect 235960 9528 235966 9540
rect 235997 9537 236009 9540
rect 236043 9537 236055 9571
rect 235997 9531 236055 9537
rect 239674 9528 239680 9580
rect 239732 9528 239738 9580
rect 241238 9528 241244 9580
rect 241296 9528 241302 9580
rect 241348 9540 241652 9568
rect 235442 9500 235448 9512
rect 229572 9472 235448 9500
rect 235442 9460 235448 9472
rect 235500 9500 235506 9512
rect 235828 9500 235856 9528
rect 241348 9500 241376 9540
rect 235500 9472 235856 9500
rect 235920 9472 241376 9500
rect 235500 9460 235506 9472
rect 198240 9404 218376 9432
rect 218425 9435 218483 9441
rect 198240 9392 198246 9404
rect 218425 9401 218437 9435
rect 218471 9432 218483 9435
rect 219158 9432 219164 9444
rect 218471 9404 219164 9432
rect 218471 9401 218483 9404
rect 218425 9395 218483 9401
rect 219158 9392 219164 9404
rect 219216 9392 219222 9444
rect 221001 9435 221059 9441
rect 221001 9401 221013 9435
rect 221047 9432 221059 9435
rect 222102 9432 222108 9444
rect 221047 9404 222108 9432
rect 221047 9401 221059 9404
rect 221001 9395 221059 9401
rect 222102 9392 222108 9404
rect 222160 9392 222166 9444
rect 222194 9392 222200 9444
rect 222252 9432 222258 9444
rect 234614 9432 234620 9444
rect 222252 9404 234620 9432
rect 222252 9392 222258 9404
rect 234614 9392 234620 9404
rect 234672 9392 234678 9444
rect 235534 9392 235540 9444
rect 235592 9432 235598 9444
rect 235920 9432 235948 9472
rect 241514 9460 241520 9512
rect 241572 9460 241578 9512
rect 241624 9500 241652 9540
rect 242710 9528 242716 9580
rect 242768 9568 242774 9580
rect 243541 9571 243599 9577
rect 243541 9568 243553 9571
rect 242768 9540 243553 9568
rect 242768 9528 242774 9540
rect 243541 9537 243553 9540
rect 243587 9537 243599 9571
rect 243541 9531 243599 9537
rect 244918 9528 244924 9580
rect 244976 9568 244982 9580
rect 246117 9571 246175 9577
rect 246117 9568 246129 9571
rect 244976 9540 246129 9568
rect 244976 9528 244982 9540
rect 246117 9537 246129 9540
rect 246163 9537 246175 9571
rect 246117 9531 246175 9537
rect 247862 9528 247868 9580
rect 247920 9568 247926 9580
rect 248693 9571 248751 9577
rect 248693 9568 248705 9571
rect 247920 9540 248705 9568
rect 247920 9528 247926 9540
rect 248693 9537 248705 9540
rect 248739 9537 248751 9571
rect 248693 9531 248751 9537
rect 250070 9528 250076 9580
rect 250128 9568 250134 9580
rect 251269 9571 251327 9577
rect 251269 9568 251281 9571
rect 250128 9540 251281 9568
rect 250128 9528 250134 9540
rect 251269 9537 251281 9540
rect 251315 9537 251327 9571
rect 251269 9531 251327 9537
rect 253106 9528 253112 9580
rect 253164 9568 253170 9580
rect 253845 9571 253903 9577
rect 253845 9568 253857 9571
rect 253164 9540 253857 9568
rect 253164 9528 253170 9540
rect 253845 9537 253857 9540
rect 253891 9537 253903 9571
rect 253845 9531 253903 9537
rect 255866 9528 255872 9580
rect 255924 9528 255930 9580
rect 257890 9528 257896 9580
rect 257948 9528 257954 9580
rect 257985 9571 258043 9577
rect 257985 9537 257997 9571
rect 258031 9568 258043 9571
rect 259178 9568 259184 9580
rect 258031 9540 259184 9568
rect 258031 9537 258043 9540
rect 257985 9531 258043 9537
rect 259178 9528 259184 9540
rect 259236 9528 259242 9580
rect 259365 9571 259423 9577
rect 259365 9537 259377 9571
rect 259411 9568 259423 9571
rect 259825 9571 259883 9577
rect 259825 9568 259837 9571
rect 259411 9540 259837 9568
rect 259411 9537 259423 9540
rect 259365 9531 259423 9537
rect 259825 9537 259837 9540
rect 259871 9537 259883 9571
rect 259825 9531 259883 9537
rect 259914 9528 259920 9580
rect 259972 9568 259978 9580
rect 260650 9568 260656 9580
rect 259972 9540 260656 9568
rect 259972 9528 259978 9540
rect 260650 9528 260656 9540
rect 260708 9528 260714 9580
rect 260837 9571 260895 9577
rect 260837 9537 260849 9571
rect 260883 9568 260895 9571
rect 261202 9568 261208 9580
rect 260883 9540 261208 9568
rect 260883 9537 260895 9540
rect 260837 9531 260895 9537
rect 261202 9528 261208 9540
rect 261260 9568 261266 9580
rect 262232 9577 262260 9608
rect 264698 9596 264704 9648
rect 264756 9636 264762 9648
rect 268102 9636 268108 9648
rect 264756 9608 268108 9636
rect 264756 9596 264762 9608
rect 268102 9596 268108 9608
rect 268160 9596 268166 9648
rect 261757 9571 261815 9577
rect 261757 9568 261769 9571
rect 261260 9540 261769 9568
rect 261260 9528 261266 9540
rect 261757 9537 261769 9540
rect 261803 9537 261815 9571
rect 261757 9531 261815 9537
rect 262217 9571 262275 9577
rect 262217 9537 262229 9571
rect 262263 9537 262275 9571
rect 262217 9531 262275 9537
rect 262858 9528 262864 9580
rect 262916 9568 262922 9580
rect 263229 9571 263287 9577
rect 263229 9568 263241 9571
rect 262916 9540 263241 9568
rect 262916 9528 262922 9540
rect 263229 9537 263241 9540
rect 263275 9537 263287 9571
rect 263229 9531 263287 9537
rect 263962 9528 263968 9580
rect 264020 9568 264026 9580
rect 264149 9571 264207 9577
rect 264149 9568 264161 9571
rect 264020 9540 264161 9568
rect 264020 9528 264026 9540
rect 264149 9537 264161 9540
rect 264195 9537 264207 9571
rect 264149 9531 264207 9537
rect 264333 9571 264391 9577
rect 264333 9537 264345 9571
rect 264379 9568 264391 9571
rect 265066 9568 265072 9580
rect 264379 9540 265072 9568
rect 264379 9537 264391 9540
rect 264333 9531 264391 9537
rect 265066 9528 265072 9540
rect 265124 9568 265130 9580
rect 265161 9571 265219 9577
rect 265161 9568 265173 9571
rect 265124 9540 265173 9568
rect 265124 9528 265130 9540
rect 265161 9537 265173 9540
rect 265207 9568 265219 9571
rect 265986 9568 265992 9580
rect 265207 9540 265992 9568
rect 265207 9537 265219 9540
rect 265161 9531 265219 9537
rect 265986 9528 265992 9540
rect 266044 9528 266050 9580
rect 267093 9571 267151 9577
rect 267093 9537 267105 9571
rect 267139 9568 267151 9571
rect 267826 9568 267832 9580
rect 267139 9540 267832 9568
rect 267139 9537 267151 9540
rect 267093 9531 267151 9537
rect 267826 9528 267832 9540
rect 267884 9528 267890 9580
rect 268212 9577 268240 9676
rect 268197 9571 268255 9577
rect 268197 9537 268209 9571
rect 268243 9568 268255 9571
rect 268838 9568 268844 9580
rect 268243 9540 268844 9568
rect 268243 9537 268255 9540
rect 268197 9531 268255 9537
rect 268838 9528 268844 9540
rect 268896 9528 268902 9580
rect 269482 9528 269488 9580
rect 269540 9528 269546 9580
rect 270129 9571 270187 9577
rect 270129 9537 270141 9571
rect 270175 9568 270187 9571
rect 271230 9568 271236 9580
rect 270175 9540 271236 9568
rect 270175 9537 270187 9540
rect 270129 9531 270187 9537
rect 271230 9528 271236 9540
rect 271288 9528 271294 9580
rect 241624 9472 243676 9500
rect 243538 9432 243544 9444
rect 235592 9404 235948 9432
rect 236104 9404 243544 9432
rect 235592 9392 235598 9404
rect 178000 9336 187188 9364
rect 178000 9324 178006 9336
rect 190914 9324 190920 9376
rect 190972 9324 190978 9376
rect 195514 9324 195520 9376
rect 195572 9364 195578 9376
rect 200666 9364 200672 9376
rect 195572 9336 200672 9364
rect 195572 9324 195578 9336
rect 200666 9324 200672 9336
rect 200724 9324 200730 9376
rect 206373 9367 206431 9373
rect 206373 9333 206385 9367
rect 206419 9364 206431 9367
rect 207382 9364 207388 9376
rect 206419 9336 207388 9364
rect 206419 9333 206431 9336
rect 206373 9327 206431 9333
rect 207382 9324 207388 9336
rect 207440 9324 207446 9376
rect 208118 9324 208124 9376
rect 208176 9324 208182 9376
rect 208762 9324 208768 9376
rect 208820 9324 208826 9376
rect 210050 9324 210056 9376
rect 210108 9324 210114 9376
rect 210697 9367 210755 9373
rect 210697 9333 210709 9367
rect 210743 9364 210755 9367
rect 211246 9364 211252 9376
rect 210743 9336 211252 9364
rect 210743 9333 210755 9336
rect 210697 9327 210755 9333
rect 211246 9324 211252 9336
rect 211304 9324 211310 9376
rect 211341 9367 211399 9373
rect 211341 9333 211353 9367
rect 211387 9364 211399 9367
rect 212718 9364 212724 9376
rect 211387 9336 212724 9364
rect 211387 9333 211399 9336
rect 211341 9327 211399 9333
rect 212718 9324 212724 9336
rect 212776 9324 212782 9376
rect 213270 9324 213276 9376
rect 213328 9324 213334 9376
rect 213914 9324 213920 9376
rect 213972 9324 213978 9376
rect 214466 9324 214472 9376
rect 214524 9364 214530 9376
rect 215205 9367 215263 9373
rect 215205 9364 215217 9367
rect 214524 9336 215217 9364
rect 214524 9324 214530 9336
rect 215205 9333 215217 9336
rect 215251 9333 215263 9367
rect 215205 9327 215263 9333
rect 215386 9324 215392 9376
rect 215444 9364 215450 9376
rect 215849 9367 215907 9373
rect 215849 9364 215861 9367
rect 215444 9336 215861 9364
rect 215444 9324 215450 9336
rect 215849 9333 215861 9336
rect 215895 9333 215907 9367
rect 215849 9327 215907 9333
rect 216493 9367 216551 9373
rect 216493 9333 216505 9367
rect 216539 9364 216551 9367
rect 217686 9364 217692 9376
rect 216539 9336 217692 9364
rect 216539 9333 216551 9336
rect 216493 9327 216551 9333
rect 217686 9324 217692 9336
rect 217744 9324 217750 9376
rect 217778 9324 217784 9376
rect 217836 9324 217842 9376
rect 219069 9367 219127 9373
rect 219069 9333 219081 9367
rect 219115 9364 219127 9367
rect 219342 9364 219348 9376
rect 219115 9336 219348 9364
rect 219115 9333 219127 9336
rect 219069 9327 219127 9333
rect 219342 9324 219348 9336
rect 219400 9324 219406 9376
rect 220354 9324 220360 9376
rect 220412 9324 220418 9376
rect 221645 9367 221703 9373
rect 221645 9333 221657 9367
rect 221691 9364 221703 9367
rect 222838 9364 222844 9376
rect 221691 9336 222844 9364
rect 221691 9333 221703 9336
rect 221645 9327 221703 9333
rect 222838 9324 222844 9336
rect 222896 9324 222902 9376
rect 222930 9324 222936 9376
rect 222988 9324 222994 9376
rect 223577 9367 223635 9373
rect 223577 9333 223589 9367
rect 223623 9364 223635 9367
rect 225138 9364 225144 9376
rect 223623 9336 225144 9364
rect 223623 9333 223635 9336
rect 223577 9327 223635 9333
rect 225138 9324 225144 9336
rect 225196 9324 225202 9376
rect 225690 9324 225696 9376
rect 225748 9364 225754 9376
rect 228082 9364 228088 9376
rect 225748 9336 228088 9364
rect 225748 9324 225754 9336
rect 228082 9324 228088 9336
rect 228140 9324 228146 9376
rect 228266 9324 228272 9376
rect 228324 9364 228330 9376
rect 228361 9367 228419 9373
rect 228361 9364 228373 9367
rect 228324 9336 228373 9364
rect 228324 9324 228330 9336
rect 228361 9333 228373 9336
rect 228407 9333 228419 9367
rect 228361 9327 228419 9333
rect 229830 9324 229836 9376
rect 229888 9364 229894 9376
rect 230845 9367 230903 9373
rect 230845 9364 230857 9367
rect 229888 9336 230857 9364
rect 229888 9324 229894 9336
rect 230845 9333 230857 9336
rect 230891 9333 230903 9367
rect 230845 9327 230903 9333
rect 231578 9324 231584 9376
rect 231636 9324 231642 9376
rect 232866 9324 232872 9376
rect 232924 9364 232930 9376
rect 236104 9364 236132 9404
rect 243538 9392 243544 9404
rect 243596 9392 243602 9444
rect 243648 9432 243676 9472
rect 243814 9460 243820 9512
rect 243872 9460 243878 9512
rect 245654 9460 245660 9512
rect 245712 9500 245718 9512
rect 246393 9503 246451 9509
rect 246393 9500 246405 9503
rect 245712 9472 246405 9500
rect 245712 9460 245718 9472
rect 246393 9469 246405 9472
rect 246439 9469 246451 9503
rect 246393 9463 246451 9469
rect 248966 9460 248972 9512
rect 249024 9460 249030 9512
rect 251450 9460 251456 9512
rect 251508 9500 251514 9512
rect 251545 9503 251603 9509
rect 251545 9500 251557 9503
rect 251508 9472 251557 9500
rect 251508 9460 251514 9472
rect 251545 9469 251557 9472
rect 251591 9469 251603 9503
rect 251545 9463 251603 9469
rect 254026 9460 254032 9512
rect 254084 9500 254090 9512
rect 254121 9503 254179 9509
rect 254121 9500 254133 9503
rect 254084 9472 254133 9500
rect 254084 9460 254090 9472
rect 254121 9469 254133 9472
rect 254167 9469 254179 9503
rect 254121 9463 254179 9469
rect 255222 9460 255228 9512
rect 255280 9500 255286 9512
rect 256421 9503 256479 9509
rect 256421 9500 256433 9503
rect 255280 9472 256433 9500
rect 255280 9460 255286 9472
rect 256421 9469 256433 9472
rect 256467 9469 256479 9503
rect 256421 9463 256479 9469
rect 256697 9503 256755 9509
rect 256697 9469 256709 9503
rect 256743 9500 256755 9503
rect 256786 9500 256792 9512
rect 256743 9472 256792 9500
rect 256743 9469 256755 9472
rect 256697 9463 256755 9469
rect 256786 9460 256792 9472
rect 256844 9460 256850 9512
rect 258166 9460 258172 9512
rect 258224 9500 258230 9512
rect 258224 9472 258672 9500
rect 258224 9460 258230 9472
rect 246666 9432 246672 9444
rect 243648 9404 246672 9432
rect 246666 9392 246672 9404
rect 246724 9392 246730 9444
rect 246758 9392 246764 9444
rect 246816 9432 246822 9444
rect 257982 9432 257988 9444
rect 246816 9404 257988 9432
rect 246816 9392 246822 9404
rect 257982 9392 257988 9404
rect 258040 9392 258046 9444
rect 232924 9336 236132 9364
rect 232924 9324 232930 9336
rect 236178 9324 236184 9376
rect 236236 9324 236242 9376
rect 236546 9324 236552 9376
rect 236604 9364 236610 9376
rect 237190 9364 237196 9376
rect 236604 9336 237196 9364
rect 236604 9324 236610 9336
rect 237190 9324 237196 9336
rect 237248 9324 237254 9376
rect 238110 9324 238116 9376
rect 238168 9364 238174 9376
rect 240321 9367 240379 9373
rect 240321 9364 240333 9367
rect 238168 9336 240333 9364
rect 238168 9324 238174 9336
rect 240321 9333 240333 9336
rect 240367 9333 240379 9367
rect 240321 9327 240379 9333
rect 243170 9324 243176 9376
rect 243228 9364 243234 9376
rect 254118 9364 254124 9376
rect 243228 9336 254124 9364
rect 243228 9324 243234 9336
rect 254118 9324 254124 9336
rect 254176 9324 254182 9376
rect 258074 9324 258080 9376
rect 258132 9364 258138 9376
rect 258169 9367 258227 9373
rect 258169 9364 258181 9367
rect 258132 9336 258181 9364
rect 258132 9324 258138 9336
rect 258169 9333 258181 9336
rect 258215 9333 258227 9367
rect 258644 9364 258672 9472
rect 258718 9460 258724 9512
rect 258776 9500 258782 9512
rect 258997 9503 259055 9509
rect 258997 9500 259009 9503
rect 258776 9472 259009 9500
rect 258776 9460 258782 9472
rect 258997 9469 259009 9472
rect 259043 9469 259055 9503
rect 258997 9463 259055 9469
rect 261478 9460 261484 9512
rect 261536 9500 261542 9512
rect 261573 9503 261631 9509
rect 261573 9500 261585 9503
rect 261536 9472 261585 9500
rect 261536 9460 261542 9472
rect 261573 9469 261585 9472
rect 261619 9469 261631 9503
rect 261573 9463 261631 9469
rect 262122 9460 262128 9512
rect 262180 9500 262186 9512
rect 264977 9503 265035 9509
rect 264977 9500 264989 9503
rect 262180 9472 264989 9500
rect 262180 9460 262186 9472
rect 264977 9469 264989 9472
rect 265023 9500 265035 9503
rect 265342 9500 265348 9512
rect 265023 9472 265348 9500
rect 265023 9469 265035 9472
rect 264977 9463 265035 9469
rect 265342 9460 265348 9472
rect 265400 9460 265406 9512
rect 265805 9503 265863 9509
rect 265805 9469 265817 9503
rect 265851 9500 265863 9503
rect 265894 9500 265900 9512
rect 265851 9472 265900 9500
rect 265851 9469 265863 9472
rect 265805 9463 265863 9469
rect 265894 9460 265900 9472
rect 265952 9460 265958 9512
rect 266722 9460 266728 9512
rect 266780 9500 266786 9512
rect 267642 9500 267648 9512
rect 266780 9472 267648 9500
rect 266780 9460 266786 9472
rect 267642 9460 267648 9472
rect 267700 9460 267706 9512
rect 267844 9500 267872 9528
rect 268470 9500 268476 9512
rect 267844 9472 268476 9500
rect 268470 9460 268476 9472
rect 268528 9460 268534 9512
rect 268654 9460 268660 9512
rect 268712 9500 268718 9512
rect 269301 9503 269359 9509
rect 269301 9500 269313 9503
rect 268712 9472 269313 9500
rect 268712 9460 268718 9472
rect 269301 9469 269313 9472
rect 269347 9469 269359 9503
rect 269301 9463 269359 9469
rect 270402 9460 270408 9512
rect 270460 9460 270466 9512
rect 263686 9392 263692 9444
rect 263744 9432 263750 9444
rect 263744 9404 270448 9432
rect 263744 9392 263750 9404
rect 270420 9376 270448 9404
rect 261478 9364 261484 9376
rect 258644 9336 261484 9364
rect 258169 9327 258227 9333
rect 261478 9324 261484 9336
rect 261536 9324 261542 9376
rect 261570 9324 261576 9376
rect 261628 9364 261634 9376
rect 261941 9367 261999 9373
rect 261941 9364 261953 9367
rect 261628 9336 261953 9364
rect 261628 9324 261634 9336
rect 261941 9333 261953 9336
rect 261987 9333 261999 9367
rect 261941 9327 261999 9333
rect 262030 9324 262036 9376
rect 262088 9364 262094 9376
rect 263778 9364 263784 9376
rect 262088 9336 263784 9364
rect 262088 9324 262094 9336
rect 263778 9324 263784 9336
rect 263836 9324 263842 9376
rect 264054 9324 264060 9376
rect 264112 9364 264118 9376
rect 264517 9367 264575 9373
rect 264517 9364 264529 9367
rect 264112 9336 264529 9364
rect 264112 9324 264118 9336
rect 264517 9333 264529 9336
rect 264563 9333 264575 9367
rect 264517 9327 264575 9333
rect 265345 9367 265403 9373
rect 265345 9333 265357 9367
rect 265391 9364 265403 9367
rect 265526 9364 265532 9376
rect 265391 9336 265532 9364
rect 265391 9333 265403 9336
rect 265345 9327 265403 9333
rect 265526 9324 265532 9336
rect 265584 9324 265590 9376
rect 265618 9324 265624 9376
rect 265676 9364 265682 9376
rect 266173 9367 266231 9373
rect 266173 9364 266185 9367
rect 265676 9336 266185 9364
rect 265676 9324 265682 9336
rect 266173 9333 266185 9336
rect 266219 9333 266231 9367
rect 266173 9327 266231 9333
rect 266998 9324 267004 9376
rect 267056 9364 267062 9376
rect 267185 9367 267243 9373
rect 267185 9364 267197 9367
rect 267056 9336 267197 9364
rect 267056 9324 267062 9336
rect 267185 9333 267197 9336
rect 267231 9333 267243 9367
rect 267185 9327 267243 9333
rect 268194 9324 268200 9376
rect 268252 9364 268258 9376
rect 268473 9367 268531 9373
rect 268473 9364 268485 9367
rect 268252 9336 268485 9364
rect 268252 9324 268258 9336
rect 268473 9333 268485 9336
rect 268519 9364 268531 9367
rect 269298 9364 269304 9376
rect 268519 9336 269304 9364
rect 268519 9333 268531 9336
rect 268473 9327 268531 9333
rect 269298 9324 269304 9336
rect 269356 9324 269362 9376
rect 269669 9367 269727 9373
rect 269669 9333 269681 9367
rect 269715 9364 269727 9367
rect 269850 9364 269856 9376
rect 269715 9336 269856 9364
rect 269715 9333 269727 9336
rect 269669 9327 269727 9333
rect 269850 9324 269856 9336
rect 269908 9324 269914 9376
rect 270402 9324 270408 9376
rect 270460 9324 270466 9376
rect 1104 9274 271492 9296
rect 1104 9222 34748 9274
rect 34800 9222 34812 9274
rect 34864 9222 34876 9274
rect 34928 9222 34940 9274
rect 34992 9222 35004 9274
rect 35056 9222 102345 9274
rect 102397 9222 102409 9274
rect 102461 9222 102473 9274
rect 102525 9222 102537 9274
rect 102589 9222 102601 9274
rect 102653 9222 169942 9274
rect 169994 9222 170006 9274
rect 170058 9222 170070 9274
rect 170122 9222 170134 9274
rect 170186 9222 170198 9274
rect 170250 9222 237539 9274
rect 237591 9222 237603 9274
rect 237655 9222 237667 9274
rect 237719 9222 237731 9274
rect 237783 9222 237795 9274
rect 237847 9222 271492 9274
rect 1104 9200 271492 9222
rect 1394 9120 1400 9172
rect 1452 9160 1458 9172
rect 1765 9163 1823 9169
rect 1765 9160 1777 9163
rect 1452 9132 1777 9160
rect 1452 9120 1458 9132
rect 1765 9129 1777 9132
rect 1811 9129 1823 9163
rect 1765 9123 1823 9129
rect 2406 9120 2412 9172
rect 2464 9160 2470 9172
rect 23106 9160 23112 9172
rect 2464 9132 23112 9160
rect 2464 9120 2470 9132
rect 23106 9120 23112 9132
rect 23164 9120 23170 9172
rect 23201 9163 23259 9169
rect 23201 9129 23213 9163
rect 23247 9160 23259 9163
rect 25130 9160 25136 9172
rect 23247 9132 25136 9160
rect 23247 9129 23259 9132
rect 23201 9123 23259 9129
rect 25130 9120 25136 9132
rect 25188 9120 25194 9172
rect 27706 9120 27712 9172
rect 27764 9160 27770 9172
rect 27764 9132 31432 9160
rect 27764 9120 27770 9132
rect 12802 9052 12808 9104
rect 12860 9092 12866 9104
rect 31294 9092 31300 9104
rect 12860 9064 31300 9092
rect 12860 9052 12866 9064
rect 31294 9052 31300 9064
rect 31352 9052 31358 9104
rect 2498 8984 2504 9036
rect 2556 9024 2562 9036
rect 22738 9024 22744 9036
rect 2556 8996 22744 9024
rect 2556 8984 2562 8996
rect 22738 8984 22744 8996
rect 22796 8984 22802 9036
rect 22830 8984 22836 9036
rect 22888 8984 22894 9036
rect 23661 9027 23719 9033
rect 23661 8993 23673 9027
rect 23707 9024 23719 9027
rect 23934 9024 23940 9036
rect 23707 8996 23940 9024
rect 23707 8993 23719 8996
rect 23661 8987 23719 8993
rect 23934 8984 23940 8996
rect 23992 8984 23998 9036
rect 24854 8984 24860 9036
rect 24912 9024 24918 9036
rect 24912 8996 25176 9024
rect 24912 8984 24918 8996
rect 3142 8916 3148 8968
rect 3200 8916 3206 8968
rect 8202 8916 8208 8968
rect 8260 8956 8266 8968
rect 8297 8959 8355 8965
rect 8297 8956 8309 8959
rect 8260 8928 8309 8956
rect 8260 8916 8266 8928
rect 8297 8925 8309 8928
rect 8343 8925 8355 8959
rect 8297 8919 8355 8925
rect 10502 8916 10508 8968
rect 10560 8916 10566 8968
rect 11238 8916 11244 8968
rect 11296 8916 11302 8968
rect 13446 8916 13452 8968
rect 13504 8916 13510 8968
rect 23017 8959 23075 8965
rect 23017 8925 23029 8959
rect 23063 8956 23075 8959
rect 23842 8956 23848 8968
rect 23063 8928 23848 8956
rect 23063 8925 23075 8928
rect 23017 8919 23075 8925
rect 23842 8916 23848 8928
rect 23900 8956 23906 8968
rect 24118 8956 24124 8968
rect 23900 8928 24124 8956
rect 23900 8916 23906 8928
rect 24118 8916 24124 8928
rect 24176 8956 24182 8968
rect 25038 8956 25044 8968
rect 24176 8928 25044 8956
rect 24176 8916 24182 8928
rect 25038 8916 25044 8928
rect 25096 8916 25102 8968
rect 25148 8956 25176 8996
rect 26234 8984 26240 9036
rect 26292 9024 26298 9036
rect 27157 9027 27215 9033
rect 27157 9024 27169 9027
rect 26292 8996 27169 9024
rect 26292 8984 26298 8996
rect 27157 8993 27169 8996
rect 27203 8993 27215 9027
rect 31404 9024 31432 9132
rect 31754 9120 31760 9172
rect 31812 9160 31818 9172
rect 33597 9163 33655 9169
rect 33597 9160 33609 9163
rect 31812 9132 33609 9160
rect 31812 9120 31818 9132
rect 33597 9129 33609 9132
rect 33643 9129 33655 9163
rect 33597 9123 33655 9129
rect 35158 9120 35164 9172
rect 35216 9120 35222 9172
rect 41230 9120 41236 9172
rect 41288 9160 41294 9172
rect 41874 9160 41880 9172
rect 41288 9132 41880 9160
rect 41288 9120 41294 9132
rect 41874 9120 41880 9132
rect 41932 9120 41938 9172
rect 53190 9120 53196 9172
rect 53248 9120 53254 9172
rect 56410 9160 56416 9172
rect 55324 9132 56416 9160
rect 31478 9052 31484 9104
rect 31536 9092 31542 9104
rect 45922 9092 45928 9104
rect 31536 9064 45928 9092
rect 31536 9052 31542 9064
rect 45922 9052 45928 9064
rect 45980 9052 45986 9104
rect 46198 9052 46204 9104
rect 46256 9092 46262 9104
rect 55324 9092 55352 9132
rect 56410 9120 56416 9132
rect 56468 9120 56474 9172
rect 57514 9120 57520 9172
rect 57572 9120 57578 9172
rect 59170 9120 59176 9172
rect 59228 9120 59234 9172
rect 59998 9120 60004 9172
rect 60056 9120 60062 9172
rect 62758 9120 62764 9172
rect 62816 9120 62822 9172
rect 64046 9120 64052 9172
rect 64104 9160 64110 9172
rect 64104 9132 64874 9160
rect 64104 9120 64110 9132
rect 46256 9064 55352 9092
rect 46256 9052 46262 9064
rect 55398 9052 55404 9104
rect 55456 9092 55462 9104
rect 64690 9092 64696 9104
rect 55456 9064 64696 9092
rect 55456 9052 55462 9064
rect 64690 9052 64696 9064
rect 64748 9052 64754 9104
rect 64846 9092 64874 9132
rect 66346 9120 66352 9172
rect 66404 9120 66410 9172
rect 66456 9132 67220 9160
rect 66456 9092 66484 9132
rect 64846 9064 66484 9092
rect 67192 9092 67220 9132
rect 67266 9120 67272 9172
rect 67324 9160 67330 9172
rect 88242 9160 88248 9172
rect 67324 9132 88248 9160
rect 67324 9120 67330 9132
rect 88242 9120 88248 9132
rect 88300 9120 88306 9172
rect 88334 9120 88340 9172
rect 88392 9160 88398 9172
rect 88429 9163 88487 9169
rect 88429 9160 88441 9163
rect 88392 9132 88441 9160
rect 88392 9120 88398 9132
rect 88429 9129 88441 9132
rect 88475 9129 88487 9163
rect 88429 9123 88487 9129
rect 90174 9120 90180 9172
rect 90232 9120 90238 9172
rect 90560 9132 96108 9160
rect 90560 9092 90588 9132
rect 67192 9064 90588 9092
rect 96080 9092 96108 9132
rect 96154 9120 96160 9172
rect 96212 9120 96218 9172
rect 97166 9120 97172 9172
rect 97224 9160 97230 9172
rect 97224 9132 97488 9160
rect 97224 9120 97230 9132
rect 97460 9092 97488 9132
rect 97994 9120 98000 9172
rect 98052 9120 98058 9172
rect 98086 9120 98092 9172
rect 98144 9160 98150 9172
rect 100110 9160 100116 9172
rect 98144 9132 100116 9160
rect 98144 9120 98150 9132
rect 100110 9120 100116 9132
rect 100168 9120 100174 9172
rect 102686 9120 102692 9172
rect 102744 9160 102750 9172
rect 107562 9160 107568 9172
rect 102744 9132 107568 9160
rect 102744 9120 102750 9132
rect 107562 9120 107568 9132
rect 107620 9120 107626 9172
rect 107654 9120 107660 9172
rect 107712 9160 107718 9172
rect 112714 9160 112720 9172
rect 107712 9132 112720 9160
rect 107712 9120 107718 9132
rect 112714 9120 112720 9132
rect 112772 9120 112778 9172
rect 120997 9163 121055 9169
rect 120997 9129 121009 9163
rect 121043 9160 121055 9163
rect 121362 9160 121368 9172
rect 121043 9132 121368 9160
rect 121043 9129 121055 9132
rect 120997 9123 121055 9129
rect 121362 9120 121368 9132
rect 121420 9120 121426 9172
rect 121917 9163 121975 9169
rect 121917 9129 121929 9163
rect 121963 9160 121975 9163
rect 122466 9160 122472 9172
rect 121963 9132 122472 9160
rect 121963 9129 121975 9132
rect 121917 9123 121975 9129
rect 122466 9120 122472 9132
rect 122524 9120 122530 9172
rect 122742 9120 122748 9172
rect 122800 9160 122806 9172
rect 123205 9163 123263 9169
rect 123205 9160 123217 9163
rect 122800 9132 123217 9160
rect 122800 9120 122806 9132
rect 123205 9129 123217 9132
rect 123251 9129 123263 9163
rect 123205 9123 123263 9129
rect 124582 9120 124588 9172
rect 124640 9120 124646 9172
rect 127802 9120 127808 9172
rect 127860 9120 127866 9172
rect 131390 9120 131396 9172
rect 131448 9120 131454 9172
rect 155494 9160 155500 9172
rect 132466 9132 155500 9160
rect 105446 9092 105452 9104
rect 96080 9064 97396 9092
rect 97460 9064 105452 9092
rect 55858 9024 55864 9036
rect 27157 8987 27215 8993
rect 29012 8996 31248 9024
rect 31404 8996 55864 9024
rect 29012 8968 29040 8996
rect 26881 8959 26939 8965
rect 25148 8928 26556 8956
rect 3326 8848 3332 8900
rect 3384 8848 3390 8900
rect 8478 8848 8484 8900
rect 8536 8848 8542 8900
rect 10689 8891 10747 8897
rect 10689 8857 10701 8891
rect 10735 8888 10747 8891
rect 17218 8888 17224 8900
rect 10735 8860 17224 8888
rect 10735 8857 10747 8860
rect 10689 8851 10747 8857
rect 17218 8848 17224 8860
rect 17276 8848 17282 8900
rect 21450 8848 21456 8900
rect 21508 8888 21514 8900
rect 21508 8860 24164 8888
rect 21508 8848 21514 8860
rect 11330 8780 11336 8832
rect 11388 8780 11394 8832
rect 13538 8780 13544 8832
rect 13596 8780 13602 8832
rect 24026 8780 24032 8832
rect 24084 8780 24090 8832
rect 24136 8820 24164 8860
rect 25130 8848 25136 8900
rect 25188 8848 25194 8900
rect 26053 8891 26111 8897
rect 26053 8857 26065 8891
rect 26099 8888 26111 8891
rect 26418 8888 26424 8900
rect 26099 8860 26424 8888
rect 26099 8857 26111 8860
rect 26053 8851 26111 8857
rect 26418 8848 26424 8860
rect 26476 8848 26482 8900
rect 26528 8888 26556 8928
rect 26881 8925 26893 8959
rect 26927 8956 26939 8959
rect 27522 8956 27528 8968
rect 26927 8928 27528 8956
rect 26927 8925 26939 8928
rect 26881 8919 26939 8925
rect 27522 8916 27528 8928
rect 27580 8916 27586 8968
rect 28905 8959 28963 8965
rect 28905 8925 28917 8959
rect 28951 8925 28963 8959
rect 28905 8919 28963 8925
rect 27062 8888 27068 8900
rect 26528 8860 27068 8888
rect 27062 8848 27068 8860
rect 27120 8848 27126 8900
rect 28920 8888 28948 8919
rect 28994 8916 29000 8968
rect 29052 8916 29058 8968
rect 30208 8965 30236 8996
rect 30101 8959 30159 8965
rect 30101 8925 30113 8959
rect 30147 8925 30159 8959
rect 30101 8919 30159 8925
rect 30193 8959 30251 8965
rect 30193 8925 30205 8959
rect 30239 8925 30251 8959
rect 30193 8919 30251 8925
rect 29546 8888 29552 8900
rect 28920 8860 29552 8888
rect 29546 8848 29552 8860
rect 29604 8888 29610 8900
rect 29914 8888 29920 8900
rect 29604 8860 29920 8888
rect 29604 8848 29610 8860
rect 29914 8848 29920 8860
rect 29972 8848 29978 8900
rect 30116 8888 30144 8919
rect 30374 8916 30380 8968
rect 30432 8916 30438 8968
rect 31110 8916 31116 8968
rect 31168 8916 31174 8968
rect 31220 8965 31248 8996
rect 55858 8984 55864 8996
rect 55916 8984 55922 9036
rect 67174 9024 67180 9036
rect 56336 8996 59860 9024
rect 31205 8959 31263 8965
rect 31205 8925 31217 8959
rect 31251 8956 31263 8959
rect 31251 8928 31754 8956
rect 31251 8925 31263 8928
rect 31205 8919 31263 8925
rect 30392 8888 30420 8916
rect 30116 8860 30420 8888
rect 31726 8888 31754 8928
rect 31938 8916 31944 8968
rect 31996 8916 32002 8968
rect 32033 8959 32091 8965
rect 32033 8925 32045 8959
rect 32079 8925 32091 8959
rect 32033 8919 32091 8925
rect 32217 8959 32275 8965
rect 32217 8925 32229 8959
rect 32263 8956 32275 8959
rect 33413 8959 33471 8965
rect 33413 8956 33425 8959
rect 32263 8928 33425 8956
rect 32263 8925 32275 8928
rect 32217 8919 32275 8925
rect 33413 8925 33425 8928
rect 33459 8925 33471 8959
rect 33413 8919 33471 8925
rect 32048 8888 32076 8919
rect 40310 8916 40316 8968
rect 40368 8916 40374 8968
rect 45462 8916 45468 8968
rect 45520 8916 45526 8968
rect 53009 8959 53067 8965
rect 53009 8925 53021 8959
rect 53055 8956 53067 8959
rect 53374 8956 53380 8968
rect 53055 8928 53380 8956
rect 53055 8925 53067 8928
rect 53009 8919 53067 8925
rect 53374 8916 53380 8928
rect 53432 8916 53438 8968
rect 53466 8916 53472 8968
rect 53524 8956 53530 8968
rect 53745 8959 53803 8965
rect 53745 8956 53757 8959
rect 53524 8928 53757 8956
rect 53524 8916 53530 8928
rect 53745 8925 53757 8928
rect 53791 8925 53803 8959
rect 53745 8919 53803 8925
rect 53929 8959 53987 8965
rect 53929 8925 53941 8959
rect 53975 8956 53987 8959
rect 53975 8928 54064 8956
rect 53975 8925 53987 8928
rect 53929 8919 53987 8925
rect 54036 8900 54064 8928
rect 54386 8916 54392 8968
rect 54444 8956 54450 8968
rect 54573 8959 54631 8965
rect 54573 8956 54585 8959
rect 54444 8928 54585 8956
rect 54444 8916 54450 8928
rect 54573 8925 54585 8928
rect 54619 8925 54631 8959
rect 54573 8919 54631 8925
rect 54757 8959 54815 8965
rect 54757 8925 54769 8959
rect 54803 8925 54815 8959
rect 54757 8919 54815 8925
rect 32769 8891 32827 8897
rect 31726 8860 32536 8888
rect 32508 8832 32536 8860
rect 32769 8857 32781 8891
rect 32815 8888 32827 8891
rect 36998 8888 37004 8900
rect 32815 8860 37004 8888
rect 32815 8857 32827 8860
rect 32769 8851 32827 8857
rect 36998 8848 37004 8860
rect 37056 8848 37062 8900
rect 54018 8848 54024 8900
rect 54076 8888 54082 8900
rect 54772 8888 54800 8919
rect 55398 8916 55404 8968
rect 55456 8956 55462 8968
rect 55493 8959 55551 8965
rect 55493 8956 55505 8959
rect 55456 8928 55505 8956
rect 55456 8916 55462 8928
rect 55493 8925 55505 8928
rect 55539 8925 55551 8959
rect 55493 8919 55551 8925
rect 55677 8959 55735 8965
rect 55677 8925 55689 8959
rect 55723 8956 55735 8959
rect 56336 8956 56364 8996
rect 55723 8928 56364 8956
rect 55723 8925 55735 8928
rect 55677 8919 55735 8925
rect 55692 8888 55720 8919
rect 56410 8916 56416 8968
rect 56468 8916 56474 8968
rect 56520 8965 56548 8996
rect 56505 8959 56563 8965
rect 56505 8925 56517 8959
rect 56551 8925 56563 8959
rect 56505 8919 56563 8925
rect 57146 8916 57152 8968
rect 57204 8916 57210 8968
rect 57348 8965 57376 8996
rect 58176 8965 58204 8996
rect 57333 8959 57391 8965
rect 57333 8925 57345 8959
rect 57379 8925 57391 8959
rect 57333 8919 57391 8925
rect 58069 8959 58127 8965
rect 58069 8925 58081 8959
rect 58115 8925 58127 8959
rect 58069 8919 58127 8925
rect 58161 8959 58219 8965
rect 58161 8925 58173 8959
rect 58207 8925 58219 8959
rect 58161 8919 58219 8925
rect 54076 8860 55720 8888
rect 58084 8888 58112 8919
rect 58894 8916 58900 8968
rect 58952 8916 58958 8968
rect 59004 8965 59032 8996
rect 59832 8968 59860 8996
rect 59924 8996 67180 9024
rect 58989 8959 59047 8965
rect 58989 8925 59001 8959
rect 59035 8925 59047 8959
rect 58989 8919 59047 8925
rect 59630 8916 59636 8968
rect 59688 8916 59694 8968
rect 59814 8916 59820 8968
rect 59872 8916 59878 8968
rect 58526 8888 58532 8900
rect 58084 8860 58532 8888
rect 54076 8848 54082 8860
rect 58526 8848 58532 8860
rect 58584 8888 58590 8900
rect 59924 8888 59952 8996
rect 67174 8984 67180 8996
rect 67232 8984 67238 9036
rect 69566 8984 69572 9036
rect 69624 8984 69630 9036
rect 72050 8984 72056 9036
rect 72108 8984 72114 9036
rect 73430 8984 73436 9036
rect 73488 8984 73494 9036
rect 74718 8984 74724 9036
rect 74776 8984 74782 9036
rect 74994 8984 75000 9036
rect 75052 8984 75058 9036
rect 77202 8984 77208 9036
rect 77260 8984 77266 9036
rect 77478 8984 77484 9036
rect 77536 8984 77542 9036
rect 78582 8984 78588 9036
rect 78640 8984 78646 9036
rect 79873 9027 79931 9033
rect 79873 8993 79885 9027
rect 79919 9024 79931 9027
rect 79962 9024 79968 9036
rect 79919 8996 79968 9024
rect 79919 8993 79931 8996
rect 79873 8987 79931 8993
rect 79962 8984 79968 8996
rect 80020 8984 80026 9036
rect 82354 8984 82360 9036
rect 82412 8984 82418 9036
rect 83826 8984 83832 9036
rect 83884 8984 83890 9036
rect 89349 9027 89407 9033
rect 89349 9024 89361 9027
rect 83936 8996 88196 9024
rect 60090 8916 60096 8968
rect 60148 8956 60154 8968
rect 60642 8956 60648 8968
rect 60148 8928 60648 8956
rect 60148 8916 60154 8928
rect 60642 8916 60648 8928
rect 60700 8956 60706 8968
rect 60737 8959 60795 8965
rect 60737 8956 60749 8959
rect 60700 8928 60749 8956
rect 60700 8916 60706 8928
rect 60737 8925 60749 8928
rect 60783 8925 60795 8959
rect 60737 8919 60795 8925
rect 60918 8916 60924 8968
rect 60976 8916 60982 8968
rect 61470 8916 61476 8968
rect 61528 8956 61534 8968
rect 61565 8959 61623 8965
rect 61565 8956 61577 8959
rect 61528 8928 61577 8956
rect 61528 8916 61534 8928
rect 61565 8925 61577 8928
rect 61611 8925 61623 8959
rect 61565 8919 61623 8925
rect 61749 8959 61807 8965
rect 61749 8925 61761 8959
rect 61795 8925 61807 8959
rect 61749 8919 61807 8925
rect 58584 8860 59952 8888
rect 60936 8888 60964 8916
rect 61764 8888 61792 8919
rect 62390 8916 62396 8968
rect 62448 8916 62454 8968
rect 62577 8959 62635 8965
rect 62577 8925 62589 8959
rect 62623 8925 62635 8959
rect 62577 8919 62635 8925
rect 62592 8888 62620 8919
rect 63218 8916 63224 8968
rect 63276 8916 63282 8968
rect 63405 8959 63463 8965
rect 63405 8925 63417 8959
rect 63451 8925 63463 8959
rect 63405 8919 63463 8925
rect 63420 8888 63448 8919
rect 64046 8916 64052 8968
rect 64104 8916 64110 8968
rect 64233 8959 64291 8965
rect 64233 8925 64245 8959
rect 64279 8925 64291 8959
rect 64233 8919 64291 8925
rect 64248 8888 64276 8919
rect 64966 8916 64972 8968
rect 65024 8916 65030 8968
rect 65061 8959 65119 8965
rect 65061 8925 65073 8959
rect 65107 8925 65119 8959
rect 65061 8919 65119 8925
rect 65076 8888 65104 8919
rect 65978 8916 65984 8968
rect 66036 8916 66042 8968
rect 66165 8959 66223 8965
rect 66165 8925 66177 8959
rect 66211 8925 66223 8959
rect 66165 8919 66223 8925
rect 66809 8959 66867 8965
rect 66809 8925 66821 8959
rect 66855 8956 66867 8959
rect 66898 8956 66904 8968
rect 66855 8928 66904 8956
rect 66855 8925 66867 8928
rect 66809 8919 66867 8925
rect 66180 8888 66208 8919
rect 66898 8916 66904 8928
rect 66956 8916 66962 8968
rect 67085 8959 67143 8965
rect 67085 8925 67097 8959
rect 67131 8925 67143 8959
rect 67085 8919 67143 8925
rect 67100 8888 67128 8919
rect 69842 8916 69848 8968
rect 69900 8916 69906 8968
rect 72329 8959 72387 8965
rect 72329 8925 72341 8959
rect 72375 8925 72387 8959
rect 72329 8919 72387 8925
rect 60936 8860 67128 8888
rect 58584 8848 58590 8860
rect 66824 8832 66852 8860
rect 25225 8823 25283 8829
rect 25225 8820 25237 8823
rect 24136 8792 25237 8820
rect 25225 8789 25237 8792
rect 25271 8789 25283 8823
rect 25225 8783 25283 8789
rect 26142 8780 26148 8832
rect 26200 8780 26206 8832
rect 26878 8780 26884 8832
rect 26936 8820 26942 8832
rect 29086 8820 29092 8832
rect 26936 8792 29092 8820
rect 26936 8780 26942 8792
rect 29086 8780 29092 8792
rect 29144 8780 29150 8832
rect 29181 8823 29239 8829
rect 29181 8789 29193 8823
rect 29227 8820 29239 8823
rect 29454 8820 29460 8832
rect 29227 8792 29460 8820
rect 29227 8789 29239 8792
rect 29181 8783 29239 8789
rect 29454 8780 29460 8792
rect 29512 8780 29518 8832
rect 30282 8780 30288 8832
rect 30340 8820 30346 8832
rect 30377 8823 30435 8829
rect 30377 8820 30389 8823
rect 30340 8792 30389 8820
rect 30340 8780 30346 8792
rect 30377 8789 30389 8792
rect 30423 8789 30435 8823
rect 30377 8783 30435 8789
rect 31110 8780 31116 8832
rect 31168 8820 31174 8832
rect 31389 8823 31447 8829
rect 31389 8820 31401 8823
rect 31168 8792 31401 8820
rect 31168 8780 31174 8792
rect 31389 8789 31401 8792
rect 31435 8789 31447 8823
rect 31389 8783 31447 8789
rect 32490 8780 32496 8832
rect 32548 8820 32554 8832
rect 32861 8823 32919 8829
rect 32861 8820 32873 8823
rect 32548 8792 32873 8820
rect 32548 8780 32554 8792
rect 32861 8789 32873 8792
rect 32907 8789 32919 8823
rect 32861 8783 32919 8789
rect 40126 8780 40132 8832
rect 40184 8780 40190 8832
rect 43438 8780 43444 8832
rect 43496 8820 43502 8832
rect 45281 8823 45339 8829
rect 45281 8820 45293 8823
rect 43496 8792 45293 8820
rect 43496 8780 43502 8792
rect 45281 8789 45293 8792
rect 45327 8789 45339 8823
rect 45281 8783 45339 8789
rect 54113 8823 54171 8829
rect 54113 8789 54125 8823
rect 54159 8820 54171 8823
rect 54570 8820 54576 8832
rect 54159 8792 54576 8820
rect 54159 8789 54171 8792
rect 54113 8783 54171 8789
rect 54570 8780 54576 8792
rect 54628 8780 54634 8832
rect 54941 8823 54999 8829
rect 54941 8789 54953 8823
rect 54987 8820 54999 8823
rect 55306 8820 55312 8832
rect 54987 8792 55312 8820
rect 54987 8789 54999 8792
rect 54941 8783 54999 8789
rect 55306 8780 55312 8792
rect 55364 8780 55370 8832
rect 55861 8823 55919 8829
rect 55861 8789 55873 8823
rect 55907 8820 55919 8823
rect 56042 8820 56048 8832
rect 55907 8792 56048 8820
rect 55907 8789 55919 8792
rect 55861 8783 55919 8789
rect 56042 8780 56048 8792
rect 56100 8780 56106 8832
rect 56689 8823 56747 8829
rect 56689 8789 56701 8823
rect 56735 8820 56747 8823
rect 56870 8820 56876 8832
rect 56735 8792 56876 8820
rect 56735 8789 56747 8792
rect 56689 8783 56747 8789
rect 56870 8780 56876 8792
rect 56928 8780 56934 8832
rect 58345 8823 58403 8829
rect 58345 8789 58357 8823
rect 58391 8820 58403 8823
rect 58434 8820 58440 8832
rect 58391 8792 58440 8820
rect 58391 8789 58403 8792
rect 58345 8783 58403 8789
rect 58434 8780 58440 8792
rect 58492 8780 58498 8832
rect 61105 8823 61163 8829
rect 61105 8789 61117 8823
rect 61151 8820 61163 8823
rect 61378 8820 61384 8832
rect 61151 8792 61384 8820
rect 61151 8789 61163 8792
rect 61105 8783 61163 8789
rect 61378 8780 61384 8792
rect 61436 8780 61442 8832
rect 61933 8823 61991 8829
rect 61933 8789 61945 8823
rect 61979 8820 61991 8823
rect 62114 8820 62120 8832
rect 61979 8792 62120 8820
rect 61979 8789 61991 8792
rect 61933 8783 61991 8789
rect 62114 8780 62120 8792
rect 62172 8780 62178 8832
rect 63586 8780 63592 8832
rect 63644 8780 63650 8832
rect 64414 8780 64420 8832
rect 64472 8780 64478 8832
rect 65242 8780 65248 8832
rect 65300 8780 65306 8832
rect 66806 8780 66812 8832
rect 66864 8780 66870 8832
rect 72344 8820 72372 8919
rect 73706 8916 73712 8968
rect 73764 8916 73770 8968
rect 78858 8916 78864 8968
rect 78916 8916 78922 8968
rect 80146 8916 80152 8968
rect 80204 8916 80210 8968
rect 82630 8916 82636 8968
rect 82688 8916 82694 8968
rect 72418 8848 72424 8900
rect 72476 8888 72482 8900
rect 83936 8888 83964 8996
rect 84102 8916 84108 8968
rect 84160 8916 84166 8968
rect 85390 8916 85396 8968
rect 85448 8916 85454 8968
rect 86494 8916 86500 8968
rect 86552 8916 86558 8968
rect 72476 8860 83964 8888
rect 72476 8848 72482 8860
rect 85574 8848 85580 8900
rect 85632 8848 85638 8900
rect 88168 8888 88196 8996
rect 88260 8996 89361 9024
rect 88260 8965 88288 8996
rect 89349 8993 89361 8996
rect 89395 8993 89407 9027
rect 89349 8987 89407 8993
rect 89686 8996 94360 9024
rect 88245 8959 88303 8965
rect 88245 8925 88257 8959
rect 88291 8925 88303 8959
rect 88245 8919 88303 8925
rect 88978 8916 88984 8968
rect 89036 8916 89042 8968
rect 89162 8916 89168 8968
rect 89220 8956 89226 8968
rect 89686 8956 89714 8996
rect 89220 8928 89714 8956
rect 89220 8916 89226 8928
rect 89898 8916 89904 8968
rect 89956 8916 89962 8968
rect 90008 8965 90036 8996
rect 89993 8959 90051 8965
rect 89993 8925 90005 8959
rect 90039 8925 90051 8959
rect 89993 8919 90051 8925
rect 90726 8916 90732 8968
rect 90784 8916 90790 8968
rect 90836 8965 90864 8996
rect 90821 8959 90879 8965
rect 90821 8925 90833 8959
rect 90867 8925 90879 8959
rect 90821 8919 90879 8925
rect 91002 8916 91008 8968
rect 91060 8956 91066 8968
rect 91848 8965 91876 8996
rect 91649 8959 91707 8965
rect 91649 8956 91661 8959
rect 91060 8928 91661 8956
rect 91060 8916 91066 8928
rect 91649 8925 91661 8928
rect 91695 8925 91707 8959
rect 91649 8919 91707 8925
rect 91833 8959 91891 8965
rect 91833 8925 91845 8959
rect 91879 8925 91891 8959
rect 91833 8919 91891 8925
rect 92014 8916 92020 8968
rect 92072 8956 92078 8968
rect 92382 8956 92388 8968
rect 92072 8928 92388 8956
rect 92072 8916 92078 8928
rect 92382 8916 92388 8928
rect 92440 8956 92446 8968
rect 92676 8965 92704 8996
rect 93504 8968 93532 8996
rect 94332 8968 94360 8996
rect 94958 8984 94964 9036
rect 95016 8984 95022 9036
rect 95050 8984 95056 9036
rect 95108 9024 95114 9036
rect 95789 9027 95847 9033
rect 95789 9024 95801 9027
rect 95108 8996 95801 9024
rect 95108 8984 95114 8996
rect 95789 8993 95801 8996
rect 95835 8993 95847 9027
rect 95789 8987 95847 8993
rect 96706 8984 96712 9036
rect 96764 9024 96770 9036
rect 96801 9027 96859 9033
rect 96801 9024 96813 9027
rect 96764 8996 96813 9024
rect 96764 8984 96770 8996
rect 96801 8993 96813 8996
rect 96847 9024 96859 9027
rect 96890 9024 96896 9036
rect 96847 8996 96896 9024
rect 96847 8993 96859 8996
rect 96801 8987 96859 8993
rect 96890 8984 96896 8996
rect 96948 8984 96954 9036
rect 92477 8959 92535 8965
rect 92477 8956 92489 8959
rect 92440 8928 92489 8956
rect 92440 8916 92446 8928
rect 92477 8925 92489 8928
rect 92523 8925 92535 8959
rect 92477 8919 92535 8925
rect 92661 8959 92719 8965
rect 92661 8925 92673 8959
rect 92707 8925 92719 8959
rect 92661 8919 92719 8925
rect 93394 8916 93400 8968
rect 93452 8916 93458 8968
rect 93486 8916 93492 8968
rect 93544 8916 93550 8968
rect 93670 8916 93676 8968
rect 93728 8916 93734 8968
rect 94133 8959 94191 8965
rect 94133 8925 94145 8959
rect 94179 8925 94191 8959
rect 94133 8919 94191 8925
rect 94148 8888 94176 8919
rect 94314 8916 94320 8968
rect 94372 8916 94378 8968
rect 95145 8959 95203 8965
rect 95145 8925 95157 8959
rect 95191 8925 95203 8959
rect 95145 8919 95203 8925
rect 95973 8959 96031 8965
rect 95973 8925 95985 8959
rect 96019 8956 96031 8959
rect 96985 8959 97043 8965
rect 96019 8928 96660 8956
rect 96019 8925 96031 8928
rect 95973 8919 96031 8925
rect 94222 8888 94228 8900
rect 86512 8860 86724 8888
rect 88168 8860 94228 8888
rect 86512 8820 86540 8860
rect 72344 8792 86540 8820
rect 86586 8780 86592 8832
rect 86644 8780 86650 8832
rect 86696 8820 86724 8860
rect 94222 8848 94228 8860
rect 94280 8848 94286 8900
rect 95160 8888 95188 8919
rect 95988 8888 96016 8919
rect 96632 8900 96660 8928
rect 96985 8925 96997 8959
rect 97031 8925 97043 8959
rect 97368 8956 97396 9064
rect 105446 9052 105452 9064
rect 105504 9052 105510 9104
rect 106090 9052 106096 9104
rect 106148 9092 106154 9104
rect 112165 9095 112223 9101
rect 112165 9092 112177 9095
rect 106148 9064 112177 9092
rect 106148 9052 106154 9064
rect 112165 9061 112177 9064
rect 112211 9061 112223 9095
rect 112165 9055 112223 9061
rect 121270 9052 121276 9104
rect 121328 9092 121334 9104
rect 132466 9092 132494 9132
rect 155494 9120 155500 9132
rect 155552 9120 155558 9172
rect 156138 9120 156144 9172
rect 156196 9120 156202 9172
rect 156966 9120 156972 9172
rect 157024 9120 157030 9172
rect 157794 9120 157800 9172
rect 157852 9120 157858 9172
rect 159818 9120 159824 9172
rect 159876 9160 159882 9172
rect 163406 9160 163412 9172
rect 159876 9132 163412 9160
rect 159876 9120 159882 9132
rect 163406 9120 163412 9132
rect 163464 9120 163470 9172
rect 164786 9120 164792 9172
rect 164844 9120 164850 9172
rect 169018 9120 169024 9172
rect 169076 9160 169082 9172
rect 170493 9163 170551 9169
rect 170493 9160 170505 9163
rect 169076 9132 170505 9160
rect 169076 9120 169082 9132
rect 170493 9129 170505 9132
rect 170539 9129 170551 9163
rect 170493 9123 170551 9129
rect 170582 9120 170588 9172
rect 170640 9160 170646 9172
rect 189718 9160 189724 9172
rect 170640 9132 189724 9160
rect 170640 9120 170646 9132
rect 189718 9120 189724 9132
rect 189776 9120 189782 9172
rect 192386 9120 192392 9172
rect 192444 9160 192450 9172
rect 193585 9163 193643 9169
rect 193585 9160 193597 9163
rect 192444 9132 193597 9160
rect 192444 9120 192450 9132
rect 193585 9129 193597 9132
rect 193631 9129 193643 9163
rect 193585 9123 193643 9129
rect 195790 9120 195796 9172
rect 195848 9120 195854 9172
rect 197906 9120 197912 9172
rect 197964 9160 197970 9172
rect 198921 9163 198979 9169
rect 198921 9160 198933 9163
rect 197964 9132 198933 9160
rect 197964 9120 197970 9132
rect 198921 9129 198933 9132
rect 198967 9129 198979 9163
rect 198921 9123 198979 9129
rect 199838 9120 199844 9172
rect 199896 9160 199902 9172
rect 200945 9163 201003 9169
rect 200945 9160 200957 9163
rect 199896 9132 200957 9160
rect 199896 9120 199902 9132
rect 200945 9129 200957 9132
rect 200991 9129 201003 9163
rect 200945 9123 201003 9129
rect 201972 9132 203748 9160
rect 121328 9064 132494 9092
rect 121328 9052 121334 9064
rect 133414 9052 133420 9104
rect 133472 9052 133478 9104
rect 133966 9052 133972 9104
rect 134024 9092 134030 9104
rect 134024 9064 134196 9092
rect 134024 9052 134030 9064
rect 97626 8984 97632 9036
rect 97684 8984 97690 9036
rect 98270 9024 98276 9036
rect 97736 8996 98276 9024
rect 97736 8956 97764 8996
rect 98270 8984 98276 8996
rect 98328 9024 98334 9036
rect 98454 9024 98460 9036
rect 98328 8996 98460 9024
rect 98328 8984 98334 8996
rect 98454 8984 98460 8996
rect 98512 8984 98518 9036
rect 99282 8984 99288 9036
rect 99340 8984 99346 9036
rect 100018 9024 100024 9036
rect 99484 8996 100024 9024
rect 99484 8968 99512 8996
rect 100018 8984 100024 8996
rect 100076 9024 100082 9036
rect 100389 9027 100447 9033
rect 100389 9024 100401 9027
rect 100076 8996 100401 9024
rect 100076 8984 100082 8996
rect 100389 8993 100401 8996
rect 100435 8993 100447 9027
rect 100389 8987 100447 8993
rect 104342 8984 104348 9036
rect 104400 9024 104406 9036
rect 108206 9024 108212 9036
rect 104400 8996 108212 9024
rect 104400 8984 104406 8996
rect 108206 8984 108212 8996
rect 108264 8984 108270 9036
rect 127158 9024 127164 9036
rect 118666 8996 127164 9024
rect 97368 8928 97764 8956
rect 97813 8959 97871 8965
rect 96985 8919 97043 8925
rect 97813 8925 97825 8959
rect 97859 8925 97871 8959
rect 97813 8919 97871 8925
rect 98641 8959 98699 8965
rect 98641 8925 98653 8959
rect 98687 8925 98699 8959
rect 99466 8956 99472 8968
rect 98641 8919 98699 8925
rect 99346 8928 99472 8956
rect 95160 8860 96016 8888
rect 96614 8848 96620 8900
rect 96672 8888 96678 8900
rect 97000 8888 97028 8919
rect 97828 8888 97856 8919
rect 98656 8888 98684 8919
rect 99346 8888 99374 8928
rect 99466 8916 99472 8928
rect 99524 8916 99530 8968
rect 100110 8916 100116 8968
rect 100168 8916 100174 8968
rect 101674 8916 101680 8968
rect 101732 8956 101738 8968
rect 106274 8956 106280 8968
rect 101732 8928 106280 8956
rect 101732 8916 101738 8928
rect 106274 8916 106280 8928
rect 106332 8916 106338 8968
rect 107194 8916 107200 8968
rect 107252 8916 107258 8968
rect 112346 8916 112352 8968
rect 112404 8916 112410 8968
rect 117314 8916 117320 8968
rect 117372 8956 117378 8968
rect 117501 8959 117559 8965
rect 117501 8956 117513 8959
rect 117372 8928 117513 8956
rect 117372 8916 117378 8928
rect 117501 8925 117513 8928
rect 117547 8925 117559 8959
rect 117501 8919 117559 8925
rect 96672 8860 99374 8888
rect 96672 8848 96678 8860
rect 100478 8848 100484 8900
rect 100536 8888 100542 8900
rect 100536 8860 100800 8888
rect 100536 8848 100542 8860
rect 89622 8820 89628 8832
rect 86696 8792 89628 8820
rect 89622 8780 89628 8792
rect 89680 8780 89686 8832
rect 90910 8780 90916 8832
rect 90968 8820 90974 8832
rect 91005 8823 91063 8829
rect 91005 8820 91017 8823
rect 90968 8792 91017 8820
rect 90968 8780 90974 8792
rect 91005 8789 91017 8792
rect 91051 8789 91063 8823
rect 91005 8783 91063 8789
rect 91646 8780 91652 8832
rect 91704 8820 91710 8832
rect 92017 8823 92075 8829
rect 92017 8820 92029 8823
rect 91704 8792 92029 8820
rect 91704 8780 91710 8792
rect 92017 8789 92029 8792
rect 92063 8789 92075 8823
rect 92017 8783 92075 8789
rect 92382 8780 92388 8832
rect 92440 8820 92446 8832
rect 92845 8823 92903 8829
rect 92845 8820 92857 8823
rect 92440 8792 92857 8820
rect 92440 8780 92446 8792
rect 92845 8789 92857 8792
rect 92891 8789 92903 8823
rect 92845 8783 92903 8789
rect 94406 8780 94412 8832
rect 94464 8820 94470 8832
rect 94501 8823 94559 8829
rect 94501 8820 94513 8823
rect 94464 8792 94513 8820
rect 94464 8780 94470 8792
rect 94501 8789 94513 8792
rect 94547 8789 94559 8823
rect 94501 8783 94559 8789
rect 95142 8780 95148 8832
rect 95200 8820 95206 8832
rect 95329 8823 95387 8829
rect 95329 8820 95341 8823
rect 95200 8792 95341 8820
rect 95200 8780 95206 8792
rect 95329 8789 95341 8792
rect 95375 8789 95387 8823
rect 95329 8783 95387 8789
rect 97169 8823 97227 8829
rect 97169 8789 97181 8823
rect 97215 8820 97227 8823
rect 97258 8820 97264 8832
rect 97215 8792 97264 8820
rect 97215 8789 97227 8792
rect 97169 8783 97227 8789
rect 97258 8780 97264 8792
rect 97316 8780 97322 8832
rect 98454 8780 98460 8832
rect 98512 8820 98518 8832
rect 98825 8823 98883 8829
rect 98825 8820 98837 8823
rect 98512 8792 98837 8820
rect 98512 8780 98518 8792
rect 98825 8789 98837 8792
rect 98871 8789 98883 8823
rect 98825 8783 98883 8789
rect 99282 8780 99288 8832
rect 99340 8820 99346 8832
rect 99558 8820 99564 8832
rect 99340 8792 99564 8820
rect 99340 8780 99346 8792
rect 99558 8780 99564 8792
rect 99616 8780 99622 8832
rect 99653 8823 99711 8829
rect 99653 8789 99665 8823
rect 99699 8820 99711 8823
rect 100662 8820 100668 8832
rect 99699 8792 100668 8820
rect 99699 8789 99711 8792
rect 99653 8783 99711 8789
rect 100662 8780 100668 8792
rect 100720 8780 100726 8832
rect 100772 8820 100800 8860
rect 104158 8848 104164 8900
rect 104216 8888 104222 8900
rect 118666 8888 118694 8996
rect 127158 8984 127164 8996
rect 127216 8984 127222 9036
rect 128725 9027 128783 9033
rect 128725 9024 128737 9027
rect 127636 8996 128737 9024
rect 120810 8916 120816 8968
rect 120868 8916 120874 8968
rect 121638 8916 121644 8968
rect 121696 8916 121702 8968
rect 121730 8916 121736 8968
rect 121788 8956 121794 8968
rect 121788 8928 122604 8956
rect 121788 8916 121794 8928
rect 104216 8860 118694 8888
rect 122576 8888 122604 8928
rect 122650 8916 122656 8968
rect 122708 8916 122714 8968
rect 122745 8959 122803 8965
rect 122745 8925 122757 8959
rect 122791 8956 122803 8959
rect 122791 8928 123248 8956
rect 122791 8925 122803 8928
rect 122745 8919 122803 8925
rect 122852 8888 122880 8928
rect 122576 8860 122880 8888
rect 123220 8888 123248 8928
rect 123294 8916 123300 8968
rect 123352 8956 123358 8968
rect 123389 8959 123447 8965
rect 123389 8956 123401 8959
rect 123352 8928 123401 8956
rect 123352 8916 123358 8928
rect 123389 8925 123401 8928
rect 123435 8925 123447 8959
rect 123389 8919 123447 8925
rect 123573 8959 123631 8965
rect 123573 8925 123585 8959
rect 123619 8925 123631 8959
rect 123573 8919 123631 8925
rect 123588 8888 123616 8919
rect 124122 8916 124128 8968
rect 124180 8956 124186 8968
rect 124217 8959 124275 8965
rect 124217 8956 124229 8959
rect 124180 8928 124229 8956
rect 124180 8916 124186 8928
rect 124217 8925 124229 8928
rect 124263 8925 124275 8959
rect 124217 8919 124275 8925
rect 124401 8959 124459 8965
rect 124401 8925 124413 8959
rect 124447 8925 124459 8959
rect 124401 8919 124459 8925
rect 124416 8888 124444 8919
rect 125042 8916 125048 8968
rect 125100 8916 125106 8968
rect 125229 8959 125287 8965
rect 125229 8925 125241 8959
rect 125275 8925 125287 8959
rect 125229 8919 125287 8925
rect 125244 8888 125272 8919
rect 125870 8916 125876 8968
rect 125928 8916 125934 8968
rect 126057 8959 126115 8965
rect 126057 8925 126069 8959
rect 126103 8925 126115 8959
rect 126057 8919 126115 8925
rect 126072 8888 126100 8919
rect 126698 8916 126704 8968
rect 126756 8916 126762 8968
rect 127636 8965 127664 8996
rect 128725 8993 128737 8996
rect 128771 8993 128783 9027
rect 128725 8987 128783 8993
rect 129274 8984 129280 9036
rect 129332 8984 129338 9036
rect 130378 9024 130384 9036
rect 129568 8996 130384 9024
rect 129568 8968 129596 8996
rect 130378 8984 130384 8996
rect 130436 9024 130442 9036
rect 134168 9024 134196 9064
rect 134242 9052 134248 9104
rect 134300 9052 134306 9104
rect 134886 9052 134892 9104
rect 134944 9052 134950 9104
rect 154945 9095 155003 9101
rect 154945 9061 154957 9095
rect 154991 9092 155003 9095
rect 158346 9092 158352 9104
rect 154991 9064 158352 9092
rect 154991 9061 155003 9064
rect 154945 9055 155003 9061
rect 158346 9052 158352 9064
rect 158404 9052 158410 9104
rect 159744 9064 159956 9092
rect 159744 9024 159772 9064
rect 130436 8996 134104 9024
rect 134168 8996 159772 9024
rect 159928 9024 159956 9064
rect 160002 9052 160008 9104
rect 160060 9092 160066 9104
rect 184566 9092 184572 9104
rect 160060 9064 184572 9092
rect 160060 9052 160066 9064
rect 184566 9052 184572 9064
rect 184624 9052 184630 9104
rect 197170 9092 197176 9104
rect 184676 9064 197176 9092
rect 159928 8996 164832 9024
rect 130436 8984 130442 8996
rect 126885 8959 126943 8965
rect 126885 8925 126897 8959
rect 126931 8925 126943 8959
rect 126885 8919 126943 8925
rect 127621 8959 127679 8965
rect 127621 8925 127633 8959
rect 127667 8925 127679 8959
rect 127621 8919 127679 8925
rect 126900 8888 126928 8919
rect 128262 8916 128268 8968
rect 128320 8956 128326 8968
rect 128357 8959 128415 8965
rect 128357 8956 128369 8959
rect 128320 8928 128369 8956
rect 128320 8916 128326 8928
rect 128357 8925 128369 8928
rect 128403 8925 128415 8959
rect 128357 8919 128415 8925
rect 128541 8959 128599 8965
rect 128541 8925 128553 8959
rect 128587 8925 128599 8959
rect 128541 8919 128599 8925
rect 127802 8888 127808 8900
rect 123220 8860 127808 8888
rect 104216 8848 104222 8860
rect 127802 8848 127808 8860
rect 127860 8888 127866 8900
rect 128556 8888 128584 8919
rect 129550 8916 129556 8968
rect 129608 8916 129614 8968
rect 131025 8959 131083 8965
rect 131025 8925 131037 8959
rect 131071 8956 131083 8959
rect 131114 8956 131120 8968
rect 131071 8928 131120 8956
rect 131071 8925 131083 8928
rect 131025 8919 131083 8925
rect 131114 8916 131120 8928
rect 131172 8916 131178 8968
rect 131224 8965 131252 8996
rect 131209 8959 131267 8965
rect 131209 8925 131221 8959
rect 131255 8925 131267 8959
rect 131209 8919 131267 8925
rect 131850 8916 131856 8968
rect 131908 8916 131914 8968
rect 132052 8965 132080 8996
rect 132037 8959 132095 8965
rect 132037 8925 132049 8959
rect 132083 8925 132095 8959
rect 132037 8919 132095 8925
rect 132954 8916 132960 8968
rect 133012 8956 133018 8968
rect 133049 8959 133107 8965
rect 133049 8956 133061 8959
rect 133012 8928 133061 8956
rect 133012 8916 133018 8928
rect 133049 8925 133061 8928
rect 133095 8925 133107 8959
rect 133049 8919 133107 8925
rect 133138 8916 133144 8968
rect 133196 8956 133202 8968
rect 133248 8965 133276 8996
rect 133233 8959 133291 8965
rect 133233 8956 133245 8959
rect 133196 8928 133245 8956
rect 133196 8916 133202 8928
rect 133233 8925 133245 8928
rect 133279 8925 133291 8959
rect 133233 8919 133291 8925
rect 133966 8916 133972 8968
rect 134024 8916 134030 8968
rect 134076 8965 134104 8996
rect 134061 8959 134119 8965
rect 134061 8925 134073 8959
rect 134107 8925 134119 8959
rect 134061 8919 134119 8925
rect 134518 8916 134524 8968
rect 134576 8956 134582 8968
rect 134705 8959 134763 8965
rect 134705 8956 134717 8959
rect 134576 8928 134717 8956
rect 134576 8916 134582 8928
rect 134705 8925 134717 8928
rect 134751 8925 134763 8959
rect 134705 8919 134763 8925
rect 139762 8916 139768 8968
rect 139820 8916 139826 8968
rect 144730 8916 144736 8968
rect 144788 8956 144794 8968
rect 144917 8959 144975 8965
rect 144917 8956 144929 8959
rect 144788 8928 144929 8956
rect 144788 8916 144794 8928
rect 144917 8925 144929 8928
rect 144963 8925 144975 8959
rect 144917 8919 144975 8925
rect 150066 8916 150072 8968
rect 150124 8916 150130 8968
rect 155126 8916 155132 8968
rect 155184 8916 155190 8968
rect 155678 8916 155684 8968
rect 155736 8916 155742 8968
rect 155773 8959 155831 8965
rect 155773 8925 155785 8959
rect 155819 8925 155831 8959
rect 155773 8919 155831 8925
rect 155957 8959 156015 8965
rect 155957 8925 155969 8959
rect 156003 8925 156015 8959
rect 155957 8919 156015 8925
rect 127860 8860 128584 8888
rect 127860 8848 127866 8860
rect 128722 8848 128728 8900
rect 128780 8888 128786 8900
rect 137278 8888 137284 8900
rect 128780 8860 137284 8888
rect 128780 8848 128786 8860
rect 137278 8848 137284 8860
rect 137336 8848 137342 8900
rect 137370 8848 137376 8900
rect 137428 8888 137434 8900
rect 155696 8888 155724 8916
rect 137428 8860 155724 8888
rect 137428 8848 137434 8860
rect 155788 8832 155816 8919
rect 155972 8888 156000 8919
rect 156690 8916 156696 8968
rect 156748 8916 156754 8968
rect 156785 8959 156843 8965
rect 156785 8925 156797 8959
rect 156831 8925 156843 8959
rect 156785 8919 156843 8925
rect 156800 8888 156828 8919
rect 157518 8916 157524 8968
rect 157576 8916 157582 8968
rect 157610 8916 157616 8968
rect 157668 8916 157674 8968
rect 158625 8959 158683 8965
rect 158625 8925 158637 8959
rect 158671 8956 158683 8959
rect 158671 8928 159772 8956
rect 158671 8925 158683 8928
rect 158625 8919 158683 8925
rect 157628 8888 157656 8916
rect 155972 8860 157656 8888
rect 158714 8848 158720 8900
rect 158772 8888 158778 8900
rect 159177 8891 159235 8897
rect 159177 8888 159189 8891
rect 158772 8860 159189 8888
rect 158772 8848 158778 8860
rect 159177 8857 159189 8860
rect 159223 8888 159235 8891
rect 159634 8888 159640 8900
rect 159223 8860 159640 8888
rect 159223 8857 159235 8860
rect 159177 8851 159235 8857
rect 159634 8848 159640 8860
rect 159692 8848 159698 8900
rect 159744 8888 159772 8928
rect 159818 8916 159824 8968
rect 159876 8916 159882 8968
rect 159910 8916 159916 8968
rect 159968 8956 159974 8968
rect 160189 8959 160247 8965
rect 160189 8956 160201 8959
rect 159968 8928 160201 8956
rect 159968 8916 159974 8928
rect 160189 8925 160201 8928
rect 160235 8925 160247 8959
rect 160189 8919 160247 8925
rect 160296 8928 160784 8956
rect 160296 8888 160324 8928
rect 159744 8860 160324 8888
rect 160756 8888 160784 8928
rect 160830 8916 160836 8968
rect 160888 8916 160894 8968
rect 161198 8916 161204 8968
rect 161256 8916 161262 8968
rect 161845 8959 161903 8965
rect 161308 8928 161796 8956
rect 161308 8888 161336 8928
rect 160756 8860 161336 8888
rect 161768 8888 161796 8928
rect 161845 8925 161857 8959
rect 161891 8956 161903 8959
rect 162210 8956 162216 8968
rect 161891 8928 162216 8956
rect 161891 8925 161903 8928
rect 161845 8919 161903 8925
rect 162210 8916 162216 8928
rect 162268 8916 162274 8968
rect 162578 8916 162584 8968
rect 162636 8916 162642 8968
rect 163777 8959 163835 8965
rect 163777 8925 163789 8959
rect 163823 8956 163835 8959
rect 164694 8956 164700 8968
rect 163823 8928 164700 8956
rect 163823 8925 163835 8928
rect 163777 8919 163835 8925
rect 164694 8916 164700 8928
rect 164752 8916 164758 8968
rect 161768 8860 162716 8888
rect 107013 8823 107071 8829
rect 107013 8820 107025 8823
rect 100772 8792 107025 8820
rect 107013 8789 107025 8792
rect 107059 8789 107071 8823
rect 107013 8783 107071 8789
rect 107102 8780 107108 8832
rect 107160 8820 107166 8832
rect 109862 8820 109868 8832
rect 107160 8792 109868 8820
rect 107160 8780 107166 8792
rect 109862 8780 109868 8792
rect 109920 8780 109926 8832
rect 115566 8780 115572 8832
rect 115624 8820 115630 8832
rect 117317 8823 117375 8829
rect 117317 8820 117329 8823
rect 115624 8792 117329 8820
rect 115624 8780 115630 8792
rect 117317 8789 117329 8792
rect 117363 8789 117375 8823
rect 117317 8783 117375 8789
rect 122929 8823 122987 8829
rect 122929 8789 122941 8823
rect 122975 8820 122987 8823
rect 123018 8820 123024 8832
rect 122975 8792 123024 8820
rect 122975 8789 122987 8792
rect 122929 8783 122987 8789
rect 123018 8780 123024 8792
rect 123076 8780 123082 8832
rect 123754 8780 123760 8832
rect 123812 8780 123818 8832
rect 125410 8780 125416 8832
rect 125468 8780 125474 8832
rect 126146 8780 126152 8832
rect 126204 8820 126210 8832
rect 126241 8823 126299 8829
rect 126241 8820 126253 8823
rect 126204 8792 126253 8820
rect 126204 8780 126210 8792
rect 126241 8789 126253 8792
rect 126287 8789 126299 8823
rect 126241 8783 126299 8789
rect 126882 8780 126888 8832
rect 126940 8820 126946 8832
rect 127069 8823 127127 8829
rect 127069 8820 127081 8823
rect 126940 8792 127081 8820
rect 126940 8780 126946 8792
rect 127069 8789 127081 8792
rect 127115 8789 127127 8823
rect 127069 8783 127127 8789
rect 127158 8780 127164 8832
rect 127216 8820 127222 8832
rect 128262 8820 128268 8832
rect 127216 8792 128268 8820
rect 127216 8780 127222 8792
rect 128262 8780 128268 8792
rect 128320 8820 128326 8832
rect 128998 8820 129004 8832
rect 128320 8792 129004 8820
rect 128320 8780 128326 8792
rect 128998 8780 129004 8792
rect 129056 8780 129062 8832
rect 132126 8780 132132 8832
rect 132184 8820 132190 8832
rect 132221 8823 132279 8829
rect 132221 8820 132233 8823
rect 132184 8792 132233 8820
rect 132184 8780 132190 8792
rect 132221 8789 132233 8792
rect 132267 8789 132279 8823
rect 132221 8783 132279 8789
rect 134242 8780 134248 8832
rect 134300 8820 134306 8832
rect 135441 8823 135499 8829
rect 135441 8820 135453 8823
rect 134300 8792 135453 8820
rect 134300 8780 134306 8792
rect 135441 8789 135453 8792
rect 135487 8789 135499 8823
rect 135441 8783 135499 8789
rect 139581 8823 139639 8829
rect 139581 8789 139593 8823
rect 139627 8820 139639 8823
rect 140406 8820 140412 8832
rect 139627 8792 140412 8820
rect 139627 8789 139639 8792
rect 139581 8783 139639 8789
rect 140406 8780 140412 8792
rect 140464 8780 140470 8832
rect 144733 8823 144791 8829
rect 144733 8789 144745 8823
rect 144779 8820 144791 8823
rect 147766 8820 147772 8832
rect 144779 8792 147772 8820
rect 144779 8789 144791 8792
rect 144733 8783 144791 8789
rect 147766 8780 147772 8792
rect 147824 8780 147830 8832
rect 149882 8780 149888 8832
rect 149940 8780 149946 8832
rect 155494 8780 155500 8832
rect 155552 8820 155558 8832
rect 155770 8820 155776 8832
rect 155552 8792 155776 8820
rect 155552 8780 155558 8792
rect 155770 8780 155776 8792
rect 155828 8780 155834 8832
rect 156690 8780 156696 8832
rect 156748 8820 156754 8832
rect 157150 8820 157156 8832
rect 156748 8792 157156 8820
rect 156748 8780 156754 8792
rect 157150 8780 157156 8792
rect 157208 8780 157214 8832
rect 157242 8780 157248 8832
rect 157300 8820 157306 8832
rect 162394 8820 162400 8832
rect 157300 8792 162400 8820
rect 157300 8780 157306 8792
rect 162394 8780 162400 8792
rect 162452 8780 162458 8832
rect 162688 8820 162716 8860
rect 163866 8848 163872 8900
rect 163924 8888 163930 8900
rect 164142 8888 164148 8900
rect 163924 8860 164148 8888
rect 163924 8848 163930 8860
rect 164142 8848 164148 8860
rect 164200 8848 164206 8900
rect 164234 8820 164240 8832
rect 162688 8792 164240 8820
rect 164234 8780 164240 8792
rect 164292 8780 164298 8832
rect 164804 8820 164832 8996
rect 165338 8984 165344 9036
rect 165396 8984 165402 9036
rect 177206 9024 177212 9036
rect 166644 8996 177212 9024
rect 165157 8959 165215 8965
rect 165157 8925 165169 8959
rect 165203 8956 165215 8959
rect 165246 8956 165252 8968
rect 165203 8928 165252 8956
rect 165203 8925 165215 8928
rect 165157 8919 165215 8925
rect 165246 8916 165252 8928
rect 165304 8916 165310 8968
rect 166644 8965 166672 8996
rect 177206 8984 177212 8996
rect 177264 8984 177270 9036
rect 179598 8984 179604 9036
rect 179656 8984 179662 9036
rect 180334 8984 180340 9036
rect 180392 9024 180398 9036
rect 180889 9027 180947 9033
rect 180889 9024 180901 9027
rect 180392 8996 180901 9024
rect 180392 8984 180398 8996
rect 180889 8993 180901 8996
rect 180935 8993 180947 9027
rect 180889 8987 180947 8993
rect 181806 8984 181812 9036
rect 181864 9024 181870 9036
rect 182177 9027 182235 9033
rect 182177 9024 182189 9027
rect 181864 8996 182189 9024
rect 181864 8984 181870 8996
rect 182177 8993 182189 8996
rect 182223 8993 182235 9027
rect 182177 8987 182235 8993
rect 182450 8984 182456 9036
rect 182508 8984 182514 9036
rect 184290 8984 184296 9036
rect 184348 8984 184354 9036
rect 166629 8959 166687 8965
rect 166629 8925 166641 8959
rect 166675 8925 166687 8959
rect 166629 8919 166687 8925
rect 167730 8916 167736 8968
rect 167788 8956 167794 8968
rect 167917 8959 167975 8965
rect 167917 8956 167929 8959
rect 167788 8928 167929 8956
rect 167788 8916 167794 8928
rect 167917 8925 167929 8928
rect 167963 8925 167975 8959
rect 167917 8919 167975 8925
rect 168098 8916 168104 8968
rect 168156 8916 168162 8968
rect 168282 8916 168288 8968
rect 168340 8956 168346 8968
rect 169021 8959 169079 8965
rect 168340 8928 168512 8956
rect 168340 8916 168346 8928
rect 166258 8848 166264 8900
rect 166316 8888 166322 8900
rect 167273 8891 167331 8897
rect 167273 8888 167285 8891
rect 166316 8860 167285 8888
rect 166316 8848 166322 8860
rect 167273 8857 167285 8860
rect 167319 8857 167331 8891
rect 167273 8851 167331 8857
rect 167362 8848 167368 8900
rect 167420 8888 167426 8900
rect 168484 8888 168512 8928
rect 169021 8925 169033 8959
rect 169067 8956 169079 8959
rect 169846 8956 169852 8968
rect 169067 8928 169852 8956
rect 169067 8925 169079 8928
rect 169021 8919 169079 8925
rect 169846 8916 169852 8928
rect 169904 8916 169910 8968
rect 169938 8916 169944 8968
rect 169996 8956 170002 8968
rect 170309 8959 170367 8965
rect 170309 8956 170321 8959
rect 169996 8928 170321 8956
rect 169996 8916 170002 8928
rect 170309 8925 170321 8928
rect 170355 8925 170367 8959
rect 170309 8919 170367 8925
rect 173710 8916 173716 8968
rect 173768 8956 173774 8968
rect 174081 8959 174139 8965
rect 174081 8956 174093 8959
rect 173768 8928 174093 8956
rect 173768 8916 173774 8928
rect 174081 8925 174093 8928
rect 174127 8925 174139 8959
rect 174081 8919 174139 8925
rect 176626 8928 176884 8956
rect 169665 8891 169723 8897
rect 169665 8888 169677 8891
rect 167420 8860 168420 8888
rect 168484 8860 169677 8888
rect 167420 8848 167426 8860
rect 167546 8820 167552 8832
rect 164804 8792 167552 8820
rect 167546 8780 167552 8792
rect 167604 8780 167610 8832
rect 167638 8780 167644 8832
rect 167696 8820 167702 8832
rect 168285 8823 168343 8829
rect 168285 8820 168297 8823
rect 167696 8792 168297 8820
rect 167696 8780 167702 8792
rect 168285 8789 168297 8792
rect 168331 8789 168343 8823
rect 168392 8820 168420 8860
rect 169665 8857 169677 8860
rect 169711 8857 169723 8891
rect 176626 8888 176654 8928
rect 169665 8851 169723 8857
rect 169772 8860 176654 8888
rect 169772 8820 169800 8860
rect 176746 8848 176752 8900
rect 176804 8848 176810 8900
rect 176856 8888 176884 8928
rect 177482 8916 177488 8968
rect 177540 8916 177546 8968
rect 179874 8916 179880 8968
rect 179932 8916 179938 8968
rect 181162 8916 181168 8968
rect 181220 8916 181226 8968
rect 184566 8916 184572 8968
rect 184624 8916 184630 8968
rect 184676 8888 184704 9064
rect 197170 9052 197176 9064
rect 197228 9052 197234 9104
rect 198090 9052 198096 9104
rect 198148 9092 198154 9104
rect 200114 9092 200120 9104
rect 198148 9064 200120 9092
rect 198148 9052 198154 9064
rect 200114 9052 200120 9064
rect 200172 9052 200178 9104
rect 201972 9092 202000 9132
rect 200592 9064 202000 9092
rect 184750 8984 184756 9036
rect 184808 9024 184814 9036
rect 185581 9027 185639 9033
rect 185581 9024 185593 9027
rect 184808 8996 185593 9024
rect 184808 8984 184814 8996
rect 185581 8993 185593 8996
rect 185627 8993 185639 9027
rect 185581 8987 185639 8993
rect 186222 8984 186228 9036
rect 186280 9024 186286 9036
rect 186869 9027 186927 9033
rect 186869 9024 186881 9027
rect 186280 8996 186881 9024
rect 186280 8984 186286 8996
rect 186869 8993 186881 8996
rect 186915 8993 186927 9027
rect 186869 8987 186927 8993
rect 189442 8984 189448 9036
rect 189500 8984 189506 9036
rect 190822 8984 190828 9036
rect 190880 9024 190886 9036
rect 197265 9027 197323 9033
rect 197265 9024 197277 9027
rect 190880 8996 197277 9024
rect 190880 8984 190886 8996
rect 197265 8993 197277 8996
rect 197311 8993 197323 9027
rect 197265 8987 197323 8993
rect 197556 8996 199976 9024
rect 185854 8916 185860 8968
rect 185912 8916 185918 8968
rect 187145 8959 187203 8965
rect 187145 8925 187157 8959
rect 187191 8925 187203 8959
rect 187145 8919 187203 8925
rect 176856 8860 184704 8888
rect 168392 8792 169800 8820
rect 168285 8783 168343 8789
rect 169846 8780 169852 8832
rect 169904 8820 169910 8832
rect 170217 8823 170275 8829
rect 170217 8820 170229 8823
rect 169904 8792 170229 8820
rect 169904 8780 169910 8792
rect 170217 8789 170229 8792
rect 170263 8820 170275 8823
rect 170306 8820 170312 8832
rect 170263 8792 170312 8820
rect 170263 8789 170275 8792
rect 170217 8783 170275 8789
rect 170306 8780 170312 8792
rect 170364 8780 170370 8832
rect 174170 8780 174176 8832
rect 174228 8780 174234 8832
rect 176838 8780 176844 8832
rect 176896 8780 176902 8832
rect 177574 8780 177580 8832
rect 177632 8780 177638 8832
rect 177850 8780 177856 8832
rect 177908 8820 177914 8832
rect 187160 8820 187188 8919
rect 187234 8916 187240 8968
rect 187292 8956 187298 8968
rect 189721 8959 189779 8965
rect 189721 8956 189733 8959
rect 187292 8928 189733 8956
rect 187292 8916 187298 8928
rect 189721 8925 189733 8928
rect 189767 8925 189779 8959
rect 189721 8919 189779 8925
rect 190641 8959 190699 8965
rect 190641 8925 190653 8959
rect 190687 8925 190699 8959
rect 190641 8919 190699 8925
rect 190733 8959 190791 8965
rect 190733 8925 190745 8959
rect 190779 8956 190791 8959
rect 190914 8956 190920 8968
rect 190779 8928 190920 8956
rect 190779 8925 190791 8928
rect 190733 8919 190791 8925
rect 190656 8888 190684 8919
rect 190914 8916 190920 8928
rect 190972 8956 190978 8968
rect 190972 8928 191144 8956
rect 190972 8916 190978 8928
rect 190822 8888 190828 8900
rect 190656 8860 190828 8888
rect 190822 8848 190828 8860
rect 190880 8848 190886 8900
rect 191116 8888 191144 8928
rect 191190 8916 191196 8968
rect 191248 8956 191254 8968
rect 191561 8959 191619 8965
rect 191561 8956 191573 8959
rect 191248 8928 191573 8956
rect 191248 8916 191254 8928
rect 191561 8925 191573 8928
rect 191607 8925 191619 8959
rect 191561 8919 191619 8925
rect 191745 8959 191803 8965
rect 191745 8925 191757 8959
rect 191791 8925 191803 8959
rect 191745 8919 191803 8925
rect 191760 8888 191788 8919
rect 192478 8916 192484 8968
rect 192536 8916 192542 8968
rect 192573 8959 192631 8965
rect 192573 8925 192585 8959
rect 192619 8925 192631 8959
rect 192573 8919 192631 8925
rect 192588 8888 192616 8919
rect 193306 8916 193312 8968
rect 193364 8916 193370 8968
rect 193401 8959 193459 8965
rect 193401 8925 193413 8959
rect 193447 8956 193459 8959
rect 193447 8928 193536 8956
rect 193447 8925 193459 8928
rect 193401 8919 193459 8925
rect 193508 8900 193536 8928
rect 194594 8916 194600 8968
rect 194652 8916 194658 8968
rect 194781 8959 194839 8965
rect 194781 8925 194793 8959
rect 194827 8925 194839 8959
rect 194781 8919 194839 8925
rect 193490 8888 193496 8900
rect 191116 8860 193496 8888
rect 193490 8848 193496 8860
rect 193548 8888 193554 8900
rect 194796 8888 194824 8919
rect 195514 8916 195520 8968
rect 195572 8916 195578 8968
rect 195609 8959 195667 8965
rect 195609 8925 195621 8959
rect 195655 8925 195667 8959
rect 195609 8919 195667 8925
rect 195624 8888 195652 8919
rect 196250 8916 196256 8968
rect 196308 8916 196314 8968
rect 196437 8959 196495 8965
rect 196437 8925 196449 8959
rect 196483 8956 196495 8959
rect 196526 8956 196532 8968
rect 196483 8928 196532 8956
rect 196483 8925 196495 8928
rect 196437 8919 196495 8925
rect 196452 8888 196480 8919
rect 196526 8916 196532 8928
rect 196584 8916 196590 8968
rect 197354 8916 197360 8968
rect 197412 8956 197418 8968
rect 197556 8965 197584 8996
rect 197541 8959 197599 8965
rect 197541 8956 197553 8959
rect 197412 8928 197553 8956
rect 197412 8916 197418 8928
rect 197541 8925 197553 8928
rect 197587 8925 197599 8959
rect 197541 8919 197599 8925
rect 197998 8916 198004 8968
rect 198056 8956 198062 8968
rect 198642 8956 198648 8968
rect 198056 8928 198648 8956
rect 198056 8916 198062 8928
rect 198642 8916 198648 8928
rect 198700 8916 198706 8968
rect 198752 8965 198780 8996
rect 198737 8959 198795 8965
rect 198737 8925 198749 8959
rect 198783 8925 198795 8959
rect 198737 8919 198795 8925
rect 199654 8916 199660 8968
rect 199712 8956 199718 8968
rect 199948 8965 199976 8996
rect 199749 8959 199807 8965
rect 199749 8956 199761 8959
rect 199712 8928 199761 8956
rect 199712 8916 199718 8928
rect 199749 8925 199761 8928
rect 199795 8925 199807 8959
rect 199749 8919 199807 8925
rect 199933 8959 199991 8965
rect 199933 8925 199945 8959
rect 199979 8925 199991 8959
rect 199933 8919 199991 8925
rect 193548 8860 196480 8888
rect 199948 8888 199976 8919
rect 200482 8916 200488 8968
rect 200540 8956 200546 8968
rect 200592 8965 200620 9064
rect 202046 9052 202052 9104
rect 202104 9092 202110 9104
rect 203610 9092 203616 9104
rect 202104 9064 203616 9092
rect 202104 9052 202110 9064
rect 203610 9052 203616 9064
rect 203668 9052 203674 9104
rect 203720 9092 203748 9132
rect 204070 9120 204076 9172
rect 204128 9120 204134 9172
rect 225598 9160 225604 9172
rect 209746 9132 225604 9160
rect 209746 9092 209774 9132
rect 225598 9120 225604 9132
rect 225656 9120 225662 9172
rect 228358 9120 228364 9172
rect 228416 9120 228422 9172
rect 228450 9120 228456 9172
rect 228508 9160 228514 9172
rect 233786 9160 233792 9172
rect 228508 9132 233792 9160
rect 228508 9120 228514 9132
rect 233786 9120 233792 9132
rect 233844 9120 233850 9172
rect 234062 9120 234068 9172
rect 234120 9120 234126 9172
rect 234154 9120 234160 9172
rect 234212 9160 234218 9172
rect 234893 9163 234951 9169
rect 234893 9160 234905 9163
rect 234212 9132 234905 9160
rect 234212 9120 234218 9132
rect 234893 9129 234905 9132
rect 234939 9129 234951 9163
rect 234893 9123 234951 9129
rect 235994 9120 236000 9172
rect 236052 9160 236058 9172
rect 236825 9163 236883 9169
rect 236825 9160 236837 9163
rect 236052 9132 236837 9160
rect 236052 9120 236058 9132
rect 236825 9129 236837 9132
rect 236871 9129 236883 9163
rect 236825 9123 236883 9129
rect 237282 9120 237288 9172
rect 237340 9160 237346 9172
rect 237561 9163 237619 9169
rect 237561 9160 237573 9163
rect 237340 9132 237573 9160
rect 237340 9120 237346 9132
rect 237561 9129 237573 9132
rect 237607 9129 237619 9163
rect 237561 9123 237619 9129
rect 237926 9120 237932 9172
rect 237984 9160 237990 9172
rect 258810 9160 258816 9172
rect 237984 9132 258816 9160
rect 237984 9120 237990 9132
rect 258810 9120 258816 9132
rect 258868 9120 258874 9172
rect 260190 9120 260196 9172
rect 260248 9120 260254 9172
rect 260650 9120 260656 9172
rect 260708 9160 260714 9172
rect 261757 9163 261815 9169
rect 261757 9160 261769 9163
rect 260708 9132 261769 9160
rect 260708 9120 260714 9132
rect 261757 9129 261769 9132
rect 261803 9129 261815 9163
rect 261757 9123 261815 9129
rect 262950 9120 262956 9172
rect 263008 9160 263014 9172
rect 269071 9163 269129 9169
rect 269071 9160 269083 9163
rect 263008 9132 269083 9160
rect 263008 9120 263014 9132
rect 269071 9129 269083 9132
rect 269117 9129 269129 9163
rect 269071 9123 269129 9129
rect 203720 9064 209774 9092
rect 210050 9052 210056 9104
rect 210108 9092 210114 9104
rect 212166 9092 212172 9104
rect 210108 9064 212172 9092
rect 210108 9052 210114 9064
rect 212166 9052 212172 9064
rect 212224 9052 212230 9104
rect 212350 9052 212356 9104
rect 212408 9092 212414 9104
rect 214374 9092 214380 9104
rect 212408 9064 214380 9092
rect 212408 9052 212414 9064
rect 214374 9052 214380 9064
rect 214432 9052 214438 9104
rect 214558 9052 214564 9104
rect 214616 9092 214622 9104
rect 222194 9092 222200 9104
rect 214616 9064 222200 9092
rect 214616 9052 214622 9064
rect 222194 9052 222200 9064
rect 222252 9052 222258 9104
rect 223393 9095 223451 9101
rect 223393 9061 223405 9095
rect 223439 9092 223451 9095
rect 223482 9092 223488 9104
rect 223439 9064 223488 9092
rect 223439 9061 223451 9064
rect 223393 9055 223451 9061
rect 223482 9052 223488 9064
rect 223540 9052 223546 9104
rect 225874 9052 225880 9104
rect 225932 9092 225938 9104
rect 233326 9092 233332 9104
rect 225932 9064 233332 9092
rect 225932 9052 225938 9064
rect 233326 9052 233332 9064
rect 233384 9052 233390 9104
rect 233418 9052 233424 9104
rect 233476 9092 233482 9104
rect 253934 9092 253940 9104
rect 233476 9064 253940 9092
rect 233476 9052 233482 9064
rect 253934 9052 253940 9064
rect 253992 9052 253998 9104
rect 262030 9092 262036 9104
rect 254044 9064 262036 9092
rect 200666 8984 200672 9036
rect 200724 9024 200730 9036
rect 221918 9024 221924 9036
rect 200724 8996 221924 9024
rect 200724 8984 200730 8996
rect 221918 8984 221924 8996
rect 221976 8984 221982 9036
rect 224313 9027 224371 9033
rect 224313 9024 224325 9027
rect 223224 8996 224325 9024
rect 200577 8959 200635 8965
rect 200577 8956 200589 8959
rect 200540 8928 200589 8956
rect 200540 8916 200546 8928
rect 200577 8925 200589 8928
rect 200623 8925 200635 8959
rect 200577 8919 200635 8925
rect 200761 8959 200819 8965
rect 200761 8925 200773 8959
rect 200807 8925 200819 8959
rect 200761 8919 200819 8925
rect 200776 8888 200804 8919
rect 201126 8916 201132 8968
rect 201184 8956 201190 8968
rect 201405 8959 201463 8965
rect 201405 8956 201417 8959
rect 201184 8928 201417 8956
rect 201184 8916 201190 8928
rect 201405 8925 201417 8928
rect 201451 8925 201463 8959
rect 201405 8919 201463 8925
rect 201589 8959 201647 8965
rect 201589 8925 201601 8959
rect 201635 8925 201647 8959
rect 201589 8919 201647 8925
rect 201604 8888 201632 8919
rect 202046 8916 202052 8968
rect 202104 8916 202110 8968
rect 202233 8959 202291 8965
rect 202233 8925 202245 8959
rect 202279 8925 202291 8959
rect 202233 8919 202291 8925
rect 202248 8888 202276 8919
rect 202598 8916 202604 8968
rect 202656 8956 202662 8968
rect 203061 8959 203119 8965
rect 203061 8956 203073 8959
rect 202656 8928 203073 8956
rect 202656 8916 202662 8928
rect 203061 8925 203073 8928
rect 203107 8925 203119 8959
rect 203061 8919 203119 8925
rect 203245 8959 203303 8965
rect 203245 8925 203257 8959
rect 203291 8925 203303 8959
rect 203245 8919 203303 8925
rect 202506 8888 202512 8900
rect 199948 8860 202512 8888
rect 193548 8848 193554 8860
rect 202506 8848 202512 8860
rect 202564 8888 202570 8900
rect 203260 8888 203288 8919
rect 203426 8916 203432 8968
rect 203484 8916 203490 8968
rect 203518 8916 203524 8968
rect 203576 8956 203582 8968
rect 203889 8959 203947 8965
rect 203889 8956 203901 8959
rect 203576 8928 203901 8956
rect 203576 8916 203582 8928
rect 203889 8925 203901 8928
rect 203935 8925 203947 8959
rect 203889 8919 203947 8925
rect 211706 8916 211712 8968
rect 211764 8916 211770 8968
rect 213914 8916 213920 8968
rect 213972 8956 213978 8968
rect 215662 8956 215668 8968
rect 213972 8928 215668 8956
rect 213972 8916 213978 8928
rect 215662 8916 215668 8928
rect 215720 8916 215726 8968
rect 216858 8916 216864 8968
rect 216916 8916 216922 8968
rect 222010 8916 222016 8968
rect 222068 8916 222074 8968
rect 223224 8965 223252 8996
rect 224313 8993 224325 8996
rect 224359 8993 224371 9027
rect 224313 8987 224371 8993
rect 224402 8984 224408 9036
rect 224460 9024 224466 9036
rect 225966 9024 225972 9036
rect 224460 8996 225644 9024
rect 224460 8984 224466 8996
rect 225616 8968 225644 8996
rect 225800 8996 225972 9024
rect 223209 8959 223267 8965
rect 223209 8925 223221 8959
rect 223255 8925 223267 8959
rect 223209 8919 223267 8925
rect 224034 8916 224040 8968
rect 224092 8916 224098 8968
rect 224129 8959 224187 8965
rect 224129 8925 224141 8959
rect 224175 8956 224187 8959
rect 224678 8956 224684 8968
rect 224175 8928 224684 8956
rect 224175 8925 224187 8928
rect 224129 8919 224187 8925
rect 224678 8916 224684 8928
rect 224736 8916 224742 8968
rect 225598 8916 225604 8968
rect 225656 8916 225662 8968
rect 225693 8959 225751 8965
rect 225693 8925 225705 8959
rect 225739 8956 225751 8959
rect 225800 8956 225828 8996
rect 225966 8984 225972 8996
rect 226024 9024 226030 9036
rect 226024 8996 229876 9024
rect 226024 8984 226030 8996
rect 225739 8928 225828 8956
rect 225739 8925 225751 8928
rect 225693 8919 225751 8925
rect 226426 8916 226432 8968
rect 226484 8916 226490 8968
rect 226536 8965 226564 8996
rect 226521 8959 226579 8965
rect 226521 8925 226533 8959
rect 226567 8925 226579 8959
rect 226521 8919 226579 8925
rect 227254 8916 227260 8968
rect 227312 8916 227318 8968
rect 227364 8965 227392 8996
rect 227349 8959 227407 8965
rect 227349 8925 227361 8959
rect 227395 8925 227407 8959
rect 227349 8919 227407 8925
rect 228082 8916 228088 8968
rect 228140 8916 228146 8968
rect 228192 8965 228220 8996
rect 228177 8959 228235 8965
rect 228177 8925 228189 8959
rect 228223 8925 228235 8959
rect 228177 8919 228235 8925
rect 228818 8916 228824 8968
rect 228876 8916 228882 8968
rect 229020 8965 229048 8996
rect 229848 8968 229876 8996
rect 230014 8984 230020 9036
rect 230072 8984 230078 9036
rect 230842 8984 230848 9036
rect 230900 9024 230906 9036
rect 231029 9027 231087 9033
rect 231029 9024 231041 9027
rect 230900 8996 231041 9024
rect 230900 8984 230906 8996
rect 231029 8993 231041 8996
rect 231075 9024 231087 9027
rect 231075 8996 235948 9024
rect 231075 8993 231087 8996
rect 231029 8987 231087 8993
rect 229005 8959 229063 8965
rect 229005 8925 229017 8959
rect 229051 8925 229063 8959
rect 229005 8919 229063 8925
rect 229094 8916 229100 8968
rect 229152 8956 229158 8968
rect 229646 8956 229652 8968
rect 229152 8928 229652 8956
rect 229152 8916 229158 8928
rect 229646 8916 229652 8928
rect 229704 8916 229710 8968
rect 229830 8916 229836 8968
rect 229888 8916 229894 8968
rect 230198 8916 230204 8968
rect 230256 8956 230262 8968
rect 230753 8959 230811 8965
rect 230753 8956 230765 8959
rect 230256 8928 230765 8956
rect 230256 8916 230262 8928
rect 230753 8925 230765 8928
rect 230799 8925 230811 8959
rect 230753 8919 230811 8925
rect 231854 8916 231860 8968
rect 231912 8956 231918 8968
rect 232041 8959 232099 8965
rect 232041 8956 232053 8959
rect 231912 8928 232053 8956
rect 231912 8916 231918 8928
rect 232041 8925 232053 8928
rect 232087 8956 232099 8959
rect 232130 8956 232136 8968
rect 232087 8928 232136 8956
rect 232087 8925 232099 8928
rect 232041 8919 232099 8925
rect 232130 8916 232136 8928
rect 232188 8916 232194 8968
rect 232240 8965 232268 8996
rect 232225 8959 232283 8965
rect 232225 8925 232237 8959
rect 232271 8925 232283 8959
rect 232225 8919 232283 8925
rect 232498 8916 232504 8968
rect 232556 8956 232562 8968
rect 232866 8956 232872 8968
rect 232556 8928 232872 8956
rect 232556 8916 232562 8928
rect 232866 8916 232872 8928
rect 232924 8916 232930 8968
rect 233068 8965 233096 8996
rect 233053 8959 233111 8965
rect 233053 8925 233065 8959
rect 233099 8925 233111 8959
rect 233053 8919 233111 8925
rect 233694 8916 233700 8968
rect 233752 8916 233758 8968
rect 233896 8965 233924 8996
rect 233881 8959 233939 8965
rect 233881 8925 233893 8959
rect 233927 8925 233939 8959
rect 233881 8919 233939 8925
rect 234522 8916 234528 8968
rect 234580 8916 234586 8968
rect 234724 8965 234752 8996
rect 235920 8968 235948 8996
rect 236086 8984 236092 9036
rect 236144 9024 236150 9036
rect 236144 8996 237420 9024
rect 236144 8984 236150 8996
rect 234709 8959 234767 8965
rect 234709 8925 234721 8959
rect 234755 8925 234767 8959
rect 235626 8956 235632 8968
rect 234709 8919 234767 8925
rect 235000 8928 235632 8956
rect 212350 8888 212356 8900
rect 202564 8860 203288 8888
rect 203536 8860 212356 8888
rect 202564 8848 202570 8860
rect 177908 8792 187188 8820
rect 177908 8780 177914 8792
rect 190362 8780 190368 8832
rect 190420 8820 190426 8832
rect 190917 8823 190975 8829
rect 190917 8820 190929 8823
rect 190420 8792 190929 8820
rect 190420 8780 190426 8792
rect 190917 8789 190929 8792
rect 190963 8789 190975 8823
rect 190917 8783 190975 8789
rect 191098 8780 191104 8832
rect 191156 8820 191162 8832
rect 191193 8823 191251 8829
rect 191193 8820 191205 8823
rect 191156 8792 191205 8820
rect 191156 8780 191162 8792
rect 191193 8789 191205 8792
rect 191239 8789 191251 8823
rect 191193 8783 191251 8789
rect 191926 8780 191932 8832
rect 191984 8780 191990 8832
rect 192018 8780 192024 8832
rect 192076 8820 192082 8832
rect 192757 8823 192815 8829
rect 192757 8820 192769 8823
rect 192076 8792 192769 8820
rect 192076 8780 192082 8792
rect 192757 8789 192769 8792
rect 192803 8789 192815 8823
rect 192757 8783 192815 8789
rect 194042 8780 194048 8832
rect 194100 8820 194106 8832
rect 194965 8823 195023 8829
rect 194965 8820 194977 8823
rect 194100 8792 194977 8820
rect 194100 8780 194106 8792
rect 194965 8789 194977 8792
rect 195011 8789 195023 8823
rect 194965 8783 195023 8789
rect 196342 8780 196348 8832
rect 196400 8820 196406 8832
rect 196621 8823 196679 8829
rect 196621 8820 196633 8823
rect 196400 8792 196633 8820
rect 196400 8780 196406 8792
rect 196621 8789 196633 8792
rect 196667 8789 196679 8823
rect 196621 8783 196679 8789
rect 199286 8780 199292 8832
rect 199344 8820 199350 8832
rect 200117 8823 200175 8829
rect 200117 8820 200129 8823
rect 199344 8792 200129 8820
rect 199344 8780 199350 8792
rect 200117 8789 200129 8792
rect 200163 8789 200175 8823
rect 200117 8783 200175 8789
rect 201034 8780 201040 8832
rect 201092 8820 201098 8832
rect 201773 8823 201831 8829
rect 201773 8820 201785 8823
rect 201092 8792 201785 8820
rect 201092 8780 201098 8792
rect 201773 8789 201785 8792
rect 201819 8789 201831 8823
rect 201773 8783 201831 8789
rect 202414 8780 202420 8832
rect 202472 8780 202478 8832
rect 202598 8780 202604 8832
rect 202656 8820 202662 8832
rect 202693 8823 202751 8829
rect 202693 8820 202705 8823
rect 202656 8792 202705 8820
rect 202656 8780 202662 8792
rect 202693 8789 202705 8792
rect 202739 8820 202751 8823
rect 203536 8820 203564 8860
rect 212350 8848 212356 8860
rect 212408 8848 212414 8900
rect 212442 8848 212448 8900
rect 212500 8888 212506 8900
rect 235000 8888 235028 8928
rect 235626 8916 235632 8928
rect 235684 8916 235690 8968
rect 235810 8916 235816 8968
rect 235868 8916 235874 8968
rect 235902 8916 235908 8968
rect 235960 8956 235966 8968
rect 237392 8965 237420 8996
rect 241974 8984 241980 9036
rect 242032 8984 242038 9036
rect 243446 8984 243452 9036
rect 243504 8984 243510 9036
rect 243538 8984 243544 9036
rect 243596 9024 243602 9036
rect 254044 9024 254072 9064
rect 262030 9052 262036 9064
rect 262088 9052 262094 9104
rect 263870 9052 263876 9104
rect 263928 9092 263934 9104
rect 264698 9092 264704 9104
rect 263928 9064 264704 9092
rect 263928 9052 263934 9064
rect 264698 9052 264704 9064
rect 264756 9052 264762 9104
rect 264790 9052 264796 9104
rect 264848 9052 264854 9104
rect 267550 9052 267556 9104
rect 267608 9092 267614 9104
rect 268381 9095 268439 9101
rect 268381 9092 268393 9095
rect 267608 9064 268393 9092
rect 267608 9052 267614 9064
rect 268381 9061 268393 9064
rect 268427 9061 268439 9095
rect 268381 9055 268439 9061
rect 243596 8996 254072 9024
rect 243596 8984 243602 8996
rect 254118 8984 254124 9036
rect 254176 8984 254182 9036
rect 256418 8984 256424 9036
rect 256476 8984 256482 9036
rect 257706 8984 257712 9036
rect 257764 8984 257770 9036
rect 258166 8984 258172 9036
rect 258224 9024 258230 9036
rect 263965 9027 264023 9033
rect 258224 8996 263594 9024
rect 258224 8984 258230 8996
rect 235997 8959 236055 8965
rect 235997 8956 236009 8959
rect 235960 8928 236009 8956
rect 235960 8916 235966 8928
rect 235997 8925 236009 8928
rect 236043 8925 236055 8959
rect 235997 8919 236055 8925
rect 236181 8959 236239 8965
rect 236181 8925 236193 8959
rect 236227 8956 236239 8959
rect 236641 8959 236699 8965
rect 236227 8950 236500 8956
rect 236641 8950 236653 8959
rect 236227 8928 236653 8950
rect 236227 8925 236239 8928
rect 236181 8919 236239 8925
rect 236472 8925 236653 8928
rect 236687 8925 236699 8959
rect 236472 8922 236699 8925
rect 236641 8919 236699 8922
rect 237377 8959 237435 8965
rect 237377 8925 237389 8959
rect 237423 8925 237435 8959
rect 237377 8919 237435 8925
rect 238754 8916 238760 8968
rect 238812 8956 238818 8968
rect 242253 8959 242311 8965
rect 242253 8956 242265 8959
rect 238812 8928 242265 8956
rect 238812 8916 238818 8928
rect 242253 8925 242265 8928
rect 242299 8925 242311 8959
rect 242253 8919 242311 8925
rect 243722 8916 243728 8968
rect 243780 8916 243786 8968
rect 244182 8916 244188 8968
rect 244240 8956 244246 8968
rect 244737 8959 244795 8965
rect 244737 8956 244749 8959
rect 244240 8928 244749 8956
rect 244240 8916 244246 8928
rect 244737 8925 244749 8928
rect 244783 8925 244795 8959
rect 244737 8919 244795 8925
rect 245010 8916 245016 8968
rect 245068 8916 245074 8968
rect 246114 8916 246120 8968
rect 246172 8916 246178 8968
rect 246206 8916 246212 8968
rect 246264 8956 246270 8968
rect 246393 8959 246451 8965
rect 246393 8956 246405 8959
rect 246264 8928 246405 8956
rect 246264 8916 246270 8928
rect 246393 8925 246405 8928
rect 246439 8925 246451 8959
rect 246393 8919 246451 8925
rect 247402 8916 247408 8968
rect 247460 8916 247466 8968
rect 247681 8959 247739 8965
rect 247681 8925 247693 8959
rect 247727 8925 247739 8959
rect 247681 8919 247739 8925
rect 212500 8860 235028 8888
rect 235276 8860 244274 8888
rect 212500 8848 212506 8860
rect 202739 8792 203564 8820
rect 202739 8789 202751 8792
rect 202693 8783 202751 8789
rect 203610 8780 203616 8832
rect 203668 8820 203674 8832
rect 211062 8820 211068 8832
rect 203668 8792 211068 8820
rect 203668 8780 203674 8792
rect 211062 8780 211068 8792
rect 211120 8780 211126 8832
rect 211525 8823 211583 8829
rect 211525 8789 211537 8823
rect 211571 8820 211583 8823
rect 214374 8820 214380 8832
rect 211571 8792 214380 8820
rect 211571 8789 211583 8792
rect 211525 8783 211583 8789
rect 214374 8780 214380 8792
rect 214432 8780 214438 8832
rect 216674 8780 216680 8832
rect 216732 8780 216738 8832
rect 221826 8780 221832 8832
rect 221884 8780 221890 8832
rect 221918 8780 221924 8832
rect 221976 8820 221982 8832
rect 225690 8820 225696 8832
rect 221976 8792 225696 8820
rect 221976 8780 221982 8792
rect 225690 8780 225696 8792
rect 225748 8780 225754 8832
rect 225782 8780 225788 8832
rect 225840 8820 225846 8832
rect 225877 8823 225935 8829
rect 225877 8820 225889 8823
rect 225840 8792 225889 8820
rect 225840 8780 225846 8792
rect 225877 8789 225889 8792
rect 225923 8789 225935 8823
rect 225877 8783 225935 8789
rect 226518 8780 226524 8832
rect 226576 8820 226582 8832
rect 226705 8823 226763 8829
rect 226705 8820 226717 8823
rect 226576 8792 226717 8820
rect 226576 8780 226582 8792
rect 226705 8789 226717 8792
rect 226751 8789 226763 8823
rect 226705 8783 226763 8789
rect 227533 8823 227591 8829
rect 227533 8789 227545 8823
rect 227579 8820 227591 8823
rect 228082 8820 228088 8832
rect 227579 8792 228088 8820
rect 227579 8789 227591 8792
rect 227533 8783 227591 8789
rect 228082 8780 228088 8792
rect 228140 8780 228146 8832
rect 228910 8780 228916 8832
rect 228968 8820 228974 8832
rect 229189 8823 229247 8829
rect 229189 8820 229201 8823
rect 228968 8792 229201 8820
rect 228968 8780 228974 8792
rect 229189 8789 229201 8792
rect 229235 8789 229247 8823
rect 229189 8783 229247 8789
rect 231762 8780 231768 8832
rect 231820 8820 231826 8832
rect 232409 8823 232467 8829
rect 232409 8820 232421 8823
rect 231820 8792 232421 8820
rect 231820 8780 231826 8792
rect 232409 8789 232421 8792
rect 232455 8789 232467 8823
rect 232409 8783 232467 8789
rect 233234 8780 233240 8832
rect 233292 8780 233298 8832
rect 233326 8780 233332 8832
rect 233384 8820 233390 8832
rect 234062 8820 234068 8832
rect 233384 8792 234068 8820
rect 233384 8780 233390 8792
rect 234062 8780 234068 8792
rect 234120 8820 234126 8832
rect 234522 8820 234528 8832
rect 234120 8792 234528 8820
rect 234120 8780 234126 8792
rect 234522 8780 234528 8792
rect 234580 8820 234586 8832
rect 235276 8820 235304 8860
rect 234580 8792 235304 8820
rect 234580 8780 234586 8792
rect 235626 8780 235632 8832
rect 235684 8820 235690 8832
rect 236362 8820 236368 8832
rect 235684 8792 236368 8820
rect 235684 8780 235690 8792
rect 236362 8780 236368 8792
rect 236420 8780 236426 8832
rect 236546 8780 236552 8832
rect 236604 8780 236610 8832
rect 244246 8820 244274 8860
rect 246482 8848 246488 8900
rect 246540 8888 246546 8900
rect 247696 8888 247724 8919
rect 248690 8916 248696 8968
rect 248748 8916 248754 8968
rect 248969 8959 249027 8965
rect 248969 8925 248981 8959
rect 249015 8925 249027 8959
rect 248969 8919 249027 8925
rect 246540 8860 247724 8888
rect 246540 8848 246546 8860
rect 247770 8848 247776 8900
rect 247828 8888 247834 8900
rect 248984 8888 249012 8919
rect 250806 8916 250812 8968
rect 250864 8956 250870 8968
rect 251269 8959 251327 8965
rect 251269 8956 251281 8959
rect 250864 8928 251281 8956
rect 250864 8916 250870 8928
rect 251269 8925 251281 8928
rect 251315 8925 251327 8959
rect 251269 8919 251327 8925
rect 251358 8916 251364 8968
rect 251416 8956 251422 8968
rect 251545 8959 251603 8965
rect 251545 8956 251557 8959
rect 251416 8928 251557 8956
rect 251416 8916 251422 8928
rect 251545 8925 251557 8928
rect 251591 8925 251603 8959
rect 251545 8919 251603 8925
rect 252278 8916 252284 8968
rect 252336 8956 252342 8968
rect 252557 8959 252615 8965
rect 252557 8956 252569 8959
rect 252336 8928 252569 8956
rect 252336 8916 252342 8928
rect 252557 8925 252569 8928
rect 252603 8925 252615 8959
rect 252557 8919 252615 8925
rect 252830 8916 252836 8968
rect 252888 8916 252894 8968
rect 253842 8916 253848 8968
rect 253900 8916 253906 8968
rect 256697 8959 256755 8965
rect 256697 8925 256709 8959
rect 256743 8956 256755 8959
rect 256878 8956 256884 8968
rect 256743 8928 256884 8956
rect 256743 8925 256755 8928
rect 256697 8919 256755 8925
rect 256878 8916 256884 8928
rect 256936 8916 256942 8968
rect 257062 8916 257068 8968
rect 257120 8956 257126 8968
rect 257985 8959 258043 8965
rect 257985 8956 257997 8959
rect 257120 8928 257997 8956
rect 257120 8916 257126 8928
rect 257985 8925 257997 8928
rect 258031 8925 258043 8959
rect 257985 8919 258043 8925
rect 258350 8916 258356 8968
rect 258408 8956 258414 8968
rect 258408 8928 260236 8956
rect 258408 8916 258414 8928
rect 247828 8860 249012 8888
rect 247828 8848 247834 8860
rect 253934 8848 253940 8900
rect 253992 8888 253998 8900
rect 258718 8888 258724 8900
rect 253992 8860 258724 8888
rect 253992 8848 253998 8860
rect 258718 8848 258724 8860
rect 258776 8888 258782 8900
rect 258776 8860 259040 8888
rect 258776 8848 258782 8860
rect 258902 8820 258908 8832
rect 244246 8792 258908 8820
rect 258902 8780 258908 8792
rect 258960 8780 258966 8832
rect 259012 8820 259040 8860
rect 259086 8848 259092 8900
rect 259144 8848 259150 8900
rect 260098 8848 260104 8900
rect 260156 8848 260162 8900
rect 259181 8823 259239 8829
rect 259181 8820 259193 8823
rect 259012 8792 259193 8820
rect 259181 8789 259193 8792
rect 259227 8789 259239 8823
rect 260208 8820 260236 8928
rect 260374 8916 260380 8968
rect 260432 8956 260438 8968
rect 263566 8956 263594 8996
rect 263965 8993 263977 9027
rect 264011 9024 264023 9027
rect 265066 9024 265072 9036
rect 264011 8996 265072 9024
rect 264011 8993 264023 8996
rect 263965 8987 264023 8993
rect 265066 8984 265072 8996
rect 265124 8984 265130 9036
rect 265158 8984 265164 9036
rect 265216 9024 265222 9036
rect 267921 9027 267979 9033
rect 267921 9024 267933 9027
rect 265216 8996 267933 9024
rect 265216 8984 265222 8996
rect 267921 8993 267933 8996
rect 267967 8993 267979 9027
rect 267921 8987 267979 8993
rect 268841 9027 268899 9033
rect 268841 8993 268853 9027
rect 268887 9024 268899 9027
rect 270586 9024 270592 9036
rect 268887 8996 270592 9024
rect 268887 8993 268899 8996
rect 268841 8987 268899 8993
rect 270586 8984 270592 8996
rect 270644 8984 270650 9036
rect 263689 8959 263747 8965
rect 263689 8956 263701 8959
rect 260432 8928 262720 8956
rect 263566 8928 263701 8956
rect 260432 8916 260438 8928
rect 260650 8848 260656 8900
rect 260708 8888 260714 8900
rect 261665 8891 261723 8897
rect 261665 8888 261677 8891
rect 260708 8860 261677 8888
rect 260708 8848 260714 8860
rect 261665 8857 261677 8860
rect 261711 8857 261723 8891
rect 261665 8851 261723 8857
rect 262582 8848 262588 8900
rect 262640 8848 262646 8900
rect 262692 8888 262720 8928
rect 263689 8925 263701 8928
rect 263735 8925 263747 8959
rect 263689 8919 263747 8925
rect 263778 8916 263784 8968
rect 263836 8956 263842 8968
rect 265802 8956 265808 8968
rect 263836 8928 265808 8956
rect 263836 8916 263842 8928
rect 265802 8916 265808 8928
rect 265860 8916 265866 8968
rect 265986 8916 265992 8968
rect 266044 8956 266050 8968
rect 266044 8928 267412 8956
rect 266044 8916 266050 8928
rect 267384 8900 267412 8928
rect 267458 8916 267464 8968
rect 267516 8956 267522 8968
rect 268013 8959 268071 8965
rect 268013 8956 268025 8959
rect 267516 8928 268025 8956
rect 267516 8916 267522 8928
rect 268013 8925 268025 8928
rect 268059 8925 268071 8959
rect 268013 8919 268071 8925
rect 268286 8916 268292 8968
rect 268344 8956 268350 8968
rect 270129 8959 270187 8965
rect 268344 8928 269620 8956
rect 268344 8916 268350 8928
rect 265158 8888 265164 8900
rect 262692 8860 265164 8888
rect 265158 8848 265164 8860
rect 265216 8848 265222 8900
rect 265253 8891 265311 8897
rect 265253 8857 265265 8891
rect 265299 8857 265311 8891
rect 265253 8851 265311 8857
rect 261846 8820 261852 8832
rect 260208 8792 261852 8820
rect 259181 8783 259239 8789
rect 261846 8780 261852 8792
rect 261904 8820 261910 8832
rect 262677 8823 262735 8829
rect 262677 8820 262689 8823
rect 261904 8792 262689 8820
rect 261904 8780 261910 8792
rect 262677 8789 262689 8792
rect 262723 8789 262735 8823
rect 262677 8783 262735 8789
rect 264790 8780 264796 8832
rect 264848 8820 264854 8832
rect 265268 8820 265296 8851
rect 266814 8848 266820 8900
rect 266872 8888 266878 8900
rect 267182 8888 267188 8900
rect 266872 8860 267188 8888
rect 266872 8848 266878 8860
rect 267182 8848 267188 8860
rect 267240 8848 267246 8900
rect 267366 8848 267372 8900
rect 267424 8888 267430 8900
rect 269482 8888 269488 8900
rect 267424 8860 269488 8888
rect 267424 8848 267430 8860
rect 269482 8848 269488 8860
rect 269540 8848 269546 8900
rect 269592 8888 269620 8928
rect 270129 8925 270141 8959
rect 270175 8956 270187 8959
rect 270310 8956 270316 8968
rect 270175 8928 270316 8956
rect 270175 8925 270187 8928
rect 270129 8919 270187 8925
rect 270310 8916 270316 8928
rect 270368 8916 270374 8968
rect 270402 8916 270408 8968
rect 270460 8916 270466 8968
rect 270770 8888 270776 8900
rect 269592 8860 270776 8888
rect 270770 8848 270776 8860
rect 270828 8848 270834 8900
rect 264848 8792 265296 8820
rect 264848 8780 264854 8792
rect 265342 8780 265348 8832
rect 265400 8780 265406 8832
rect 266630 8780 266636 8832
rect 266688 8820 266694 8832
rect 266909 8823 266967 8829
rect 266909 8820 266921 8823
rect 266688 8792 266921 8820
rect 266688 8780 266694 8792
rect 266909 8789 266921 8792
rect 266955 8789 266967 8823
rect 266909 8783 266967 8789
rect 267734 8780 267740 8832
rect 267792 8820 267798 8832
rect 268562 8820 268568 8832
rect 267792 8792 268568 8820
rect 267792 8780 267798 8792
rect 268562 8780 268568 8792
rect 268620 8780 268626 8832
rect 269298 8780 269304 8832
rect 269356 8820 269362 8832
rect 271046 8820 271052 8832
rect 269356 8792 271052 8820
rect 269356 8780 269362 8792
rect 271046 8780 271052 8792
rect 271104 8780 271110 8832
rect 1104 8730 271651 8752
rect 1104 8678 68546 8730
rect 68598 8678 68610 8730
rect 68662 8678 68674 8730
rect 68726 8678 68738 8730
rect 68790 8678 68802 8730
rect 68854 8678 136143 8730
rect 136195 8678 136207 8730
rect 136259 8678 136271 8730
rect 136323 8678 136335 8730
rect 136387 8678 136399 8730
rect 136451 8678 203740 8730
rect 203792 8678 203804 8730
rect 203856 8678 203868 8730
rect 203920 8678 203932 8730
rect 203984 8678 203996 8730
rect 204048 8678 271337 8730
rect 271389 8678 271401 8730
rect 271453 8678 271465 8730
rect 271517 8678 271529 8730
rect 271581 8678 271593 8730
rect 271645 8678 271651 8730
rect 1104 8656 271651 8678
rect 6914 8576 6920 8628
rect 6972 8616 6978 8628
rect 23290 8616 23296 8628
rect 6972 8588 23296 8616
rect 6972 8576 6978 8588
rect 23290 8576 23296 8588
rect 23348 8576 23354 8628
rect 23474 8576 23480 8628
rect 23532 8576 23538 8628
rect 25225 8619 25283 8625
rect 25225 8585 25237 8619
rect 25271 8616 25283 8619
rect 25271 8588 27292 8616
rect 25271 8585 25283 8588
rect 25225 8579 25283 8585
rect 23106 8508 23112 8560
rect 23164 8548 23170 8560
rect 23164 8520 23980 8548
rect 23164 8508 23170 8520
rect 23293 8483 23351 8489
rect 23293 8449 23305 8483
rect 23339 8449 23351 8483
rect 23293 8443 23351 8449
rect 13538 8304 13544 8356
rect 13596 8344 13602 8356
rect 23198 8344 23204 8356
rect 13596 8316 23204 8344
rect 13596 8304 13602 8316
rect 23198 8304 23204 8316
rect 23256 8304 23262 8356
rect 23308 8344 23336 8443
rect 23750 8440 23756 8492
rect 23808 8480 23814 8492
rect 23845 8483 23903 8489
rect 23845 8480 23857 8483
rect 23808 8452 23857 8480
rect 23808 8440 23814 8452
rect 23845 8449 23857 8452
rect 23891 8449 23903 8483
rect 23845 8443 23903 8449
rect 23952 8412 23980 8520
rect 25682 8508 25688 8560
rect 25740 8548 25746 8560
rect 25777 8551 25835 8557
rect 25777 8548 25789 8551
rect 25740 8520 25789 8548
rect 25740 8508 25746 8520
rect 25777 8517 25789 8520
rect 25823 8517 25835 8551
rect 25777 8511 25835 8517
rect 25958 8508 25964 8560
rect 26016 8548 26022 8560
rect 26145 8551 26203 8557
rect 26145 8548 26157 8551
rect 26016 8520 26157 8548
rect 26016 8508 26022 8520
rect 26145 8517 26157 8520
rect 26191 8517 26203 8551
rect 26145 8511 26203 8517
rect 26234 8508 26240 8560
rect 26292 8548 26298 8560
rect 27264 8557 27292 8588
rect 28718 8576 28724 8628
rect 28776 8576 28782 8628
rect 29638 8576 29644 8628
rect 29696 8576 29702 8628
rect 30190 8576 30196 8628
rect 30248 8616 30254 8628
rect 30469 8619 30527 8625
rect 30469 8616 30481 8619
rect 30248 8588 30481 8616
rect 30248 8576 30254 8588
rect 30469 8585 30481 8588
rect 30515 8585 30527 8619
rect 30469 8579 30527 8585
rect 31294 8576 31300 8628
rect 31352 8576 31358 8628
rect 31938 8576 31944 8628
rect 31996 8616 32002 8628
rect 32582 8616 32588 8628
rect 31996 8588 32588 8616
rect 31996 8576 32002 8588
rect 32582 8576 32588 8588
rect 32640 8576 32646 8628
rect 32674 8576 32680 8628
rect 32732 8576 32738 8628
rect 54110 8576 54116 8628
rect 54168 8576 54174 8628
rect 54754 8576 54760 8628
rect 54812 8576 54818 8628
rect 55490 8576 55496 8628
rect 55548 8576 55554 8628
rect 56226 8576 56232 8628
rect 56284 8576 56290 8628
rect 57054 8576 57060 8628
rect 57112 8576 57118 8628
rect 58618 8576 58624 8628
rect 58676 8576 58682 8628
rect 59814 8576 59820 8628
rect 59872 8576 59878 8628
rect 60734 8576 60740 8628
rect 60792 8576 60798 8628
rect 61562 8576 61568 8628
rect 61620 8576 61626 8628
rect 62298 8576 62304 8628
rect 62356 8576 62362 8628
rect 63770 8576 63776 8628
rect 63828 8576 63834 8628
rect 64598 8576 64604 8628
rect 64656 8576 64662 8628
rect 64690 8576 64696 8628
rect 64748 8616 64754 8628
rect 64748 8588 84194 8616
rect 64748 8576 64754 8588
rect 27249 8551 27307 8557
rect 26292 8520 26464 8548
rect 26292 8508 26298 8520
rect 24026 8440 24032 8492
rect 24084 8440 24090 8492
rect 24136 8452 24992 8480
rect 24136 8412 24164 8452
rect 23952 8384 24164 8412
rect 24210 8372 24216 8424
rect 24268 8372 24274 8424
rect 24581 8415 24639 8421
rect 24581 8381 24593 8415
rect 24627 8412 24639 8415
rect 24854 8412 24860 8424
rect 24627 8384 24860 8412
rect 24627 8381 24639 8384
rect 24581 8375 24639 8381
rect 24854 8372 24860 8384
rect 24912 8372 24918 8424
rect 24964 8412 24992 8452
rect 25038 8440 25044 8492
rect 25096 8440 25102 8492
rect 26436 8489 26464 8520
rect 27249 8517 27261 8551
rect 27295 8517 27307 8551
rect 29730 8548 29736 8560
rect 27249 8511 27307 8517
rect 28184 8520 29736 8548
rect 26421 8483 26479 8489
rect 26421 8449 26433 8483
rect 26467 8449 26479 8483
rect 26421 8443 26479 8449
rect 26605 8483 26663 8489
rect 26605 8449 26617 8483
rect 26651 8480 26663 8483
rect 28184 8480 28212 8520
rect 29730 8508 29736 8520
rect 29788 8508 29794 8560
rect 36354 8548 36360 8560
rect 31726 8520 36360 8548
rect 26651 8452 28212 8480
rect 26651 8449 26663 8452
rect 26605 8443 26663 8449
rect 28442 8440 28448 8492
rect 28500 8440 28506 8492
rect 28537 8483 28595 8489
rect 28537 8449 28549 8483
rect 28583 8480 28595 8483
rect 28994 8480 29000 8492
rect 28583 8452 29000 8480
rect 28583 8449 28595 8452
rect 28537 8443 28595 8449
rect 28994 8440 29000 8452
rect 29052 8440 29058 8492
rect 29454 8440 29460 8492
rect 29512 8440 29518 8492
rect 30282 8440 30288 8492
rect 30340 8440 30346 8492
rect 31110 8440 31116 8492
rect 31168 8440 31174 8492
rect 24964 8384 25360 8412
rect 25222 8344 25228 8356
rect 23308 8316 25228 8344
rect 25222 8304 25228 8316
rect 25280 8304 25286 8356
rect 25332 8344 25360 8384
rect 25498 8372 25504 8424
rect 25556 8412 25562 8424
rect 25774 8412 25780 8424
rect 25556 8384 25780 8412
rect 25556 8372 25562 8384
rect 25774 8372 25780 8384
rect 25832 8412 25838 8424
rect 26237 8415 26295 8421
rect 26237 8412 26249 8415
rect 25832 8384 26249 8412
rect 25832 8372 25838 8384
rect 26237 8381 26249 8384
rect 26283 8381 26295 8415
rect 26237 8375 26295 8381
rect 31726 8344 31754 8520
rect 36354 8508 36360 8520
rect 36412 8508 36418 8560
rect 65702 8548 65708 8560
rect 41386 8520 65708 8548
rect 32490 8440 32496 8492
rect 32548 8440 32554 8492
rect 32582 8440 32588 8492
rect 32640 8480 32646 8492
rect 41386 8480 41414 8520
rect 65702 8508 65708 8520
rect 65760 8548 65766 8560
rect 65978 8548 65984 8560
rect 65760 8520 65984 8548
rect 65760 8508 65766 8520
rect 65978 8508 65984 8520
rect 66036 8508 66042 8560
rect 66990 8508 66996 8560
rect 67048 8508 67054 8560
rect 84166 8548 84194 8588
rect 88334 8576 88340 8628
rect 88392 8616 88398 8628
rect 88981 8619 89039 8625
rect 88981 8616 88993 8619
rect 88392 8588 88993 8616
rect 88392 8576 88398 8588
rect 88981 8585 88993 8588
rect 89027 8585 89039 8619
rect 88981 8579 89039 8585
rect 90450 8576 90456 8628
rect 90508 8616 90514 8628
rect 91097 8619 91155 8625
rect 91097 8616 91109 8619
rect 90508 8588 91109 8616
rect 90508 8576 90514 8588
rect 91097 8585 91109 8588
rect 91143 8585 91155 8619
rect 91097 8579 91155 8585
rect 91830 8576 91836 8628
rect 91888 8576 91894 8628
rect 91922 8576 91928 8628
rect 91980 8616 91986 8628
rect 92569 8619 92627 8625
rect 92569 8616 92581 8619
rect 91980 8588 92581 8616
rect 91980 8576 91986 8588
rect 92569 8585 92581 8588
rect 92615 8585 92627 8619
rect 92569 8579 92627 8585
rect 94590 8576 94596 8628
rect 94648 8576 94654 8628
rect 94866 8576 94872 8628
rect 94924 8616 94930 8628
rect 95329 8619 95387 8625
rect 95329 8616 95341 8619
rect 94924 8588 95341 8616
rect 94924 8576 94930 8588
rect 95329 8585 95341 8588
rect 95375 8585 95387 8619
rect 95329 8579 95387 8585
rect 96798 8576 96804 8628
rect 96856 8576 96862 8628
rect 97442 8576 97448 8628
rect 97500 8576 97506 8628
rect 98638 8576 98644 8628
rect 98696 8576 98702 8628
rect 100202 8576 100208 8628
rect 100260 8576 100266 8628
rect 100294 8576 100300 8628
rect 100352 8616 100358 8628
rect 100849 8619 100907 8625
rect 100849 8616 100861 8619
rect 100352 8588 100861 8616
rect 100352 8576 100358 8588
rect 100849 8585 100861 8588
rect 100895 8585 100907 8619
rect 100849 8579 100907 8585
rect 120810 8576 120816 8628
rect 120868 8616 120874 8628
rect 121917 8619 121975 8625
rect 121917 8616 121929 8619
rect 120868 8588 121929 8616
rect 120868 8576 120874 8588
rect 121917 8585 121929 8588
rect 121963 8585 121975 8619
rect 121917 8579 121975 8585
rect 123202 8576 123208 8628
rect 123260 8576 123266 8628
rect 123938 8576 123944 8628
rect 123996 8576 124002 8628
rect 125318 8576 125324 8628
rect 125376 8616 125382 8628
rect 125597 8619 125655 8625
rect 125597 8616 125609 8619
rect 125376 8588 125609 8616
rect 125376 8576 125382 8588
rect 125597 8585 125609 8588
rect 125643 8585 125655 8619
rect 125597 8579 125655 8585
rect 126330 8576 126336 8628
rect 126388 8576 126394 8628
rect 126790 8576 126796 8628
rect 126848 8616 126854 8628
rect 127069 8619 127127 8625
rect 127069 8616 127081 8619
rect 126848 8588 127081 8616
rect 126848 8576 126854 8588
rect 127069 8585 127081 8588
rect 127115 8585 127127 8619
rect 127069 8579 127127 8585
rect 127986 8576 127992 8628
rect 128044 8576 128050 8628
rect 128630 8576 128636 8628
rect 128688 8616 128694 8628
rect 129461 8619 129519 8625
rect 129461 8616 129473 8619
rect 128688 8588 129473 8616
rect 128688 8576 128694 8588
rect 129461 8585 129473 8588
rect 129507 8585 129519 8619
rect 129461 8579 129519 8585
rect 130470 8576 130476 8628
rect 130528 8616 130534 8628
rect 131577 8619 131635 8625
rect 131577 8616 131589 8619
rect 130528 8588 131589 8616
rect 130528 8576 130534 8588
rect 131577 8585 131589 8588
rect 131623 8585 131635 8619
rect 131577 8579 131635 8585
rect 132310 8576 132316 8628
rect 132368 8576 132374 8628
rect 134518 8576 134524 8628
rect 134576 8576 134582 8628
rect 137278 8576 137284 8628
rect 137336 8616 137342 8628
rect 156877 8619 156935 8625
rect 137336 8588 149100 8616
rect 137336 8576 137342 8588
rect 89990 8548 89996 8560
rect 84166 8520 89996 8548
rect 89990 8508 89996 8520
rect 90048 8548 90054 8560
rect 90726 8548 90732 8560
rect 90048 8520 90732 8548
rect 90048 8508 90054 8520
rect 90726 8508 90732 8520
rect 90784 8548 90790 8560
rect 124122 8548 124128 8560
rect 90784 8520 124128 8548
rect 90784 8508 90790 8520
rect 124122 8508 124128 8520
rect 124180 8508 124186 8560
rect 125870 8508 125876 8560
rect 125928 8548 125934 8560
rect 128722 8548 128728 8560
rect 125928 8520 128728 8548
rect 125928 8508 125934 8520
rect 128722 8508 128728 8520
rect 128780 8508 128786 8560
rect 149072 8548 149100 8588
rect 156877 8585 156889 8619
rect 156923 8616 156935 8619
rect 157426 8616 157432 8628
rect 156923 8588 157432 8616
rect 156923 8585 156935 8588
rect 156877 8579 156935 8585
rect 157426 8576 157432 8588
rect 157484 8576 157490 8628
rect 158349 8619 158407 8625
rect 158349 8585 158361 8619
rect 158395 8616 158407 8619
rect 159266 8616 159272 8628
rect 158395 8588 159272 8616
rect 158395 8585 158407 8588
rect 158349 8579 158407 8585
rect 159266 8576 159272 8588
rect 159324 8576 159330 8628
rect 159358 8576 159364 8628
rect 159416 8576 159422 8628
rect 159818 8576 159824 8628
rect 159876 8616 159882 8628
rect 161198 8616 161204 8628
rect 159876 8588 161204 8616
rect 159876 8576 159882 8588
rect 161198 8576 161204 8588
rect 161256 8576 161262 8628
rect 161860 8588 164234 8616
rect 159836 8548 159864 8576
rect 128832 8520 138014 8548
rect 149072 8520 159864 8548
rect 32640 8452 41414 8480
rect 53929 8483 53987 8489
rect 32640 8440 32646 8452
rect 53929 8449 53941 8483
rect 53975 8480 53987 8483
rect 54018 8480 54024 8492
rect 53975 8452 54024 8480
rect 53975 8449 53987 8452
rect 53929 8443 53987 8449
rect 54018 8440 54024 8452
rect 54076 8440 54082 8492
rect 54570 8440 54576 8492
rect 54628 8440 54634 8492
rect 55306 8440 55312 8492
rect 55364 8440 55370 8492
rect 56042 8440 56048 8492
rect 56100 8440 56106 8492
rect 56870 8440 56876 8492
rect 56928 8440 56934 8492
rect 58434 8440 58440 8492
rect 58492 8440 58498 8492
rect 59725 8483 59783 8489
rect 59725 8449 59737 8483
rect 59771 8480 59783 8483
rect 60553 8483 60611 8489
rect 59771 8452 60504 8480
rect 59771 8449 59783 8452
rect 59725 8443 59783 8449
rect 32309 8415 32367 8421
rect 32309 8381 32321 8415
rect 32355 8412 32367 8415
rect 33137 8415 33195 8421
rect 33137 8412 33149 8415
rect 32355 8384 33149 8412
rect 32355 8381 32367 8384
rect 32309 8375 32367 8381
rect 33137 8381 33149 8384
rect 33183 8381 33195 8415
rect 33137 8375 33195 8381
rect 53745 8415 53803 8421
rect 53745 8381 53757 8415
rect 53791 8412 53803 8415
rect 54110 8412 54116 8424
rect 53791 8384 54116 8412
rect 53791 8381 53803 8384
rect 53745 8375 53803 8381
rect 54110 8372 54116 8384
rect 54168 8372 54174 8424
rect 60366 8372 60372 8424
rect 60424 8372 60430 8424
rect 60476 8412 60504 8452
rect 60553 8449 60565 8483
rect 60599 8480 60611 8483
rect 60918 8480 60924 8492
rect 60599 8452 60924 8480
rect 60599 8449 60611 8452
rect 60553 8443 60611 8449
rect 60918 8440 60924 8452
rect 60976 8440 60982 8492
rect 61378 8440 61384 8492
rect 61436 8440 61442 8492
rect 62114 8440 62120 8492
rect 62172 8440 62178 8492
rect 63586 8440 63592 8492
rect 63644 8440 63650 8492
rect 64414 8440 64420 8492
rect 64472 8440 64478 8492
rect 65242 8440 65248 8492
rect 65300 8440 65306 8492
rect 66806 8440 66812 8492
rect 66864 8440 66870 8492
rect 71314 8440 71320 8492
rect 71372 8440 71378 8492
rect 74258 8440 74264 8492
rect 74316 8440 74322 8492
rect 76466 8440 76472 8492
rect 76524 8440 76530 8492
rect 76742 8440 76748 8492
rect 76800 8440 76806 8492
rect 79410 8440 79416 8492
rect 79468 8440 79474 8492
rect 81618 8440 81624 8492
rect 81676 8440 81682 8492
rect 88794 8440 88800 8492
rect 88852 8440 88858 8492
rect 89162 8440 89168 8492
rect 89220 8480 89226 8492
rect 89901 8483 89959 8489
rect 89901 8480 89913 8483
rect 89220 8452 89913 8480
rect 89220 8440 89226 8452
rect 89901 8449 89913 8452
rect 89947 8449 89959 8483
rect 89901 8443 89959 8449
rect 90910 8440 90916 8492
rect 90968 8440 90974 8492
rect 91646 8440 91652 8492
rect 91704 8440 91710 8492
rect 92382 8440 92388 8492
rect 92440 8440 92446 8492
rect 93210 8440 93216 8492
rect 93268 8440 93274 8492
rect 93305 8483 93363 8489
rect 93305 8449 93317 8483
rect 93351 8480 93363 8483
rect 93486 8480 93492 8492
rect 93351 8452 93492 8480
rect 93351 8449 93363 8452
rect 93305 8443 93363 8449
rect 93486 8440 93492 8452
rect 93544 8440 93550 8492
rect 94406 8440 94412 8492
rect 94464 8440 94470 8492
rect 95142 8440 95148 8492
rect 95200 8440 95206 8492
rect 95970 8440 95976 8492
rect 96028 8480 96034 8492
rect 96430 8480 96436 8492
rect 96028 8452 96436 8480
rect 96028 8440 96034 8452
rect 96430 8440 96436 8452
rect 96488 8440 96494 8492
rect 96614 8440 96620 8492
rect 96672 8440 96678 8492
rect 97258 8440 97264 8492
rect 97316 8440 97322 8492
rect 98454 8440 98460 8492
rect 98512 8440 98518 8492
rect 99926 8440 99932 8492
rect 99984 8440 99990 8492
rect 100018 8440 100024 8492
rect 100076 8440 100082 8492
rect 100662 8440 100668 8492
rect 100720 8440 100726 8492
rect 111702 8440 111708 8492
rect 111760 8480 111766 8492
rect 121270 8480 121276 8492
rect 111760 8452 121276 8480
rect 111760 8440 111766 8452
rect 121270 8440 121276 8452
rect 121328 8480 121334 8492
rect 121549 8483 121607 8489
rect 121549 8480 121561 8483
rect 121328 8452 121561 8480
rect 121328 8440 121334 8452
rect 121549 8449 121561 8452
rect 121595 8449 121607 8483
rect 121549 8443 121607 8449
rect 121730 8440 121736 8492
rect 121788 8440 121794 8492
rect 123018 8440 123024 8492
rect 123076 8440 123082 8492
rect 123754 8440 123760 8492
rect 123812 8440 123818 8492
rect 125410 8440 125416 8492
rect 125468 8440 125474 8492
rect 126146 8440 126152 8492
rect 126204 8440 126210 8492
rect 126882 8440 126888 8492
rect 126940 8440 126946 8492
rect 127618 8440 127624 8492
rect 127676 8440 127682 8492
rect 127802 8440 127808 8492
rect 127860 8440 127866 8492
rect 66625 8415 66683 8421
rect 60476 8384 66392 8412
rect 25332 8316 31754 8344
rect 32600 8316 32812 8344
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 26878 8276 26884 8288
rect 3476 8248 26884 8276
rect 3476 8236 3482 8248
rect 26878 8236 26884 8248
rect 26936 8236 26942 8288
rect 26970 8236 26976 8288
rect 27028 8276 27034 8288
rect 27341 8279 27399 8285
rect 27341 8276 27353 8279
rect 27028 8248 27353 8276
rect 27028 8236 27034 8248
rect 27341 8245 27353 8248
rect 27387 8245 27399 8279
rect 27341 8239 27399 8245
rect 27614 8236 27620 8288
rect 27672 8276 27678 8288
rect 32600 8276 32628 8316
rect 27672 8248 32628 8276
rect 32784 8276 32812 8316
rect 65426 8304 65432 8356
rect 65484 8304 65490 8356
rect 66364 8344 66392 8384
rect 66625 8381 66637 8415
rect 66671 8412 66683 8415
rect 67453 8415 67511 8421
rect 67453 8412 67465 8415
rect 66671 8384 67465 8412
rect 66671 8381 66683 8384
rect 66625 8375 66683 8381
rect 67453 8381 67465 8384
rect 67499 8381 67511 8415
rect 67453 8375 67511 8381
rect 71590 8372 71596 8424
rect 71648 8372 71654 8424
rect 74534 8372 74540 8424
rect 74592 8372 74598 8424
rect 79689 8415 79747 8421
rect 79689 8381 79701 8415
rect 79735 8381 79747 8415
rect 79689 8375 79747 8381
rect 66898 8344 66904 8356
rect 66364 8316 66904 8344
rect 66898 8304 66904 8316
rect 66956 8304 66962 8356
rect 51350 8276 51356 8288
rect 32784 8248 51356 8276
rect 27672 8236 27678 8248
rect 51350 8236 51356 8248
rect 51408 8236 51414 8288
rect 79704 8276 79732 8375
rect 81894 8372 81900 8424
rect 81952 8372 81958 8424
rect 88150 8372 88156 8424
rect 88208 8412 88214 8424
rect 89441 8415 89499 8421
rect 89441 8412 89453 8415
rect 88208 8384 89453 8412
rect 88208 8372 88214 8384
rect 89441 8381 89453 8384
rect 89487 8412 89499 8415
rect 89717 8415 89775 8421
rect 89717 8412 89729 8415
rect 89487 8384 89729 8412
rect 89487 8381 89499 8384
rect 89441 8375 89499 8381
rect 89717 8381 89729 8384
rect 89763 8412 89775 8415
rect 92934 8412 92940 8424
rect 89763 8384 92940 8412
rect 89763 8381 89775 8384
rect 89717 8375 89775 8381
rect 92934 8372 92940 8384
rect 92992 8372 92998 8424
rect 104158 8412 104164 8424
rect 96540 8384 104164 8412
rect 90008 8316 90220 8344
rect 84194 8276 84200 8288
rect 79704 8248 84200 8276
rect 84194 8236 84200 8248
rect 84252 8236 84258 8288
rect 84838 8236 84844 8288
rect 84896 8276 84902 8288
rect 90008 8276 90036 8316
rect 84896 8248 90036 8276
rect 84896 8236 84902 8248
rect 90082 8236 90088 8288
rect 90140 8236 90146 8288
rect 90192 8276 90220 8316
rect 93044 8316 93624 8344
rect 93044 8276 93072 8316
rect 90192 8248 93072 8276
rect 93118 8236 93124 8288
rect 93176 8276 93182 8288
rect 93489 8279 93547 8285
rect 93489 8276 93501 8279
rect 93176 8248 93501 8276
rect 93176 8236 93182 8248
rect 93489 8245 93501 8248
rect 93535 8245 93547 8279
rect 93596 8276 93624 8316
rect 94222 8304 94228 8356
rect 94280 8344 94286 8356
rect 96540 8344 96568 8384
rect 104158 8372 104164 8384
rect 104216 8372 104222 8424
rect 114554 8372 114560 8424
rect 114612 8412 114618 8424
rect 115842 8412 115848 8424
rect 114612 8384 115848 8412
rect 114612 8372 114618 8384
rect 115842 8372 115848 8384
rect 115900 8372 115906 8424
rect 125042 8372 125048 8424
rect 125100 8412 125106 8424
rect 128832 8412 128860 8520
rect 129090 8440 129096 8492
rect 129148 8440 129154 8492
rect 129277 8483 129335 8489
rect 129277 8449 129289 8483
rect 129323 8480 129335 8483
rect 129550 8480 129556 8492
rect 129323 8452 129556 8480
rect 129323 8449 129335 8452
rect 129277 8443 129335 8449
rect 129550 8440 129556 8452
rect 129608 8480 129614 8492
rect 130749 8483 130807 8489
rect 130749 8480 130761 8483
rect 129608 8452 130761 8480
rect 129608 8440 129614 8452
rect 130749 8449 130761 8452
rect 130795 8449 130807 8483
rect 130749 8443 130807 8449
rect 130933 8483 130991 8489
rect 130933 8449 130945 8483
rect 130979 8480 130991 8483
rect 131393 8483 131451 8489
rect 131393 8480 131405 8483
rect 130979 8452 131405 8480
rect 130979 8449 130991 8452
rect 130933 8443 130991 8449
rect 131393 8449 131405 8452
rect 131439 8449 131451 8483
rect 131393 8443 131451 8449
rect 132126 8440 132132 8492
rect 132184 8440 132190 8492
rect 132862 8440 132868 8492
rect 132920 8480 132926 8492
rect 132957 8483 133015 8489
rect 132957 8480 132969 8483
rect 132920 8452 132969 8480
rect 132920 8440 132926 8452
rect 132957 8449 132969 8452
rect 133003 8449 133015 8483
rect 132957 8443 133015 8449
rect 133138 8440 133144 8492
rect 133196 8440 133202 8492
rect 134242 8440 134248 8492
rect 134300 8440 134306 8492
rect 134337 8483 134395 8489
rect 134337 8449 134349 8483
rect 134383 8449 134395 8483
rect 134337 8443 134395 8449
rect 130562 8412 130568 8424
rect 125100 8384 128860 8412
rect 128924 8384 130568 8412
rect 125100 8372 125106 8384
rect 94280 8316 96568 8344
rect 94280 8304 94286 8316
rect 96614 8304 96620 8356
rect 96672 8344 96678 8356
rect 96672 8316 128354 8344
rect 96672 8304 96678 8316
rect 104894 8276 104900 8288
rect 93596 8248 104900 8276
rect 93489 8239 93547 8245
rect 104894 8236 104900 8248
rect 104952 8236 104958 8288
rect 105722 8236 105728 8288
rect 105780 8276 105786 8288
rect 107930 8276 107936 8288
rect 105780 8248 107936 8276
rect 105780 8236 105786 8248
rect 107930 8236 107936 8248
rect 107988 8236 107994 8288
rect 128326 8276 128354 8316
rect 128924 8276 128952 8384
rect 130562 8372 130568 8384
rect 130620 8372 130626 8424
rect 133156 8412 133184 8440
rect 134352 8412 134380 8443
rect 133156 8384 134380 8412
rect 128998 8304 129004 8356
rect 129056 8344 129062 8356
rect 137370 8344 137376 8356
rect 129056 8316 137376 8344
rect 129056 8304 129062 8316
rect 137370 8304 137376 8316
rect 137428 8304 137434 8356
rect 137986 8344 138014 8520
rect 160830 8508 160836 8560
rect 160888 8548 160894 8560
rect 161860 8548 161888 8588
rect 160888 8520 161888 8548
rect 164206 8548 164234 8588
rect 165154 8576 165160 8628
rect 165212 8576 165218 8628
rect 169938 8576 169944 8628
rect 169996 8576 170002 8628
rect 170030 8576 170036 8628
rect 170088 8616 170094 8628
rect 185854 8616 185860 8628
rect 170088 8588 185860 8616
rect 170088 8576 170094 8588
rect 185854 8576 185860 8588
rect 185912 8576 185918 8628
rect 185946 8576 185952 8628
rect 186004 8616 186010 8628
rect 186004 8588 188752 8616
rect 186004 8576 186010 8588
rect 187694 8548 187700 8560
rect 164206 8520 187700 8548
rect 160888 8508 160894 8520
rect 187694 8508 187700 8520
rect 187752 8508 187758 8560
rect 148686 8440 148692 8492
rect 148744 8480 148750 8492
rect 156693 8483 156751 8489
rect 148744 8452 156644 8480
rect 148744 8440 148750 8452
rect 156506 8372 156512 8424
rect 156564 8372 156570 8424
rect 156616 8412 156644 8452
rect 156693 8449 156705 8483
rect 156739 8480 156751 8483
rect 157610 8480 157616 8492
rect 156739 8452 157616 8480
rect 156739 8449 156751 8452
rect 156693 8443 156751 8449
rect 157610 8440 157616 8452
rect 157668 8480 157674 8492
rect 158165 8483 158223 8489
rect 158165 8480 158177 8483
rect 157668 8452 158177 8480
rect 157668 8440 157674 8452
rect 158165 8449 158177 8452
rect 158211 8480 158223 8483
rect 159177 8483 159235 8489
rect 159177 8480 159189 8483
rect 158211 8452 159189 8480
rect 158211 8449 158223 8452
rect 158165 8443 158223 8449
rect 159177 8449 159189 8452
rect 159223 8480 159235 8483
rect 160005 8483 160063 8489
rect 160005 8480 160017 8483
rect 159223 8452 160017 8480
rect 159223 8449 159235 8452
rect 159177 8443 159235 8449
rect 160005 8449 160017 8452
rect 160051 8449 160063 8483
rect 160005 8443 160063 8449
rect 161201 8483 161259 8489
rect 161201 8449 161213 8483
rect 161247 8480 161259 8483
rect 161934 8480 161940 8492
rect 161247 8452 161940 8480
rect 161247 8449 161259 8452
rect 161201 8443 161259 8449
rect 157242 8412 157248 8424
rect 156616 8384 157248 8412
rect 157242 8372 157248 8384
rect 157300 8372 157306 8424
rect 157981 8415 158039 8421
rect 157981 8381 157993 8415
rect 158027 8412 158039 8415
rect 158714 8412 158720 8424
rect 158027 8384 158720 8412
rect 158027 8381 158039 8384
rect 157981 8375 158039 8381
rect 158714 8372 158720 8384
rect 158772 8372 158778 8424
rect 158993 8415 159051 8421
rect 158993 8381 159005 8415
rect 159039 8412 159051 8415
rect 159082 8412 159088 8424
rect 159039 8384 159088 8412
rect 159039 8381 159051 8384
rect 158993 8375 159051 8381
rect 159082 8372 159088 8384
rect 159140 8372 159146 8424
rect 159818 8372 159824 8424
rect 159876 8372 159882 8424
rect 160020 8412 160048 8443
rect 161934 8440 161940 8452
rect 161992 8440 161998 8492
rect 162489 8483 162547 8489
rect 162489 8449 162501 8483
rect 162535 8480 162547 8483
rect 162670 8480 162676 8492
rect 162535 8452 162676 8480
rect 162535 8449 162547 8452
rect 162489 8443 162547 8449
rect 162670 8440 162676 8452
rect 162728 8440 162734 8492
rect 163317 8483 163375 8489
rect 163317 8449 163329 8483
rect 163363 8480 163375 8483
rect 163682 8480 163688 8492
rect 163363 8452 163688 8480
rect 163363 8449 163375 8452
rect 163317 8443 163375 8449
rect 163682 8440 163688 8452
rect 163740 8440 163746 8492
rect 164973 8483 165031 8489
rect 164973 8449 164985 8483
rect 165019 8480 165031 8483
rect 165522 8480 165528 8492
rect 165019 8452 165528 8480
rect 165019 8449 165031 8452
rect 164973 8443 165031 8449
rect 165522 8440 165528 8452
rect 165580 8440 165586 8492
rect 166813 8483 166871 8489
rect 166813 8449 166825 8483
rect 166859 8480 166871 8483
rect 167362 8480 167368 8492
rect 166859 8452 167368 8480
rect 166859 8449 166871 8452
rect 166813 8443 166871 8449
rect 167362 8440 167368 8452
rect 167420 8440 167426 8492
rect 168285 8483 168343 8489
rect 168285 8449 168297 8483
rect 168331 8480 168343 8483
rect 168331 8452 169708 8480
rect 168331 8449 168343 8452
rect 168285 8443 168343 8449
rect 161566 8412 161572 8424
rect 160020 8384 161572 8412
rect 161566 8372 161572 8384
rect 161624 8372 161630 8424
rect 161661 8415 161719 8421
rect 161661 8381 161673 8415
rect 161707 8381 161719 8415
rect 161661 8375 161719 8381
rect 159100 8344 159128 8372
rect 159910 8344 159916 8356
rect 137986 8316 159916 8344
rect 159910 8304 159916 8316
rect 159968 8304 159974 8356
rect 160922 8304 160928 8356
rect 160980 8344 160986 8356
rect 161676 8344 161704 8375
rect 161750 8372 161756 8424
rect 161808 8412 161814 8424
rect 162210 8412 162216 8424
rect 161808 8384 162216 8412
rect 161808 8372 161814 8384
rect 162210 8372 162216 8384
rect 162268 8412 162274 8424
rect 162305 8415 162363 8421
rect 162305 8412 162317 8415
rect 162268 8384 162317 8412
rect 162268 8372 162274 8384
rect 162305 8381 162317 8384
rect 162351 8412 162363 8415
rect 162762 8412 162768 8424
rect 162351 8384 162768 8412
rect 162351 8381 162363 8384
rect 162305 8375 162363 8381
rect 162762 8372 162768 8384
rect 162820 8372 162826 8424
rect 163958 8372 163964 8424
rect 164016 8412 164022 8424
rect 164142 8412 164148 8424
rect 164016 8384 164148 8412
rect 164016 8372 164022 8384
rect 164142 8372 164148 8384
rect 164200 8412 164206 8424
rect 164789 8415 164847 8421
rect 164789 8412 164801 8415
rect 164200 8384 164801 8412
rect 164200 8372 164206 8384
rect 164789 8381 164801 8384
rect 164835 8381 164847 8415
rect 164789 8375 164847 8381
rect 167086 8372 167092 8424
rect 167144 8372 167150 8424
rect 167730 8372 167736 8424
rect 167788 8412 167794 8424
rect 168098 8412 168104 8424
rect 167788 8384 168104 8412
rect 167788 8372 167794 8384
rect 168098 8372 168104 8384
rect 168156 8412 168162 8424
rect 168469 8415 168527 8421
rect 168469 8412 168481 8415
rect 168156 8384 168481 8412
rect 168156 8372 168162 8384
rect 168469 8381 168481 8384
rect 168515 8381 168527 8415
rect 168469 8375 168527 8381
rect 169570 8372 169576 8424
rect 169628 8372 169634 8424
rect 169680 8412 169708 8452
rect 169754 8440 169760 8492
rect 169812 8440 169818 8492
rect 173434 8440 173440 8492
rect 173492 8480 173498 8492
rect 173492 8452 180104 8480
rect 173492 8440 173498 8452
rect 179966 8412 179972 8424
rect 169680 8384 179972 8412
rect 179966 8372 179972 8384
rect 180024 8372 180030 8424
rect 180076 8412 180104 8452
rect 183278 8440 183284 8492
rect 183336 8440 183342 8492
rect 186958 8440 186964 8492
rect 187016 8440 187022 8492
rect 187050 8440 187056 8492
rect 187108 8480 187114 8492
rect 187237 8483 187295 8489
rect 187237 8480 187249 8483
rect 187108 8452 187249 8480
rect 187108 8440 187114 8452
rect 187237 8449 187249 8452
rect 187283 8449 187295 8483
rect 187237 8443 187295 8449
rect 188430 8440 188436 8492
rect 188488 8440 188494 8492
rect 188724 8489 188752 8588
rect 189902 8576 189908 8628
rect 189960 8616 189966 8628
rect 190549 8619 190607 8625
rect 190549 8616 190561 8619
rect 189960 8588 190561 8616
rect 189960 8576 189966 8588
rect 190549 8585 190561 8588
rect 190595 8585 190607 8619
rect 190549 8579 190607 8585
rect 191282 8576 191288 8628
rect 191340 8576 191346 8628
rect 191374 8576 191380 8628
rect 191432 8616 191438 8628
rect 192205 8619 192263 8625
rect 192205 8616 192217 8619
rect 191432 8588 192217 8616
rect 191432 8576 191438 8588
rect 192205 8585 192217 8588
rect 192251 8585 192263 8619
rect 192205 8579 192263 8585
rect 193582 8576 193588 8628
rect 193640 8576 193646 8628
rect 194226 8576 194232 8628
rect 194284 8576 194290 8628
rect 195606 8576 195612 8628
rect 195664 8576 195670 8628
rect 196618 8576 196624 8628
rect 196676 8576 196682 8628
rect 197538 8576 197544 8628
rect 197596 8576 197602 8628
rect 197909 8619 197967 8625
rect 197909 8585 197921 8619
rect 197955 8616 197967 8619
rect 198090 8616 198096 8628
rect 197955 8588 198096 8616
rect 197955 8585 197967 8588
rect 197909 8579 197967 8585
rect 198090 8576 198096 8588
rect 198148 8576 198154 8628
rect 198826 8576 198832 8628
rect 198884 8576 198890 8628
rect 199470 8576 199476 8628
rect 199528 8576 199534 8628
rect 200850 8576 200856 8628
rect 200908 8576 200914 8628
rect 200942 8576 200948 8628
rect 201000 8616 201006 8628
rect 201589 8619 201647 8625
rect 201589 8616 201601 8619
rect 201000 8588 201601 8616
rect 201000 8576 201006 8588
rect 201589 8585 201601 8588
rect 201635 8585 201647 8619
rect 201589 8579 201647 8585
rect 202690 8576 202696 8628
rect 202748 8576 202754 8628
rect 203518 8576 203524 8628
rect 203576 8576 203582 8628
rect 225874 8616 225880 8628
rect 203628 8588 225880 8616
rect 196526 8508 196532 8560
rect 196584 8548 196590 8560
rect 196584 8520 203380 8548
rect 196584 8508 196590 8520
rect 188709 8483 188767 8489
rect 188709 8449 188721 8483
rect 188755 8449 188767 8483
rect 188709 8443 188767 8449
rect 190362 8440 190368 8492
rect 190420 8440 190426 8492
rect 191101 8483 191159 8489
rect 191101 8449 191113 8483
rect 191147 8480 191159 8483
rect 191926 8480 191932 8492
rect 191147 8452 191932 8480
rect 191147 8449 191159 8452
rect 191101 8443 191159 8449
rect 191926 8440 191932 8452
rect 191984 8440 191990 8492
rect 192018 8440 192024 8492
rect 192076 8440 192082 8492
rect 193214 8440 193220 8492
rect 193272 8440 193278 8492
rect 193401 8483 193459 8489
rect 193401 8449 193413 8483
rect 193447 8480 193459 8483
rect 193490 8480 193496 8492
rect 193447 8452 193496 8480
rect 193447 8449 193459 8452
rect 193401 8443 193459 8449
rect 193490 8440 193496 8452
rect 193548 8440 193554 8492
rect 194042 8440 194048 8492
rect 194100 8440 194106 8492
rect 195425 8483 195483 8489
rect 195425 8449 195437 8483
rect 195471 8480 195483 8483
rect 196342 8480 196348 8492
rect 195471 8452 196348 8480
rect 195471 8449 195483 8452
rect 195425 8443 195483 8449
rect 196342 8440 196348 8452
rect 196400 8440 196406 8492
rect 196437 8483 196495 8489
rect 196437 8449 196449 8483
rect 196483 8480 196495 8483
rect 196544 8480 196572 8508
rect 196483 8452 196572 8480
rect 196483 8449 196495 8452
rect 196437 8443 196495 8449
rect 197354 8440 197360 8492
rect 197412 8480 197418 8492
rect 198645 8483 198703 8489
rect 198645 8480 198657 8483
rect 197412 8452 198657 8480
rect 197412 8440 197418 8452
rect 198645 8449 198657 8452
rect 198691 8449 198703 8483
rect 198645 8443 198703 8449
rect 199286 8440 199292 8492
rect 199344 8440 199350 8492
rect 200669 8483 200727 8489
rect 200669 8449 200681 8483
rect 200715 8480 200727 8483
rect 201034 8480 201040 8492
rect 200715 8452 201040 8480
rect 200715 8449 200727 8452
rect 200669 8443 200727 8449
rect 201034 8440 201040 8452
rect 201092 8440 201098 8492
rect 201405 8483 201463 8489
rect 201405 8449 201417 8483
rect 201451 8480 201463 8483
rect 202414 8480 202420 8492
rect 201451 8452 202420 8480
rect 201451 8449 201463 8452
rect 201405 8443 201463 8449
rect 202414 8440 202420 8452
rect 202472 8440 202478 8492
rect 202506 8440 202512 8492
rect 202564 8440 202570 8492
rect 203352 8489 203380 8520
rect 203337 8483 203395 8489
rect 203337 8449 203349 8483
rect 203383 8449 203395 8483
rect 203337 8443 203395 8449
rect 183557 8415 183615 8421
rect 183557 8412 183569 8415
rect 180076 8384 183569 8412
rect 183557 8381 183569 8384
rect 183603 8381 183615 8415
rect 183557 8375 183615 8381
rect 196253 8415 196311 8421
rect 196253 8381 196265 8415
rect 196299 8412 196311 8415
rect 196526 8412 196532 8424
rect 196299 8384 196532 8412
rect 196299 8381 196311 8384
rect 196253 8375 196311 8381
rect 196526 8372 196532 8384
rect 196584 8412 196590 8424
rect 196710 8412 196716 8424
rect 196584 8384 196716 8412
rect 196584 8372 196590 8384
rect 196710 8372 196716 8384
rect 196768 8372 196774 8424
rect 197173 8415 197231 8421
rect 197173 8381 197185 8415
rect 197219 8412 197231 8415
rect 197262 8412 197268 8424
rect 197219 8384 197268 8412
rect 197219 8381 197231 8384
rect 197173 8375 197231 8381
rect 197262 8372 197268 8384
rect 197320 8412 197326 8424
rect 198090 8412 198096 8424
rect 197320 8384 198096 8412
rect 197320 8372 197326 8384
rect 198090 8372 198096 8384
rect 198148 8372 198154 8424
rect 198461 8415 198519 8421
rect 198461 8381 198473 8415
rect 198507 8412 198519 8415
rect 198826 8412 198832 8424
rect 198507 8384 198832 8412
rect 198507 8381 198519 8384
rect 198461 8375 198519 8381
rect 198826 8372 198832 8384
rect 198884 8372 198890 8424
rect 202230 8372 202236 8424
rect 202288 8412 202294 8424
rect 202325 8415 202383 8421
rect 202325 8412 202337 8415
rect 202288 8384 202337 8412
rect 202288 8372 202294 8384
rect 202325 8381 202337 8384
rect 202371 8412 202383 8415
rect 202782 8412 202788 8424
rect 202371 8384 202788 8412
rect 202371 8381 202383 8384
rect 202325 8375 202383 8381
rect 202782 8372 202788 8384
rect 202840 8412 202846 8424
rect 202969 8415 203027 8421
rect 202969 8412 202981 8415
rect 202840 8384 202981 8412
rect 202840 8372 202846 8384
rect 202969 8381 202981 8384
rect 203015 8381 203027 8415
rect 202969 8375 203027 8381
rect 203150 8372 203156 8424
rect 203208 8372 203214 8424
rect 160980 8316 161704 8344
rect 160980 8304 160986 8316
rect 161934 8304 161940 8356
rect 161992 8344 161998 8356
rect 162121 8347 162179 8353
rect 162121 8344 162133 8347
rect 161992 8316 162133 8344
rect 161992 8304 161998 8316
rect 162121 8313 162133 8316
rect 162167 8344 162179 8347
rect 162167 8316 162808 8344
rect 162167 8313 162179 8316
rect 162121 8307 162179 8313
rect 128326 8248 128952 8276
rect 132862 8236 132868 8288
rect 132920 8276 132926 8288
rect 133325 8279 133383 8285
rect 133325 8276 133337 8279
rect 132920 8248 133337 8276
rect 132920 8236 132926 8248
rect 133325 8245 133337 8248
rect 133371 8245 133383 8279
rect 133325 8239 133383 8245
rect 146846 8236 146852 8288
rect 146904 8276 146910 8288
rect 151722 8276 151728 8288
rect 146904 8248 151728 8276
rect 146904 8236 146910 8248
rect 151722 8236 151728 8248
rect 151780 8236 151786 8288
rect 160094 8236 160100 8288
rect 160152 8276 160158 8288
rect 160189 8279 160247 8285
rect 160189 8276 160201 8279
rect 160152 8248 160201 8276
rect 160152 8236 160158 8248
rect 160189 8245 160201 8248
rect 160235 8245 160247 8279
rect 160189 8239 160247 8245
rect 162394 8236 162400 8288
rect 162452 8276 162458 8288
rect 162673 8279 162731 8285
rect 162673 8276 162685 8279
rect 162452 8248 162685 8276
rect 162452 8236 162458 8248
rect 162673 8245 162685 8248
rect 162719 8245 162731 8279
rect 162780 8276 162808 8316
rect 162854 8304 162860 8356
rect 162912 8344 162918 8356
rect 170030 8344 170036 8356
rect 162912 8316 170036 8344
rect 162912 8304 162918 8316
rect 170030 8304 170036 8316
rect 170088 8304 170094 8356
rect 196342 8304 196348 8356
rect 196400 8344 196406 8356
rect 196400 8316 201080 8344
rect 196400 8304 196406 8316
rect 163314 8276 163320 8288
rect 162780 8248 163320 8276
rect 162673 8239 162731 8245
rect 163314 8236 163320 8248
rect 163372 8236 163378 8288
rect 201052 8276 201080 8316
rect 201126 8304 201132 8356
rect 201184 8344 201190 8356
rect 203628 8344 203656 8588
rect 225874 8576 225880 8588
rect 225932 8576 225938 8628
rect 225966 8576 225972 8628
rect 226024 8576 226030 8628
rect 226702 8576 226708 8628
rect 226760 8576 226766 8628
rect 228266 8576 228272 8628
rect 228324 8576 228330 8628
rect 229094 8576 229100 8628
rect 229152 8576 229158 8628
rect 231026 8576 231032 8628
rect 231084 8576 231090 8628
rect 231946 8576 231952 8628
rect 232004 8576 232010 8628
rect 232866 8576 232872 8628
rect 232924 8616 232930 8628
rect 233421 8619 233479 8625
rect 233421 8616 233433 8619
rect 232924 8588 233433 8616
rect 232924 8576 232930 8588
rect 233421 8585 233433 8588
rect 233467 8585 233479 8619
rect 233421 8579 233479 8585
rect 234890 8576 234896 8628
rect 234948 8576 234954 8628
rect 235997 8619 236055 8625
rect 235997 8585 236009 8619
rect 236043 8616 236055 8619
rect 236086 8616 236092 8628
rect 236043 8588 236092 8616
rect 236043 8585 236055 8588
rect 235997 8579 236055 8585
rect 236086 8576 236092 8588
rect 236144 8576 236150 8628
rect 236638 8576 236644 8628
rect 236696 8576 236702 8628
rect 242986 8576 242992 8628
rect 243044 8616 243050 8628
rect 247770 8616 247776 8628
rect 243044 8588 247776 8616
rect 243044 8576 243050 8588
rect 247770 8576 247776 8588
rect 247828 8576 247834 8628
rect 258258 8576 258264 8628
rect 258316 8576 258322 8628
rect 262582 8616 262588 8628
rect 260116 8588 262588 8616
rect 223942 8548 223948 8560
rect 209746 8520 223948 8548
rect 209746 8480 209774 8520
rect 223942 8508 223948 8520
rect 224000 8508 224006 8560
rect 224770 8548 224776 8560
rect 224420 8520 224776 8548
rect 201184 8316 203656 8344
rect 203720 8452 209774 8480
rect 201184 8304 201190 8316
rect 203720 8276 203748 8452
rect 217962 8440 217968 8492
rect 218020 8480 218026 8492
rect 220906 8480 220912 8492
rect 218020 8452 220912 8480
rect 218020 8440 218026 8452
rect 220906 8440 220912 8452
rect 220964 8440 220970 8492
rect 221826 8440 221832 8492
rect 221884 8480 221890 8492
rect 223666 8480 223672 8492
rect 221884 8452 223672 8480
rect 221884 8440 221890 8452
rect 223666 8440 223672 8452
rect 223724 8440 223730 8492
rect 224420 8489 224448 8520
rect 224770 8508 224776 8520
rect 224828 8508 224834 8560
rect 224862 8508 224868 8560
rect 224920 8548 224926 8560
rect 224920 8520 229784 8548
rect 224920 8508 224926 8520
rect 224405 8483 224463 8489
rect 224405 8449 224417 8483
rect 224451 8449 224463 8483
rect 224405 8443 224463 8449
rect 224589 8483 224647 8489
rect 224589 8449 224601 8483
rect 224635 8480 224647 8483
rect 225049 8483 225107 8489
rect 225049 8480 225061 8483
rect 224635 8452 225061 8480
rect 224635 8449 224647 8452
rect 224589 8443 224647 8449
rect 225049 8449 225061 8452
rect 225095 8449 225107 8483
rect 225049 8443 225107 8449
rect 225782 8440 225788 8492
rect 225840 8440 225846 8492
rect 226518 8440 226524 8492
rect 226576 8440 226582 8492
rect 228082 8440 228088 8492
rect 228140 8440 228146 8492
rect 228910 8440 228916 8492
rect 228968 8440 228974 8492
rect 229462 8440 229468 8492
rect 229520 8480 229526 8492
rect 229756 8480 229784 8520
rect 229830 8508 229836 8560
rect 229888 8548 229894 8560
rect 229888 8520 230060 8548
rect 229888 8508 229894 8520
rect 229922 8480 229928 8492
rect 229520 8452 229692 8480
rect 229756 8452 229928 8480
rect 229520 8440 229526 8452
rect 212350 8372 212356 8424
rect 212408 8412 212414 8424
rect 212408 8384 218008 8412
rect 212408 8372 212414 8384
rect 201052 8248 203748 8276
rect 211062 8236 211068 8288
rect 211120 8276 211126 8288
rect 214558 8276 214564 8288
rect 211120 8248 214564 8276
rect 211120 8236 211126 8248
rect 214558 8236 214564 8248
rect 214616 8236 214622 8288
rect 217980 8276 218008 8384
rect 223482 8372 223488 8424
rect 223540 8412 223546 8424
rect 223853 8415 223911 8421
rect 223853 8412 223865 8415
rect 223540 8384 223865 8412
rect 223540 8372 223546 8384
rect 223853 8381 223865 8384
rect 223899 8412 223911 8415
rect 224221 8415 224279 8421
rect 224221 8412 224233 8415
rect 223899 8384 224233 8412
rect 223899 8381 223911 8384
rect 223853 8375 223911 8381
rect 224221 8381 224233 8384
rect 224267 8381 224279 8415
rect 229554 8412 229560 8424
rect 224221 8375 224279 8381
rect 224328 8384 229560 8412
rect 224328 8344 224356 8384
rect 229554 8372 229560 8384
rect 229612 8372 229618 8424
rect 229664 8412 229692 8452
rect 229922 8440 229928 8452
rect 229980 8440 229986 8492
rect 230032 8489 230060 8520
rect 230106 8508 230112 8560
rect 230164 8548 230170 8560
rect 260116 8548 260144 8588
rect 262582 8576 262588 8588
rect 262640 8576 262646 8628
rect 263229 8619 263287 8625
rect 263229 8585 263241 8619
rect 263275 8616 263287 8619
rect 263594 8616 263600 8628
rect 263275 8588 263600 8616
rect 263275 8585 263287 8588
rect 263229 8579 263287 8585
rect 263594 8576 263600 8588
rect 263652 8616 263658 8628
rect 264238 8616 264244 8628
rect 263652 8588 264244 8616
rect 263652 8576 263658 8588
rect 264238 8576 264244 8588
rect 264296 8576 264302 8628
rect 264882 8576 264888 8628
rect 264940 8616 264946 8628
rect 267458 8616 267464 8628
rect 264940 8588 267464 8616
rect 264940 8576 264946 8588
rect 267458 8576 267464 8588
rect 267516 8576 267522 8628
rect 267642 8576 267648 8628
rect 267700 8616 267706 8628
rect 268286 8616 268292 8628
rect 267700 8588 268292 8616
rect 267700 8576 267706 8588
rect 268286 8576 268292 8588
rect 268344 8576 268350 8628
rect 268381 8619 268439 8625
rect 268381 8585 268393 8619
rect 268427 8616 268439 8619
rect 270218 8616 270224 8628
rect 268427 8588 270224 8616
rect 268427 8585 268439 8588
rect 268381 8579 268439 8585
rect 270218 8576 270224 8588
rect 270276 8576 270282 8628
rect 230164 8520 260144 8548
rect 230164 8508 230170 8520
rect 260926 8508 260932 8560
rect 260984 8548 260990 8560
rect 266081 8551 266139 8557
rect 266081 8548 266093 8551
rect 260984 8520 266093 8548
rect 260984 8508 260990 8520
rect 266081 8517 266093 8520
rect 266127 8548 266139 8551
rect 266725 8551 266783 8557
rect 266725 8548 266737 8551
rect 266127 8520 266737 8548
rect 266127 8517 266139 8520
rect 266081 8511 266139 8517
rect 266725 8517 266737 8520
rect 266771 8548 266783 8551
rect 266906 8548 266912 8560
rect 266771 8520 266912 8548
rect 266771 8517 266783 8520
rect 266725 8511 266783 8517
rect 266906 8508 266912 8520
rect 266964 8508 266970 8560
rect 230017 8483 230075 8489
rect 230017 8449 230029 8483
rect 230063 8449 230075 8483
rect 230017 8443 230075 8449
rect 230658 8440 230664 8492
rect 230716 8440 230722 8492
rect 230842 8440 230848 8492
rect 230900 8440 230906 8492
rect 231762 8440 231768 8492
rect 231820 8440 231826 8492
rect 233234 8440 233240 8492
rect 233292 8440 233298 8492
rect 234522 8440 234528 8492
rect 234580 8440 234586 8492
rect 234709 8483 234767 8489
rect 234709 8449 234721 8483
rect 234755 8449 234767 8483
rect 234709 8443 234767 8449
rect 229830 8412 229836 8424
rect 229664 8384 229836 8412
rect 229830 8372 229836 8384
rect 229888 8372 229894 8424
rect 230676 8412 230704 8440
rect 231026 8412 231032 8424
rect 230676 8384 231032 8412
rect 231026 8372 231032 8384
rect 231084 8372 231090 8424
rect 234724 8412 234752 8443
rect 235718 8440 235724 8492
rect 235776 8440 235782 8492
rect 235813 8483 235871 8489
rect 235813 8449 235825 8483
rect 235859 8480 235871 8483
rect 235902 8480 235908 8492
rect 235859 8452 235908 8480
rect 235859 8449 235871 8452
rect 235813 8443 235871 8449
rect 235828 8412 235856 8443
rect 235902 8440 235908 8452
rect 235960 8440 235966 8492
rect 236178 8440 236184 8492
rect 236236 8480 236242 8492
rect 236457 8483 236515 8489
rect 236457 8480 236469 8483
rect 236236 8452 236469 8480
rect 236236 8440 236242 8452
rect 236457 8449 236469 8452
rect 236503 8449 236515 8483
rect 236457 8443 236515 8449
rect 246390 8440 246396 8492
rect 246448 8440 246454 8492
rect 246666 8440 246672 8492
rect 246724 8440 246730 8492
rect 249334 8440 249340 8492
rect 249392 8440 249398 8492
rect 251542 8440 251548 8492
rect 251600 8440 251606 8492
rect 254486 8440 254492 8492
rect 254544 8440 254550 8492
rect 256694 8440 256700 8492
rect 256752 8440 256758 8492
rect 258074 8440 258080 8492
rect 258132 8440 258138 8492
rect 258350 8440 258356 8492
rect 258408 8480 258414 8492
rect 259178 8480 259184 8492
rect 258408 8452 259184 8480
rect 258408 8440 258414 8452
rect 259178 8440 259184 8452
rect 259236 8480 259242 8492
rect 260193 8483 260251 8489
rect 260193 8480 260205 8483
rect 259236 8452 260205 8480
rect 259236 8440 259242 8452
rect 260193 8449 260205 8452
rect 260239 8480 260251 8483
rect 260239 8452 260604 8480
rect 260239 8449 260251 8452
rect 260193 8443 260251 8449
rect 234724 8384 235856 8412
rect 236362 8372 236368 8424
rect 236420 8412 236426 8424
rect 242894 8412 242900 8424
rect 236420 8384 242900 8412
rect 236420 8372 236426 8384
rect 242894 8372 242900 8384
rect 242952 8372 242958 8424
rect 249610 8372 249616 8424
rect 249668 8372 249674 8424
rect 251818 8372 251824 8424
rect 251876 8372 251882 8424
rect 254762 8372 254768 8424
rect 254820 8372 254826 8424
rect 256973 8415 257031 8421
rect 256973 8381 256985 8415
rect 257019 8381 257031 8415
rect 256973 8375 257031 8381
rect 223500 8316 224356 8344
rect 223500 8276 223528 8316
rect 224770 8304 224776 8356
rect 224828 8344 224834 8356
rect 225233 8347 225291 8353
rect 225233 8344 225245 8347
rect 224828 8316 225245 8344
rect 224828 8304 224834 8316
rect 225233 8313 225245 8316
rect 225279 8313 225291 8347
rect 225233 8307 225291 8313
rect 226426 8304 226432 8356
rect 226484 8344 226490 8356
rect 227070 8344 227076 8356
rect 226484 8316 227076 8344
rect 226484 8304 226490 8316
rect 227070 8304 227076 8316
rect 227128 8304 227134 8356
rect 230201 8347 230259 8353
rect 230201 8313 230213 8347
rect 230247 8344 230259 8347
rect 230566 8344 230572 8356
rect 230247 8316 230572 8344
rect 230247 8313 230259 8316
rect 230201 8307 230259 8313
rect 230566 8304 230572 8316
rect 230624 8304 230630 8356
rect 234522 8304 234528 8356
rect 234580 8344 234586 8356
rect 234890 8344 234896 8356
rect 234580 8316 234896 8344
rect 234580 8304 234586 8316
rect 234890 8304 234896 8316
rect 234948 8344 234954 8356
rect 237926 8344 237932 8356
rect 234948 8316 237932 8344
rect 234948 8304 234954 8316
rect 237926 8304 237932 8316
rect 237984 8304 237990 8356
rect 238570 8304 238576 8356
rect 238628 8344 238634 8356
rect 256988 8344 257016 8375
rect 258902 8372 258908 8424
rect 258960 8412 258966 8424
rect 258997 8415 259055 8421
rect 258997 8412 259009 8415
rect 258960 8384 259009 8412
rect 258960 8372 258966 8384
rect 258997 8381 259009 8384
rect 259043 8381 259055 8415
rect 258997 8375 259055 8381
rect 259638 8372 259644 8424
rect 259696 8412 259702 8424
rect 260009 8415 260067 8421
rect 260009 8412 260021 8415
rect 259696 8384 260021 8412
rect 259696 8372 259702 8384
rect 260009 8381 260021 8384
rect 260055 8412 260067 8415
rect 260055 8384 260236 8412
rect 260055 8381 260067 8384
rect 260009 8375 260067 8381
rect 260208 8356 260236 8384
rect 238628 8316 257016 8344
rect 238628 8304 238634 8316
rect 260190 8304 260196 8356
rect 260248 8304 260254 8356
rect 260576 8344 260604 8452
rect 261110 8440 261116 8492
rect 261168 8480 261174 8492
rect 261297 8483 261355 8489
rect 261297 8480 261309 8483
rect 261168 8452 261309 8480
rect 261168 8440 261174 8452
rect 261297 8449 261309 8452
rect 261343 8449 261355 8483
rect 261297 8443 261355 8449
rect 261478 8440 261484 8492
rect 261536 8480 261542 8492
rect 261665 8483 261723 8489
rect 261665 8480 261677 8483
rect 261536 8452 261677 8480
rect 261536 8440 261542 8452
rect 261665 8449 261677 8452
rect 261711 8449 261723 8483
rect 261665 8443 261723 8449
rect 262493 8483 262551 8489
rect 262493 8449 262505 8483
rect 262539 8480 262551 8483
rect 263594 8480 263600 8492
rect 262539 8452 263600 8480
rect 262539 8449 262551 8452
rect 262493 8443 262551 8449
rect 263594 8440 263600 8452
rect 263652 8440 263658 8492
rect 264238 8440 264244 8492
rect 264296 8480 264302 8492
rect 264514 8480 264520 8492
rect 264296 8452 264520 8480
rect 264296 8440 264302 8452
rect 264514 8440 264520 8452
rect 264572 8440 264578 8492
rect 265158 8440 265164 8492
rect 265216 8440 265222 8492
rect 265529 8483 265587 8489
rect 265529 8449 265541 8483
rect 265575 8480 265587 8483
rect 265894 8480 265900 8492
rect 265575 8452 265900 8480
rect 265575 8449 265587 8452
rect 265529 8443 265587 8449
rect 265894 8440 265900 8452
rect 265952 8440 265958 8492
rect 266446 8440 266452 8492
rect 266504 8440 266510 8492
rect 267090 8440 267096 8492
rect 267148 8480 267154 8492
rect 267369 8483 267427 8489
rect 267369 8480 267381 8483
rect 267148 8452 267381 8480
rect 267148 8440 267154 8452
rect 267369 8449 267381 8452
rect 267415 8449 267427 8483
rect 267369 8443 267427 8449
rect 267461 8483 267519 8489
rect 267461 8449 267473 8483
rect 267507 8480 267519 8483
rect 267642 8480 267648 8492
rect 267507 8452 267648 8480
rect 267507 8449 267519 8452
rect 267461 8443 267519 8449
rect 260834 8372 260840 8424
rect 260892 8412 260898 8424
rect 263505 8415 263563 8421
rect 263505 8412 263517 8415
rect 260892 8384 263517 8412
rect 260892 8372 260898 8384
rect 263505 8381 263517 8384
rect 263551 8412 263563 8415
rect 265176 8412 265204 8440
rect 263551 8384 265204 8412
rect 263551 8381 263563 8384
rect 263505 8375 263563 8381
rect 265802 8372 265808 8424
rect 265860 8412 265866 8424
rect 266464 8412 266492 8440
rect 265860 8384 266492 8412
rect 267384 8412 267412 8443
rect 267642 8440 267648 8452
rect 267700 8440 267706 8492
rect 267734 8440 267740 8492
rect 267792 8440 267798 8492
rect 268010 8440 268016 8492
rect 268068 8480 268074 8492
rect 268304 8489 268332 8576
rect 268197 8483 268255 8489
rect 268197 8480 268209 8483
rect 268068 8452 268209 8480
rect 268068 8440 268074 8452
rect 268197 8449 268209 8452
rect 268243 8449 268255 8483
rect 268197 8443 268255 8449
rect 268289 8483 268347 8489
rect 268289 8449 268301 8483
rect 268335 8449 268347 8483
rect 268289 8443 268347 8449
rect 268378 8440 268384 8492
rect 268436 8480 268442 8492
rect 268473 8483 268531 8489
rect 268473 8480 268485 8483
rect 268436 8452 268485 8480
rect 268436 8440 268442 8452
rect 268473 8449 268485 8452
rect 268519 8449 268531 8483
rect 268473 8443 268531 8449
rect 268562 8440 268568 8492
rect 268620 8440 268626 8492
rect 268657 8483 268715 8489
rect 268657 8449 268669 8483
rect 268703 8480 268715 8483
rect 268746 8480 268752 8492
rect 268703 8452 268752 8480
rect 268703 8449 268715 8452
rect 268657 8443 268715 8449
rect 268746 8440 268752 8452
rect 268804 8480 268810 8492
rect 268804 8452 269436 8480
rect 268804 8440 268810 8452
rect 268102 8412 268108 8424
rect 267384 8384 268108 8412
rect 265860 8372 265866 8384
rect 268102 8372 268108 8384
rect 268160 8372 268166 8424
rect 269298 8372 269304 8424
rect 269356 8372 269362 8424
rect 269408 8412 269436 8452
rect 269482 8440 269488 8492
rect 269540 8440 269546 8492
rect 270862 8480 270868 8492
rect 269592 8452 270868 8480
rect 269592 8412 269620 8452
rect 270862 8440 270868 8452
rect 270920 8440 270926 8492
rect 269408 8384 269620 8412
rect 269666 8372 269672 8424
rect 269724 8372 269730 8424
rect 270126 8372 270132 8424
rect 270184 8372 270190 8424
rect 270405 8415 270463 8421
rect 270405 8381 270417 8415
rect 270451 8381 270463 8415
rect 270405 8375 270463 8381
rect 261202 8344 261208 8356
rect 260576 8316 261208 8344
rect 261202 8304 261208 8316
rect 261260 8344 261266 8356
rect 261938 8344 261944 8356
rect 261260 8316 261944 8344
rect 261260 8304 261266 8316
rect 261938 8304 261944 8316
rect 261996 8304 262002 8356
rect 263962 8304 263968 8356
rect 264020 8344 264026 8356
rect 264425 8347 264483 8353
rect 264425 8344 264437 8347
rect 264020 8316 264437 8344
rect 264020 8304 264026 8316
rect 264425 8313 264437 8316
rect 264471 8313 264483 8347
rect 264425 8307 264483 8313
rect 268930 8304 268936 8356
rect 268988 8344 268994 8356
rect 270420 8344 270448 8375
rect 268988 8316 270448 8344
rect 268988 8304 268994 8316
rect 217980 8248 223528 8276
rect 223574 8236 223580 8288
rect 223632 8276 223638 8288
rect 228910 8276 228916 8288
rect 223632 8248 228916 8276
rect 223632 8236 223638 8248
rect 228910 8236 228916 8248
rect 228968 8236 228974 8288
rect 235810 8236 235816 8288
rect 235868 8276 235874 8288
rect 236546 8276 236552 8288
rect 235868 8248 236552 8276
rect 235868 8236 235874 8248
rect 236546 8236 236552 8248
rect 236604 8236 236610 8288
rect 236914 8236 236920 8288
rect 236972 8276 236978 8288
rect 243170 8276 243176 8288
rect 236972 8248 243176 8276
rect 236972 8236 236978 8248
rect 243170 8236 243176 8248
rect 243228 8236 243234 8288
rect 258810 8236 258816 8288
rect 258868 8276 258874 8288
rect 259365 8279 259423 8285
rect 259365 8276 259377 8279
rect 258868 8248 259377 8276
rect 258868 8236 258874 8248
rect 259365 8245 259377 8248
rect 259411 8245 259423 8279
rect 259365 8239 259423 8245
rect 260282 8236 260288 8288
rect 260340 8276 260346 8288
rect 260377 8279 260435 8285
rect 260377 8276 260389 8279
rect 260340 8248 260389 8276
rect 260340 8236 260346 8248
rect 260377 8245 260389 8248
rect 260423 8245 260435 8279
rect 260377 8239 260435 8245
rect 262674 8236 262680 8288
rect 262732 8276 262738 8288
rect 264238 8276 264244 8288
rect 262732 8248 264244 8276
rect 262732 8236 262738 8248
rect 264238 8236 264244 8248
rect 264296 8236 264302 8288
rect 267185 8279 267243 8285
rect 267185 8245 267197 8279
rect 267231 8276 267243 8279
rect 267458 8276 267464 8288
rect 267231 8248 267464 8276
rect 267231 8245 267243 8248
rect 267185 8239 267243 8245
rect 267458 8236 267464 8248
rect 267516 8236 267522 8288
rect 267645 8279 267703 8285
rect 267645 8245 267657 8279
rect 267691 8276 267703 8279
rect 268746 8276 268752 8288
rect 267691 8248 268752 8276
rect 267691 8245 267703 8248
rect 267645 8239 267703 8245
rect 268746 8236 268752 8248
rect 268804 8236 268810 8288
rect 1104 8186 271492 8208
rect 1104 8134 34748 8186
rect 34800 8134 34812 8186
rect 34864 8134 34876 8186
rect 34928 8134 34940 8186
rect 34992 8134 35004 8186
rect 35056 8134 102345 8186
rect 102397 8134 102409 8186
rect 102461 8134 102473 8186
rect 102525 8134 102537 8186
rect 102589 8134 102601 8186
rect 102653 8134 169942 8186
rect 169994 8134 170006 8186
rect 170058 8134 170070 8186
rect 170122 8134 170134 8186
rect 170186 8134 170198 8186
rect 170250 8134 237539 8186
rect 237591 8134 237603 8186
rect 237655 8134 237667 8186
rect 237719 8134 237731 8186
rect 237783 8134 237795 8186
rect 237847 8134 271492 8186
rect 1104 8112 271492 8134
rect 25222 8032 25228 8084
rect 25280 8032 25286 8084
rect 28350 8032 28356 8084
rect 28408 8032 28414 8084
rect 47302 8072 47308 8084
rect 28460 8044 47308 8072
rect 23198 7964 23204 8016
rect 23256 8004 23262 8016
rect 28460 8004 28488 8044
rect 47302 8032 47308 8044
rect 47360 8032 47366 8084
rect 118234 8072 118240 8084
rect 89686 8044 118240 8072
rect 23256 7976 28488 8004
rect 23256 7964 23262 7976
rect 28534 7964 28540 8016
rect 28592 8004 28598 8016
rect 48222 8004 48228 8016
rect 28592 7976 48228 8004
rect 28592 7964 28598 7976
rect 48222 7964 48228 7976
rect 48280 7964 48286 8016
rect 73706 7964 73712 8016
rect 73764 8004 73770 8016
rect 82170 8004 82176 8016
rect 73764 7976 82176 8004
rect 73764 7964 73770 7976
rect 82170 7964 82176 7976
rect 82228 7964 82234 8016
rect 85574 7964 85580 8016
rect 85632 8004 85638 8016
rect 89686 8004 89714 8044
rect 118234 8032 118240 8044
rect 118292 8032 118298 8084
rect 133046 8032 133052 8084
rect 133104 8032 133110 8084
rect 160278 8032 160284 8084
rect 160336 8032 160342 8084
rect 162302 8032 162308 8084
rect 162360 8072 162366 8084
rect 162397 8075 162455 8081
rect 162397 8072 162409 8075
rect 162360 8044 162409 8072
rect 162360 8032 162366 8044
rect 162397 8041 162409 8044
rect 162443 8041 162455 8075
rect 162397 8035 162455 8041
rect 166350 8032 166356 8084
rect 166408 8032 166414 8084
rect 166810 8032 166816 8084
rect 166868 8072 166874 8084
rect 167089 8075 167147 8081
rect 167089 8072 167101 8075
rect 166868 8044 167101 8072
rect 166868 8032 166874 8044
rect 167089 8041 167101 8044
rect 167135 8041 167147 8075
rect 167089 8035 167147 8041
rect 167822 8032 167828 8084
rect 167880 8032 167886 8084
rect 168374 8032 168380 8084
rect 168432 8072 168438 8084
rect 169021 8075 169079 8081
rect 169021 8072 169033 8075
rect 168432 8044 169033 8072
rect 168432 8032 168438 8044
rect 169021 8041 169033 8044
rect 169067 8041 169079 8075
rect 169021 8035 169079 8041
rect 208394 8032 208400 8084
rect 208452 8072 208458 8084
rect 217962 8072 217968 8084
rect 208452 8044 217968 8072
rect 208452 8032 208458 8044
rect 217962 8032 217968 8044
rect 218020 8032 218026 8084
rect 225874 8032 225880 8084
rect 225932 8072 225938 8084
rect 225932 8044 226748 8072
rect 225932 8032 225938 8044
rect 85632 7976 89714 8004
rect 85632 7964 85638 7976
rect 93302 7964 93308 8016
rect 93360 7964 93366 8016
rect 99282 7964 99288 8016
rect 99340 8004 99346 8016
rect 99561 8007 99619 8013
rect 99561 8004 99573 8007
rect 99340 7976 99573 8004
rect 99340 7964 99346 7976
rect 99561 7973 99573 7976
rect 99607 7973 99619 8007
rect 99561 7967 99619 7973
rect 107930 7964 107936 8016
rect 107988 7964 107994 8016
rect 114922 7964 114928 8016
rect 114980 8004 114986 8016
rect 150894 8004 150900 8016
rect 114980 7976 150900 8004
rect 114980 7964 114986 7976
rect 150894 7964 150900 7976
rect 150952 7964 150958 8016
rect 152826 7964 152832 8016
rect 152884 8004 152890 8016
rect 162854 8004 162860 8016
rect 152884 7976 162860 8004
rect 152884 7964 152890 7976
rect 162854 7964 162860 7976
rect 162912 7964 162918 8016
rect 162946 7964 162952 8016
rect 163004 8004 163010 8016
rect 184566 8004 184572 8016
rect 163004 7976 184572 8004
rect 163004 7964 163010 7976
rect 184566 7964 184572 7976
rect 184624 7964 184630 8016
rect 221090 7964 221096 8016
rect 221148 8004 221154 8016
rect 226720 8004 226748 8044
rect 227622 8032 227628 8084
rect 227680 8072 227686 8084
rect 230382 8072 230388 8084
rect 227680 8044 230388 8072
rect 227680 8032 227686 8044
rect 230382 8032 230388 8044
rect 230440 8032 230446 8084
rect 230842 8032 230848 8084
rect 230900 8032 230906 8084
rect 243078 8032 243084 8084
rect 243136 8072 243142 8084
rect 243136 8044 258948 8072
rect 243136 8032 243142 8044
rect 236730 8004 236736 8016
rect 221148 7976 226656 8004
rect 226720 7976 236736 8004
rect 221148 7964 221154 7976
rect 14734 7896 14740 7948
rect 14792 7936 14798 7948
rect 45738 7936 45744 7948
rect 14792 7908 45744 7936
rect 14792 7896 14798 7908
rect 45738 7896 45744 7908
rect 45796 7896 45802 7948
rect 81894 7896 81900 7948
rect 81952 7936 81958 7948
rect 94958 7936 94964 7948
rect 81952 7908 94964 7936
rect 81952 7896 81958 7908
rect 94958 7896 94964 7908
rect 95016 7896 95022 7948
rect 99926 7896 99932 7948
rect 99984 7936 99990 7948
rect 100113 7939 100171 7945
rect 100113 7936 100125 7939
rect 99984 7908 100125 7936
rect 99984 7896 99990 7908
rect 100113 7905 100125 7908
rect 100159 7905 100171 7939
rect 100113 7899 100171 7905
rect 105170 7896 105176 7948
rect 105228 7896 105234 7948
rect 105449 7939 105507 7945
rect 105449 7905 105461 7939
rect 105495 7936 105507 7939
rect 106090 7936 106096 7948
rect 105495 7908 106096 7936
rect 105495 7905 105507 7908
rect 105449 7899 105507 7905
rect 106090 7896 106096 7908
rect 106148 7896 106154 7948
rect 107746 7896 107752 7948
rect 107804 7896 107810 7948
rect 141694 7896 141700 7948
rect 141752 7936 141758 7948
rect 152550 7936 152556 7948
rect 141752 7908 152556 7936
rect 141752 7896 141758 7908
rect 152550 7896 152556 7908
rect 152608 7896 152614 7948
rect 161382 7896 161388 7948
rect 161440 7896 161446 7948
rect 161658 7896 161664 7948
rect 161716 7936 161722 7948
rect 162670 7936 162676 7948
rect 161716 7908 162676 7936
rect 161716 7896 161722 7908
rect 162670 7896 162676 7908
rect 162728 7896 162734 7948
rect 163884 7908 165476 7936
rect 24949 7871 25007 7877
rect 24949 7837 24961 7871
rect 24995 7837 25007 7871
rect 24949 7831 25007 7837
rect 24964 7800 24992 7831
rect 25038 7828 25044 7880
rect 25096 7828 25102 7880
rect 26145 7871 26203 7877
rect 26145 7837 26157 7871
rect 26191 7868 26203 7871
rect 26602 7868 26608 7880
rect 26191 7840 26608 7868
rect 26191 7837 26203 7840
rect 26145 7831 26203 7837
rect 26602 7828 26608 7840
rect 26660 7828 26666 7880
rect 26697 7871 26755 7877
rect 26697 7837 26709 7871
rect 26743 7837 26755 7871
rect 26697 7831 26755 7837
rect 24964 7772 25636 7800
rect 25608 7741 25636 7772
rect 26234 7760 26240 7812
rect 26292 7800 26298 7812
rect 26712 7800 26740 7831
rect 27338 7828 27344 7880
rect 27396 7828 27402 7880
rect 27522 7828 27528 7880
rect 27580 7828 27586 7880
rect 28166 7828 28172 7880
rect 28224 7828 28230 7880
rect 28902 7828 28908 7880
rect 28960 7828 28966 7880
rect 29086 7828 29092 7880
rect 29144 7868 29150 7880
rect 52822 7868 52828 7880
rect 29144 7840 52828 7868
rect 29144 7828 29150 7840
rect 52822 7828 52828 7840
rect 52880 7828 52886 7880
rect 89533 7871 89591 7877
rect 89533 7837 89545 7871
rect 89579 7868 89591 7871
rect 90082 7868 90088 7880
rect 89579 7840 90088 7868
rect 89579 7837 89591 7840
rect 89533 7831 89591 7837
rect 90082 7828 90088 7840
rect 90140 7828 90146 7880
rect 93118 7828 93124 7880
rect 93176 7828 93182 7880
rect 99374 7828 99380 7880
rect 99432 7828 99438 7880
rect 105630 7877 105636 7880
rect 104529 7871 104587 7877
rect 104529 7868 104541 7871
rect 103808 7840 104541 7868
rect 26292 7772 26740 7800
rect 26292 7760 26298 7772
rect 26786 7760 26792 7812
rect 26844 7800 26850 7812
rect 51718 7800 51724 7812
rect 26844 7772 51724 7800
rect 26844 7760 26850 7772
rect 51718 7760 51724 7772
rect 51776 7760 51782 7812
rect 69842 7760 69848 7812
rect 69900 7800 69906 7812
rect 85666 7800 85672 7812
rect 69900 7772 85672 7800
rect 69900 7760 69906 7772
rect 85666 7760 85672 7772
rect 85724 7760 85730 7812
rect 25593 7735 25651 7741
rect 25593 7701 25605 7735
rect 25639 7732 25651 7735
rect 25682 7732 25688 7744
rect 25639 7704 25688 7732
rect 25639 7701 25651 7704
rect 25593 7695 25651 7701
rect 25682 7692 25688 7704
rect 25740 7692 25746 7744
rect 26510 7692 26516 7744
rect 26568 7732 26574 7744
rect 26881 7735 26939 7741
rect 26881 7732 26893 7735
rect 26568 7704 26893 7732
rect 26568 7692 26574 7704
rect 26881 7701 26893 7704
rect 26927 7701 26939 7735
rect 26881 7695 26939 7701
rect 27709 7735 27767 7741
rect 27709 7701 27721 7735
rect 27755 7732 27767 7735
rect 27798 7732 27804 7744
rect 27755 7704 27804 7732
rect 27755 7701 27767 7704
rect 27709 7695 27767 7701
rect 27798 7692 27804 7704
rect 27856 7692 27862 7744
rect 27890 7692 27896 7744
rect 27948 7732 27954 7744
rect 29089 7735 29147 7741
rect 29089 7732 29101 7735
rect 27948 7704 29101 7732
rect 27948 7692 27954 7704
rect 29089 7701 29101 7704
rect 29135 7701 29147 7735
rect 29089 7695 29147 7701
rect 89714 7692 89720 7744
rect 89772 7692 89778 7744
rect 94314 7692 94320 7744
rect 94372 7732 94378 7744
rect 103808 7741 103836 7840
rect 104529 7837 104541 7840
rect 104575 7837 104587 7871
rect 104529 7831 104587 7837
rect 104713 7871 104771 7877
rect 104713 7837 104725 7871
rect 104759 7837 104771 7871
rect 104713 7831 104771 7837
rect 105587 7871 105636 7877
rect 105587 7837 105599 7871
rect 105633 7837 105636 7871
rect 105587 7831 105636 7837
rect 103793 7735 103851 7741
rect 103793 7732 103805 7735
rect 94372 7704 103805 7732
rect 94372 7692 94378 7704
rect 103793 7701 103805 7704
rect 103839 7701 103851 7735
rect 103793 7695 103851 7701
rect 104158 7692 104164 7744
rect 104216 7732 104222 7744
rect 104728 7732 104756 7831
rect 105630 7828 105636 7831
rect 105688 7828 105694 7880
rect 105722 7828 105728 7880
rect 105780 7828 105786 7880
rect 107764 7868 107792 7896
rect 108945 7871 109003 7877
rect 108945 7868 108957 7871
rect 107764 7840 108957 7868
rect 108945 7837 108957 7840
rect 108991 7837 109003 7871
rect 108945 7831 109003 7837
rect 109773 7871 109831 7877
rect 109773 7837 109785 7871
rect 109819 7868 109831 7871
rect 109862 7868 109868 7880
rect 109819 7840 109868 7868
rect 109819 7837 109831 7840
rect 109773 7831 109831 7837
rect 106550 7800 106556 7812
rect 106292 7772 106556 7800
rect 104216 7704 104756 7732
rect 104216 7692 104222 7704
rect 105630 7692 105636 7744
rect 105688 7732 105694 7744
rect 106292 7732 106320 7772
rect 106550 7760 106556 7772
rect 106608 7760 106614 7812
rect 107749 7803 107807 7809
rect 107749 7769 107761 7803
rect 107795 7800 107807 7803
rect 108390 7800 108396 7812
rect 107795 7772 108396 7800
rect 107795 7769 107807 7772
rect 107749 7763 107807 7769
rect 108390 7760 108396 7772
rect 108448 7760 108454 7812
rect 108960 7800 108988 7831
rect 109862 7828 109868 7840
rect 109920 7828 109926 7880
rect 132862 7828 132868 7880
rect 132920 7828 132926 7880
rect 138658 7828 138664 7880
rect 138716 7868 138722 7880
rect 149054 7868 149060 7880
rect 138716 7840 149060 7868
rect 138716 7828 138722 7840
rect 149054 7828 149060 7840
rect 149112 7828 149118 7880
rect 149146 7828 149152 7880
rect 149204 7868 149210 7880
rect 158622 7868 158628 7880
rect 149204 7840 158628 7868
rect 149204 7828 149210 7840
rect 158622 7828 158628 7840
rect 158680 7828 158686 7880
rect 160094 7828 160100 7880
rect 160152 7828 160158 7880
rect 161572 7871 161630 7877
rect 161572 7837 161584 7871
rect 161618 7868 161630 7871
rect 161676 7868 161704 7896
rect 161618 7840 161704 7868
rect 161753 7871 161811 7877
rect 161618 7837 161630 7840
rect 161572 7831 161630 7837
rect 161753 7837 161765 7871
rect 161799 7868 161811 7871
rect 162213 7871 162271 7877
rect 162213 7868 162225 7871
rect 161799 7840 162225 7868
rect 161799 7837 161811 7840
rect 161753 7831 161811 7837
rect 162213 7837 162225 7840
rect 162259 7837 162271 7871
rect 162213 7831 162271 7837
rect 163774 7828 163780 7880
rect 163832 7828 163838 7880
rect 163884 7877 163912 7908
rect 163869 7871 163927 7877
rect 163869 7837 163881 7871
rect 163915 7837 163927 7871
rect 163869 7831 163927 7837
rect 164326 7828 164332 7880
rect 164384 7868 164390 7880
rect 164602 7868 164608 7880
rect 164384 7840 164608 7868
rect 164384 7828 164390 7840
rect 164602 7828 164608 7840
rect 164660 7828 164666 7880
rect 164712 7877 164740 7908
rect 165448 7880 165476 7908
rect 165614 7896 165620 7948
rect 165672 7936 165678 7948
rect 165672 7908 168972 7936
rect 165672 7896 165678 7908
rect 164697 7871 164755 7877
rect 164697 7837 164709 7871
rect 164743 7837 164755 7871
rect 164697 7831 164755 7837
rect 165338 7828 165344 7880
rect 165396 7828 165402 7880
rect 165430 7828 165436 7880
rect 165488 7868 165494 7880
rect 165525 7871 165583 7877
rect 165525 7868 165537 7871
rect 165488 7840 165537 7868
rect 165488 7828 165494 7840
rect 165525 7837 165537 7840
rect 165571 7837 165583 7871
rect 165525 7831 165583 7837
rect 166166 7828 166172 7880
rect 166224 7828 166230 7880
rect 166905 7871 166963 7877
rect 166905 7837 166917 7871
rect 166951 7868 166963 7871
rect 167454 7868 167460 7880
rect 166951 7840 167460 7868
rect 166951 7837 166963 7840
rect 166905 7831 166963 7837
rect 167454 7828 167460 7840
rect 167512 7828 167518 7880
rect 167638 7828 167644 7880
rect 167696 7828 167702 7880
rect 168834 7828 168840 7880
rect 168892 7828 168898 7880
rect 168944 7868 168972 7908
rect 169570 7896 169576 7948
rect 169628 7896 169634 7948
rect 187234 7936 187240 7948
rect 171106 7908 187240 7936
rect 171106 7868 171134 7908
rect 187234 7896 187240 7908
rect 187292 7896 187298 7948
rect 202785 7939 202843 7945
rect 202785 7905 202797 7939
rect 202831 7936 202843 7939
rect 203150 7936 203156 7948
rect 202831 7908 203156 7936
rect 202831 7905 202843 7908
rect 202785 7899 202843 7905
rect 203150 7896 203156 7908
rect 203208 7896 203214 7948
rect 216306 7896 216312 7948
rect 216364 7896 216370 7948
rect 218698 7896 218704 7948
rect 218756 7936 218762 7948
rect 223390 7936 223396 7948
rect 218756 7908 223396 7936
rect 218756 7896 218762 7908
rect 223390 7896 223396 7908
rect 223448 7896 223454 7948
rect 226628 7936 226656 7976
rect 236730 7964 236736 7976
rect 236788 7964 236794 8016
rect 237190 7964 237196 8016
rect 237248 8004 237254 8016
rect 239030 8004 239036 8016
rect 237248 7976 239036 8004
rect 237248 7964 237254 7976
rect 239030 7964 239036 7976
rect 239088 7964 239094 8016
rect 242894 7964 242900 8016
rect 242952 8004 242958 8016
rect 242952 7976 258304 8004
rect 242952 7964 242958 7976
rect 254026 7936 254032 7948
rect 226628 7908 254032 7936
rect 254026 7896 254032 7908
rect 254084 7896 254090 7948
rect 258276 7936 258304 7976
rect 258350 7964 258356 8016
rect 258408 7964 258414 8016
rect 258534 7936 258540 7948
rect 258276 7908 258540 7936
rect 258534 7896 258540 7908
rect 258592 7896 258598 7948
rect 168944 7840 171134 7868
rect 177206 7828 177212 7880
rect 177264 7868 177270 7880
rect 212442 7868 212448 7880
rect 177264 7840 212448 7868
rect 177264 7828 177270 7840
rect 212442 7828 212448 7840
rect 212500 7828 212506 7880
rect 214650 7828 214656 7880
rect 214708 7868 214714 7880
rect 215849 7871 215907 7877
rect 215849 7868 215861 7871
rect 214708 7840 215861 7868
rect 214708 7828 214714 7840
rect 215849 7837 215861 7840
rect 215895 7837 215907 7871
rect 215849 7831 215907 7837
rect 217781 7871 217839 7877
rect 217781 7837 217793 7871
rect 217827 7868 217839 7871
rect 219437 7871 219495 7877
rect 219437 7868 219449 7871
rect 217827 7840 219449 7868
rect 217827 7837 217839 7840
rect 217781 7831 217839 7837
rect 219437 7837 219449 7840
rect 219483 7868 219495 7871
rect 223574 7868 223580 7880
rect 219483 7840 223580 7868
rect 219483 7837 219495 7840
rect 219437 7831 219495 7837
rect 108960 7772 110000 7800
rect 105688 7704 106320 7732
rect 105688 7692 105694 7704
rect 106366 7692 106372 7744
rect 106424 7692 106430 7744
rect 108758 7692 108764 7744
rect 108816 7732 108822 7744
rect 109972 7741 110000 7772
rect 141602 7760 141608 7812
rect 141660 7800 141666 7812
rect 146478 7800 146484 7812
rect 141660 7772 146484 7800
rect 141660 7760 141666 7772
rect 146478 7760 146484 7772
rect 146536 7760 146542 7812
rect 146662 7760 146668 7812
rect 146720 7800 146726 7812
rect 174722 7800 174728 7812
rect 146720 7772 174728 7800
rect 146720 7760 146726 7772
rect 174722 7760 174728 7772
rect 174780 7760 174786 7812
rect 189258 7760 189264 7812
rect 189316 7800 189322 7812
rect 217796 7800 217824 7831
rect 223574 7828 223580 7840
rect 223632 7828 223638 7880
rect 226058 7868 226064 7880
rect 224788 7840 226064 7868
rect 189316 7772 217824 7800
rect 189316 7760 189322 7772
rect 217962 7760 217968 7812
rect 218020 7800 218026 7812
rect 218701 7803 218759 7809
rect 218701 7800 218713 7803
rect 218020 7772 218713 7800
rect 218020 7760 218026 7772
rect 218701 7769 218713 7772
rect 218747 7800 218759 7803
rect 224788 7800 224816 7840
rect 226058 7828 226064 7840
rect 226116 7828 226122 7880
rect 230566 7828 230572 7880
rect 230624 7868 230630 7880
rect 230661 7871 230719 7877
rect 230661 7868 230673 7871
rect 230624 7840 230673 7868
rect 230624 7828 230630 7840
rect 230661 7837 230673 7840
rect 230707 7837 230719 7871
rect 230661 7831 230719 7837
rect 235718 7828 235724 7880
rect 235776 7868 235782 7880
rect 235813 7871 235871 7877
rect 235813 7868 235825 7871
rect 235776 7840 235825 7868
rect 235776 7828 235782 7840
rect 235813 7837 235825 7840
rect 235859 7837 235871 7871
rect 235813 7831 235871 7837
rect 237006 7828 237012 7880
rect 237064 7828 237070 7880
rect 237101 7871 237159 7877
rect 237101 7837 237113 7871
rect 237147 7868 237159 7871
rect 237374 7868 237380 7880
rect 237147 7840 237380 7868
rect 237147 7837 237159 7840
rect 237101 7831 237159 7837
rect 237374 7828 237380 7840
rect 237432 7828 237438 7880
rect 237834 7828 237840 7880
rect 237892 7828 237898 7880
rect 237929 7871 237987 7877
rect 237929 7837 237941 7871
rect 237975 7868 237987 7871
rect 238018 7868 238024 7880
rect 237975 7840 238024 7868
rect 237975 7837 237987 7840
rect 237929 7831 237987 7837
rect 238018 7828 238024 7840
rect 238076 7828 238082 7880
rect 239398 7828 239404 7880
rect 239456 7868 239462 7880
rect 239456 7840 258764 7868
rect 239456 7828 239462 7840
rect 227622 7800 227628 7812
rect 218747 7772 224816 7800
rect 224926 7772 227628 7800
rect 218747 7769 218759 7772
rect 218701 7763 218759 7769
rect 109037 7735 109095 7741
rect 109037 7732 109049 7735
rect 108816 7704 109049 7732
rect 108816 7692 108822 7704
rect 109037 7701 109049 7704
rect 109083 7701 109095 7735
rect 109037 7695 109095 7701
rect 109957 7735 110015 7741
rect 109957 7701 109969 7735
rect 110003 7701 110015 7735
rect 109957 7695 110015 7701
rect 110506 7692 110512 7744
rect 110564 7732 110570 7744
rect 111886 7732 111892 7744
rect 110564 7704 111892 7732
rect 110564 7692 110570 7704
rect 111886 7692 111892 7704
rect 111944 7692 111950 7744
rect 143994 7692 144000 7744
rect 144052 7732 144058 7744
rect 146386 7732 146392 7744
rect 144052 7704 146392 7732
rect 144052 7692 144058 7704
rect 146386 7692 146392 7704
rect 146444 7692 146450 7744
rect 151446 7692 151452 7744
rect 151504 7732 151510 7744
rect 160002 7732 160008 7744
rect 151504 7704 160008 7732
rect 151504 7692 151510 7704
rect 160002 7692 160008 7704
rect 160060 7692 160066 7744
rect 163866 7692 163872 7744
rect 163924 7732 163930 7744
rect 164053 7735 164111 7741
rect 164053 7732 164065 7735
rect 163924 7704 164065 7732
rect 163924 7692 163930 7704
rect 164053 7701 164065 7704
rect 164099 7701 164111 7735
rect 164053 7695 164111 7701
rect 164602 7692 164608 7744
rect 164660 7732 164666 7744
rect 164881 7735 164939 7741
rect 164881 7732 164893 7735
rect 164660 7704 164893 7732
rect 164660 7692 164666 7704
rect 164881 7701 164893 7704
rect 164927 7701 164939 7735
rect 164881 7695 164939 7701
rect 165338 7692 165344 7744
rect 165396 7732 165402 7744
rect 165709 7735 165767 7741
rect 165709 7732 165721 7735
rect 165396 7704 165721 7732
rect 165396 7692 165402 7704
rect 165709 7701 165721 7704
rect 165755 7701 165767 7735
rect 165709 7695 165767 7701
rect 214190 7692 214196 7744
rect 214248 7732 214254 7744
rect 216398 7732 216404 7744
rect 214248 7704 216404 7732
rect 214248 7692 214254 7704
rect 216398 7692 216404 7704
rect 216456 7692 216462 7744
rect 216490 7692 216496 7744
rect 216548 7732 216554 7744
rect 217873 7735 217931 7741
rect 217873 7732 217885 7735
rect 216548 7704 217885 7732
rect 216548 7692 216554 7704
rect 217873 7701 217885 7704
rect 217919 7732 217931 7735
rect 218330 7732 218336 7744
rect 217919 7704 218336 7732
rect 217919 7701 217931 7704
rect 217873 7695 217931 7701
rect 218330 7692 218336 7704
rect 218388 7692 218394 7744
rect 218422 7692 218428 7744
rect 218480 7732 218486 7744
rect 218793 7735 218851 7741
rect 218793 7732 218805 7735
rect 218480 7704 218805 7732
rect 218480 7692 218486 7704
rect 218793 7701 218805 7704
rect 218839 7701 218851 7735
rect 218793 7695 218851 7701
rect 218974 7692 218980 7744
rect 219032 7732 219038 7744
rect 219529 7735 219587 7741
rect 219529 7732 219541 7735
rect 219032 7704 219541 7732
rect 219032 7692 219038 7704
rect 219529 7701 219541 7704
rect 219575 7701 219587 7735
rect 219529 7695 219587 7701
rect 219618 7692 219624 7744
rect 219676 7732 219682 7744
rect 224926 7732 224954 7772
rect 227622 7760 227628 7772
rect 227680 7760 227686 7812
rect 231210 7760 231216 7812
rect 231268 7800 231274 7812
rect 238113 7803 238171 7809
rect 238113 7800 238125 7803
rect 231268 7772 238125 7800
rect 231268 7760 231274 7772
rect 238113 7769 238125 7772
rect 238159 7769 238171 7803
rect 238113 7763 238171 7769
rect 258166 7760 258172 7812
rect 258224 7760 258230 7812
rect 219676 7704 224954 7732
rect 219676 7692 219682 7704
rect 228082 7692 228088 7744
rect 228140 7732 228146 7744
rect 236086 7732 236092 7744
rect 228140 7704 236092 7732
rect 228140 7692 228146 7704
rect 236086 7692 236092 7704
rect 236144 7692 236150 7744
rect 236178 7692 236184 7744
rect 236236 7732 236242 7744
rect 237285 7735 237343 7741
rect 237285 7732 237297 7735
rect 236236 7704 237297 7732
rect 236236 7692 236242 7704
rect 237285 7701 237297 7704
rect 237331 7701 237343 7735
rect 237285 7695 237343 7701
rect 237650 7692 237656 7744
rect 237708 7732 237714 7744
rect 242894 7732 242900 7744
rect 237708 7704 242900 7732
rect 237708 7692 237714 7704
rect 242894 7692 242900 7704
rect 242952 7692 242958 7744
rect 258736 7732 258764 7840
rect 258810 7828 258816 7880
rect 258868 7828 258874 7880
rect 258920 7800 258948 8044
rect 258994 8032 259000 8084
rect 259052 8032 259058 8084
rect 259641 8075 259699 8081
rect 259641 8041 259653 8075
rect 259687 8072 259699 8075
rect 259822 8072 259828 8084
rect 259687 8044 259828 8072
rect 259687 8041 259699 8044
rect 259641 8035 259699 8041
rect 259822 8032 259828 8044
rect 259880 8032 259886 8084
rect 260466 8032 260472 8084
rect 260524 8032 260530 8084
rect 268010 8072 268016 8084
rect 261680 8044 268016 8072
rect 261680 8004 261708 8044
rect 268010 8032 268016 8044
rect 268068 8032 268074 8084
rect 268102 8032 268108 8084
rect 268160 8072 268166 8084
rect 269669 8075 269727 8081
rect 269669 8072 269681 8075
rect 268160 8044 269681 8072
rect 268160 8032 268166 8044
rect 269669 8041 269681 8044
rect 269715 8041 269727 8075
rect 269669 8035 269727 8041
rect 259840 7976 261708 8004
rect 263566 7976 269344 8004
rect 259840 7877 259868 7976
rect 259914 7896 259920 7948
rect 259972 7936 259978 7948
rect 263566 7936 263594 7976
rect 259972 7908 263594 7936
rect 259972 7896 259978 7908
rect 264238 7896 264244 7948
rect 264296 7936 264302 7948
rect 268197 7939 268255 7945
rect 268197 7936 268209 7939
rect 264296 7908 268209 7936
rect 264296 7896 264302 7908
rect 268197 7905 268209 7908
rect 268243 7905 268255 7939
rect 268197 7899 268255 7905
rect 268657 7939 268715 7945
rect 268657 7905 268669 7939
rect 268703 7905 268715 7939
rect 268657 7899 268715 7905
rect 259825 7871 259883 7877
rect 259825 7837 259837 7871
rect 259871 7837 259883 7871
rect 259825 7831 259883 7837
rect 260282 7828 260288 7880
rect 260340 7828 260346 7880
rect 261846 7828 261852 7880
rect 261904 7828 261910 7880
rect 261938 7828 261944 7880
rect 261996 7828 262002 7880
rect 262582 7828 262588 7880
rect 262640 7828 262646 7880
rect 262769 7871 262827 7877
rect 262769 7837 262781 7871
rect 262815 7837 262827 7871
rect 262769 7831 262827 7837
rect 260834 7800 260840 7812
rect 258920 7772 260840 7800
rect 260834 7760 260840 7772
rect 260892 7760 260898 7812
rect 261956 7800 261984 7828
rect 262784 7800 262812 7831
rect 263134 7828 263140 7880
rect 263192 7868 263198 7880
rect 263413 7871 263471 7877
rect 263413 7868 263425 7871
rect 263192 7840 263425 7868
rect 263192 7828 263198 7840
rect 263413 7837 263425 7840
rect 263459 7837 263471 7871
rect 263413 7831 263471 7837
rect 263597 7871 263655 7877
rect 263597 7837 263609 7871
rect 263643 7868 263655 7871
rect 263778 7868 263784 7880
rect 263643 7840 263784 7868
rect 263643 7837 263655 7840
rect 263597 7831 263655 7837
rect 263612 7800 263640 7831
rect 263778 7828 263784 7840
rect 263836 7828 263842 7880
rect 264425 7871 264483 7877
rect 264425 7837 264437 7871
rect 264471 7868 264483 7871
rect 264977 7871 265035 7877
rect 264624 7868 264928 7870
rect 264471 7842 264928 7868
rect 264471 7840 264652 7842
rect 264471 7837 264483 7840
rect 264425 7831 264483 7837
rect 261956 7772 263640 7800
rect 260926 7732 260932 7744
rect 258736 7704 260932 7732
rect 260926 7692 260932 7704
rect 260984 7692 260990 7744
rect 262125 7735 262183 7741
rect 262125 7701 262137 7735
rect 262171 7732 262183 7735
rect 262306 7732 262312 7744
rect 262171 7704 262312 7732
rect 262171 7701 262183 7704
rect 262125 7695 262183 7701
rect 262306 7692 262312 7704
rect 262364 7692 262370 7744
rect 262953 7735 263011 7741
rect 262953 7701 262965 7735
rect 262999 7732 263011 7735
rect 263042 7732 263048 7744
rect 262999 7704 263048 7732
rect 262999 7701 263011 7704
rect 262953 7695 263011 7701
rect 263042 7692 263048 7704
rect 263100 7692 263106 7744
rect 263781 7735 263839 7741
rect 263781 7701 263793 7735
rect 263827 7732 263839 7735
rect 264146 7732 264152 7744
rect 263827 7704 264152 7732
rect 263827 7701 263839 7704
rect 263781 7695 263839 7701
rect 264146 7692 264152 7704
rect 264204 7692 264210 7744
rect 264238 7692 264244 7744
rect 264296 7692 264302 7744
rect 264900 7732 264928 7842
rect 264977 7837 264989 7871
rect 265023 7837 265035 7871
rect 264977 7831 265035 7837
rect 265069 7871 265127 7877
rect 265069 7837 265081 7871
rect 265115 7868 265127 7871
rect 265250 7868 265256 7880
rect 265115 7840 265256 7868
rect 265115 7837 265127 7840
rect 265069 7831 265127 7837
rect 264992 7800 265020 7831
rect 265250 7828 265256 7840
rect 265308 7828 265314 7880
rect 265802 7828 265808 7880
rect 265860 7828 265866 7880
rect 265897 7871 265955 7877
rect 265897 7837 265909 7871
rect 265943 7868 265955 7871
rect 265986 7868 265992 7880
rect 265943 7840 265992 7868
rect 265943 7837 265955 7840
rect 265897 7831 265955 7837
rect 265986 7828 265992 7840
rect 266044 7828 266050 7880
rect 267458 7828 267464 7880
rect 267516 7868 267522 7880
rect 267516 7840 268240 7868
rect 267516 7828 267522 7840
rect 266170 7800 266176 7812
rect 264992 7772 266176 7800
rect 266170 7760 266176 7772
rect 266228 7760 266234 7812
rect 267274 7760 267280 7812
rect 267332 7760 267338 7812
rect 267642 7760 267648 7812
rect 267700 7760 267706 7812
rect 268212 7800 268240 7840
rect 268286 7828 268292 7880
rect 268344 7828 268350 7880
rect 268562 7800 268568 7812
rect 268212 7772 268568 7800
rect 268562 7760 268568 7772
rect 268620 7760 268626 7812
rect 265066 7732 265072 7744
rect 264900 7704 265072 7732
rect 265066 7692 265072 7704
rect 265124 7692 265130 7744
rect 265253 7735 265311 7741
rect 265253 7701 265265 7735
rect 265299 7732 265311 7735
rect 265434 7732 265440 7744
rect 265299 7704 265440 7732
rect 265299 7701 265311 7704
rect 265253 7695 265311 7701
rect 265434 7692 265440 7704
rect 265492 7692 265498 7744
rect 266078 7692 266084 7744
rect 266136 7692 266142 7744
rect 267458 7692 267464 7744
rect 267516 7732 267522 7744
rect 268672 7732 268700 7899
rect 269022 7896 269028 7948
rect 269080 7936 269086 7948
rect 269209 7939 269267 7945
rect 269209 7936 269221 7939
rect 269080 7908 269221 7936
rect 269080 7896 269086 7908
rect 269209 7905 269221 7908
rect 269255 7905 269267 7939
rect 269209 7899 269267 7905
rect 269316 7877 269344 7976
rect 270129 7939 270187 7945
rect 270129 7905 270141 7939
rect 270175 7936 270187 7939
rect 271782 7936 271788 7948
rect 270175 7908 271788 7936
rect 270175 7905 270187 7908
rect 270129 7899 270187 7905
rect 271782 7896 271788 7908
rect 271840 7896 271846 7948
rect 269301 7871 269359 7877
rect 269301 7837 269313 7871
rect 269347 7837 269359 7871
rect 269301 7831 269359 7837
rect 270405 7871 270463 7877
rect 270405 7837 270417 7871
rect 270451 7837 270463 7871
rect 270405 7831 270463 7837
rect 268746 7760 268752 7812
rect 268804 7800 268810 7812
rect 270420 7800 270448 7831
rect 268804 7772 270448 7800
rect 268804 7760 268810 7772
rect 267516 7704 268700 7732
rect 267516 7692 267522 7704
rect 1104 7642 271651 7664
rect 1104 7590 68546 7642
rect 68598 7590 68610 7642
rect 68662 7590 68674 7642
rect 68726 7590 68738 7642
rect 68790 7590 68802 7642
rect 68854 7590 136143 7642
rect 136195 7590 136207 7642
rect 136259 7590 136271 7642
rect 136323 7590 136335 7642
rect 136387 7590 136399 7642
rect 136451 7590 203740 7642
rect 203792 7590 203804 7642
rect 203856 7590 203868 7642
rect 203920 7590 203932 7642
rect 203984 7590 203996 7642
rect 204048 7590 271337 7642
rect 271389 7590 271401 7642
rect 271453 7590 271465 7642
rect 271517 7590 271529 7642
rect 271581 7590 271593 7642
rect 271645 7590 271651 7642
rect 1104 7568 271651 7590
rect 25130 7488 25136 7540
rect 25188 7528 25194 7540
rect 25593 7531 25651 7537
rect 25593 7528 25605 7531
rect 25188 7500 25605 7528
rect 25188 7488 25194 7500
rect 25593 7497 25605 7500
rect 25639 7497 25651 7531
rect 25593 7491 25651 7497
rect 26418 7488 26424 7540
rect 26476 7488 26482 7540
rect 26602 7488 26608 7540
rect 26660 7528 26666 7540
rect 26660 7500 31754 7528
rect 26660 7488 26666 7500
rect 20346 7420 20352 7472
rect 20404 7460 20410 7472
rect 26786 7460 26792 7472
rect 20404 7432 26792 7460
rect 20404 7420 20410 7432
rect 26786 7420 26792 7432
rect 26844 7420 26850 7472
rect 31726 7460 31754 7500
rect 31846 7488 31852 7540
rect 31904 7528 31910 7540
rect 41966 7528 41972 7540
rect 31904 7500 41972 7528
rect 31904 7488 31910 7500
rect 41966 7488 41972 7500
rect 42024 7488 42030 7540
rect 66898 7488 66904 7540
rect 66956 7528 66962 7540
rect 67361 7531 67419 7537
rect 67361 7528 67373 7531
rect 66956 7500 67373 7528
rect 66956 7488 66962 7500
rect 67361 7497 67373 7500
rect 67407 7497 67419 7531
rect 67361 7491 67419 7497
rect 78214 7488 78220 7540
rect 78272 7528 78278 7540
rect 104158 7528 104164 7540
rect 78272 7500 104164 7528
rect 78272 7488 78278 7500
rect 104158 7488 104164 7500
rect 104216 7488 104222 7540
rect 109037 7531 109095 7537
rect 109037 7528 109049 7531
rect 106568 7500 109049 7528
rect 59814 7460 59820 7472
rect 31726 7432 59820 7460
rect 59814 7420 59820 7432
rect 59872 7460 59878 7472
rect 60366 7460 60372 7472
rect 59872 7432 60372 7460
rect 59872 7420 59878 7432
rect 60366 7420 60372 7432
rect 60424 7420 60430 7472
rect 77570 7420 77576 7472
rect 77628 7460 77634 7472
rect 94314 7460 94320 7472
rect 77628 7432 94320 7460
rect 77628 7420 77634 7432
rect 94314 7420 94320 7432
rect 94372 7420 94378 7472
rect 94406 7420 94412 7472
rect 94464 7460 94470 7472
rect 106093 7463 106151 7469
rect 106093 7460 106105 7463
rect 94464 7432 106105 7460
rect 94464 7420 94470 7432
rect 106093 7429 106105 7432
rect 106139 7460 106151 7463
rect 106139 7432 106504 7460
rect 106139 7429 106151 7432
rect 106093 7423 106151 7429
rect 24486 7352 24492 7404
rect 24544 7352 24550 7404
rect 25038 7352 25044 7404
rect 25096 7392 25102 7404
rect 25409 7395 25467 7401
rect 25409 7392 25421 7395
rect 25096 7364 25421 7392
rect 25096 7352 25102 7364
rect 25409 7361 25421 7364
rect 25455 7392 25467 7395
rect 26234 7392 26240 7404
rect 25455 7364 26240 7392
rect 25455 7361 25467 7364
rect 25409 7355 25467 7361
rect 26234 7352 26240 7364
rect 26292 7352 26298 7404
rect 27798 7352 27804 7404
rect 27856 7352 27862 7404
rect 42797 7395 42855 7401
rect 42797 7361 42809 7395
rect 42843 7392 42855 7395
rect 67545 7395 67603 7401
rect 42843 7364 43208 7392
rect 42843 7361 42855 7364
rect 42797 7355 42855 7361
rect 25222 7284 25228 7336
rect 25280 7284 25286 7336
rect 26050 7284 26056 7336
rect 26108 7284 26114 7336
rect 23382 7216 23388 7268
rect 23440 7256 23446 7268
rect 28534 7256 28540 7268
rect 23440 7228 28540 7256
rect 23440 7216 23446 7228
rect 28534 7216 28540 7228
rect 28592 7216 28598 7268
rect 36998 7216 37004 7268
rect 37056 7256 37062 7268
rect 43180 7265 43208 7364
rect 67545 7361 67557 7395
rect 67591 7392 67603 7395
rect 79410 7392 79416 7404
rect 67591 7364 79416 7392
rect 67591 7361 67603 7364
rect 67545 7355 67603 7361
rect 79410 7352 79416 7364
rect 79468 7352 79474 7404
rect 84166 7364 96614 7392
rect 80146 7284 80152 7336
rect 80204 7324 80210 7336
rect 84166 7324 84194 7364
rect 80204 7296 84194 7324
rect 96586 7324 96614 7364
rect 100202 7352 100208 7404
rect 100260 7352 100266 7404
rect 106476 7401 106504 7432
rect 106461 7395 106519 7401
rect 106461 7361 106473 7395
rect 106507 7361 106519 7395
rect 106461 7355 106519 7361
rect 106568 7324 106596 7500
rect 109037 7497 109049 7500
rect 109083 7528 109095 7531
rect 111705 7531 111763 7537
rect 111705 7528 111717 7531
rect 109083 7500 109632 7528
rect 109083 7497 109095 7500
rect 109037 7491 109095 7497
rect 107378 7352 107384 7404
rect 107436 7352 107442 7404
rect 108390 7352 108396 7404
rect 108448 7352 108454 7404
rect 109604 7401 109632 7500
rect 109788 7500 111717 7528
rect 109788 7401 109816 7500
rect 111705 7497 111717 7500
rect 111751 7497 111763 7531
rect 111705 7491 111763 7497
rect 121181 7531 121239 7537
rect 121181 7497 121193 7531
rect 121227 7528 121239 7531
rect 121454 7528 121460 7540
rect 121227 7500 121460 7528
rect 121227 7497 121239 7500
rect 121181 7491 121239 7497
rect 121454 7488 121460 7500
rect 121512 7488 121518 7540
rect 146294 7528 146300 7540
rect 145668 7500 146300 7528
rect 109589 7395 109647 7401
rect 109589 7361 109601 7395
rect 109635 7361 109647 7395
rect 109589 7355 109647 7361
rect 109773 7395 109831 7401
rect 109773 7361 109785 7395
rect 109819 7361 109831 7395
rect 109773 7355 109831 7361
rect 96586 7296 106596 7324
rect 106645 7327 106703 7333
rect 80204 7284 80210 7296
rect 106645 7293 106657 7327
rect 106691 7324 106703 7327
rect 106826 7324 106832 7336
rect 106691 7296 106832 7324
rect 106691 7293 106703 7296
rect 106645 7287 106703 7293
rect 106826 7284 106832 7296
rect 106884 7284 106890 7336
rect 107562 7333 107568 7336
rect 107519 7327 107568 7333
rect 107519 7293 107531 7327
rect 107565 7293 107568 7327
rect 107519 7287 107568 7293
rect 107562 7284 107568 7287
rect 107620 7284 107626 7336
rect 107657 7327 107715 7333
rect 107657 7293 107669 7327
rect 107703 7324 107715 7327
rect 107838 7324 107844 7336
rect 107703 7296 107844 7324
rect 107703 7293 107715 7296
rect 107657 7287 107715 7293
rect 107838 7284 107844 7296
rect 107896 7284 107902 7336
rect 109788 7324 109816 7355
rect 110506 7352 110512 7404
rect 110564 7352 110570 7404
rect 112070 7352 112076 7404
rect 112128 7352 112134 7404
rect 120258 7352 120264 7404
rect 120316 7392 120322 7404
rect 145668 7401 145696 7500
rect 146294 7488 146300 7500
rect 146352 7488 146358 7540
rect 146754 7488 146760 7540
rect 146812 7528 146818 7540
rect 155586 7528 155592 7540
rect 146812 7500 155592 7528
rect 146812 7488 146818 7500
rect 155586 7488 155592 7500
rect 155644 7488 155650 7540
rect 161290 7488 161296 7540
rect 161348 7488 161354 7540
rect 162578 7488 162584 7540
rect 162636 7488 162642 7540
rect 162670 7488 162676 7540
rect 162728 7528 162734 7540
rect 163317 7531 163375 7537
rect 163317 7528 163329 7531
rect 162728 7500 163329 7528
rect 162728 7488 162734 7500
rect 163317 7497 163329 7500
rect 163363 7497 163375 7531
rect 163317 7491 163375 7497
rect 164050 7488 164056 7540
rect 164108 7488 164114 7540
rect 164786 7488 164792 7540
rect 164844 7488 164850 7540
rect 165522 7488 165528 7540
rect 165580 7488 165586 7540
rect 168282 7488 168288 7540
rect 168340 7528 168346 7540
rect 218698 7528 218704 7540
rect 168340 7500 218704 7528
rect 168340 7488 168346 7500
rect 218698 7488 218704 7500
rect 218756 7488 218762 7540
rect 220357 7531 220415 7537
rect 220357 7497 220369 7531
rect 220403 7528 220415 7531
rect 221458 7528 221464 7540
rect 220403 7500 221464 7528
rect 220403 7497 220415 7500
rect 220357 7491 220415 7497
rect 221458 7488 221464 7500
rect 221516 7528 221522 7540
rect 236914 7528 236920 7540
rect 221516 7500 236920 7528
rect 221516 7488 221522 7500
rect 236914 7488 236920 7500
rect 236972 7488 236978 7540
rect 237190 7488 237196 7540
rect 237248 7528 237254 7540
rect 238938 7528 238944 7540
rect 237248 7500 238944 7528
rect 237248 7488 237254 7500
rect 238938 7488 238944 7500
rect 238996 7488 239002 7540
rect 259641 7531 259699 7537
rect 259641 7497 259653 7531
rect 259687 7528 259699 7531
rect 259914 7528 259920 7540
rect 259687 7500 259920 7528
rect 259687 7497 259699 7500
rect 259641 7491 259699 7497
rect 259914 7488 259920 7500
rect 259972 7488 259978 7540
rect 260285 7531 260343 7537
rect 260285 7497 260297 7531
rect 260331 7528 260343 7531
rect 260374 7528 260380 7540
rect 260331 7500 260380 7528
rect 260331 7497 260343 7500
rect 260285 7491 260343 7497
rect 260374 7488 260380 7500
rect 260432 7488 260438 7540
rect 261754 7488 261760 7540
rect 261812 7488 261818 7540
rect 262490 7488 262496 7540
rect 262548 7488 262554 7540
rect 263226 7488 263232 7540
rect 263284 7488 263290 7540
rect 264330 7488 264336 7540
rect 264388 7488 264394 7540
rect 265897 7531 265955 7537
rect 265897 7497 265909 7531
rect 265943 7528 265955 7531
rect 270678 7528 270684 7540
rect 265943 7500 270684 7528
rect 265943 7497 265955 7500
rect 265897 7491 265955 7497
rect 270678 7488 270684 7500
rect 270736 7488 270742 7540
rect 152366 7460 152372 7472
rect 151188 7432 152372 7460
rect 146754 7401 146760 7404
rect 121365 7395 121423 7401
rect 121365 7392 121377 7395
rect 120316 7364 121377 7392
rect 120316 7352 120322 7364
rect 121365 7361 121377 7364
rect 121411 7361 121423 7395
rect 121365 7355 121423 7361
rect 145653 7395 145711 7401
rect 145653 7361 145665 7395
rect 145699 7361 145711 7395
rect 145653 7355 145711 7361
rect 146711 7395 146760 7401
rect 146711 7361 146723 7395
rect 146757 7361 146760 7395
rect 146711 7355 146760 7361
rect 146754 7352 146760 7355
rect 146812 7352 146818 7404
rect 151188 7401 151216 7432
rect 152366 7420 152372 7432
rect 152424 7420 152430 7472
rect 152550 7420 152556 7472
rect 152608 7460 152614 7472
rect 168190 7460 168196 7472
rect 152608 7432 168196 7460
rect 152608 7420 152614 7432
rect 168190 7420 168196 7432
rect 168248 7420 168254 7472
rect 217962 7460 217968 7472
rect 216416 7432 217968 7460
rect 216416 7404 216444 7432
rect 217962 7420 217968 7432
rect 218020 7420 218026 7472
rect 226978 7420 226984 7472
rect 227036 7460 227042 7472
rect 251358 7460 251364 7472
rect 227036 7432 251364 7460
rect 227036 7420 227042 7432
rect 251358 7420 251364 7432
rect 251416 7420 251422 7472
rect 268010 7460 268016 7472
rect 261128 7432 268016 7460
rect 151173 7395 151231 7401
rect 151173 7361 151185 7395
rect 151219 7361 151231 7395
rect 151173 7355 151231 7361
rect 152568 7364 157334 7392
rect 110626 7327 110684 7333
rect 110626 7324 110638 7327
rect 108040 7296 109816 7324
rect 110340 7296 110638 7324
rect 42613 7259 42671 7265
rect 42613 7256 42625 7259
rect 37056 7228 42625 7256
rect 37056 7216 37062 7228
rect 42613 7225 42625 7228
rect 42659 7225 42671 7259
rect 42613 7219 42671 7225
rect 43165 7259 43223 7265
rect 43165 7225 43177 7259
rect 43211 7256 43223 7259
rect 43211 7228 74534 7256
rect 43211 7225 43223 7228
rect 43165 7219 43223 7225
rect 23474 7148 23480 7200
rect 23532 7188 23538 7200
rect 24673 7191 24731 7197
rect 24673 7188 24685 7191
rect 23532 7160 24685 7188
rect 23532 7148 23538 7160
rect 24673 7157 24685 7160
rect 24719 7157 24731 7191
rect 24673 7151 24731 7157
rect 26234 7148 26240 7200
rect 26292 7188 26298 7200
rect 27985 7191 28043 7197
rect 27985 7188 27997 7191
rect 26292 7160 27997 7188
rect 26292 7148 26298 7160
rect 27985 7157 27997 7160
rect 28031 7157 28043 7191
rect 74506 7188 74534 7228
rect 78858 7216 78864 7268
rect 78916 7256 78922 7268
rect 94406 7256 94412 7268
rect 78916 7228 94412 7256
rect 78916 7216 78922 7228
rect 94406 7216 94412 7228
rect 94464 7216 94470 7268
rect 99346 7228 100156 7256
rect 79594 7188 79600 7200
rect 74506 7160 79600 7188
rect 27985 7151 28043 7157
rect 79594 7148 79600 7160
rect 79652 7148 79658 7200
rect 80146 7148 80152 7200
rect 80204 7188 80210 7200
rect 99346 7188 99374 7228
rect 80204 7160 99374 7188
rect 80204 7148 80210 7160
rect 100018 7148 100024 7200
rect 100076 7148 100082 7200
rect 100128 7188 100156 7228
rect 105170 7216 105176 7268
rect 105228 7256 105234 7268
rect 107102 7256 107108 7268
rect 105228 7228 107108 7256
rect 105228 7216 105234 7228
rect 107102 7216 107108 7228
rect 107160 7216 107166 7268
rect 108040 7188 108068 7296
rect 108301 7259 108359 7265
rect 108301 7225 108313 7259
rect 108347 7256 108359 7259
rect 109126 7256 109132 7268
rect 108347 7228 109132 7256
rect 108347 7225 108359 7228
rect 108301 7219 108359 7225
rect 109126 7216 109132 7228
rect 109184 7216 109190 7268
rect 110230 7216 110236 7268
rect 110288 7216 110294 7268
rect 100128 7160 108068 7188
rect 108574 7148 108580 7200
rect 108632 7148 108638 7200
rect 110340 7188 110368 7296
rect 110626 7293 110638 7296
rect 110672 7293 110684 7327
rect 110626 7287 110684 7293
rect 110785 7327 110843 7333
rect 110785 7293 110797 7327
rect 110831 7324 110843 7327
rect 110966 7324 110972 7336
rect 110831 7296 110972 7324
rect 110831 7293 110843 7296
rect 110785 7287 110843 7293
rect 110966 7284 110972 7296
rect 111024 7284 111030 7336
rect 112622 7284 112628 7336
rect 112680 7284 112686 7336
rect 145837 7327 145895 7333
rect 145837 7293 145849 7327
rect 145883 7324 145895 7327
rect 146573 7327 146631 7333
rect 146573 7324 146585 7327
rect 145883 7296 146156 7324
rect 145883 7293 145895 7296
rect 145837 7287 145895 7293
rect 146128 7268 146156 7296
rect 146404 7296 146585 7324
rect 111429 7259 111487 7265
rect 111429 7225 111441 7259
rect 111475 7256 111487 7259
rect 112438 7256 112444 7268
rect 111475 7228 112444 7256
rect 111475 7225 111487 7228
rect 111429 7219 111487 7225
rect 112438 7216 112444 7228
rect 112496 7216 112502 7268
rect 146110 7216 146116 7268
rect 146168 7216 146174 7268
rect 146294 7216 146300 7268
rect 146352 7216 146358 7268
rect 113082 7188 113088 7200
rect 110340 7160 113088 7188
rect 113082 7148 113088 7160
rect 113140 7148 113146 7200
rect 146404 7188 146432 7296
rect 146573 7293 146585 7296
rect 146619 7293 146631 7327
rect 146573 7287 146631 7293
rect 146849 7327 146907 7333
rect 146849 7293 146861 7327
rect 146895 7324 146907 7327
rect 147030 7324 147036 7336
rect 146895 7296 147036 7324
rect 146895 7293 146907 7296
rect 146849 7287 146907 7293
rect 147030 7284 147036 7296
rect 147088 7284 147094 7336
rect 150986 7284 150992 7336
rect 151044 7324 151050 7336
rect 151357 7327 151415 7333
rect 151357 7324 151369 7327
rect 151044 7296 151369 7324
rect 151044 7284 151050 7296
rect 151357 7293 151369 7296
rect 151403 7293 151415 7327
rect 151357 7287 151415 7293
rect 147861 7259 147919 7265
rect 147861 7256 147873 7259
rect 147232 7228 147873 7256
rect 147232 7188 147260 7228
rect 147861 7225 147873 7228
rect 147907 7256 147919 7259
rect 152568 7256 152596 7364
rect 153013 7327 153071 7333
rect 153013 7293 153025 7327
rect 153059 7293 153071 7327
rect 153013 7287 153071 7293
rect 147907 7228 152596 7256
rect 147907 7225 147919 7228
rect 147861 7219 147919 7225
rect 146404 7160 147260 7188
rect 147490 7148 147496 7200
rect 147548 7148 147554 7200
rect 150894 7148 150900 7200
rect 150952 7188 150958 7200
rect 153028 7188 153056 7287
rect 157306 7256 157334 7364
rect 161106 7352 161112 7404
rect 161164 7352 161170 7404
rect 162394 7352 162400 7404
rect 162452 7352 162458 7404
rect 163225 7395 163283 7401
rect 163225 7361 163237 7395
rect 163271 7361 163283 7395
rect 163225 7355 163283 7361
rect 158622 7284 158628 7336
rect 158680 7324 158686 7336
rect 162946 7324 162952 7336
rect 158680 7296 162952 7324
rect 158680 7284 158686 7296
rect 162946 7284 162952 7296
rect 163004 7284 163010 7336
rect 163240 7324 163268 7355
rect 163866 7352 163872 7404
rect 163924 7352 163930 7404
rect 164602 7352 164608 7404
rect 164660 7352 164666 7404
rect 165338 7352 165344 7404
rect 165396 7352 165402 7404
rect 169297 7395 169355 7401
rect 169297 7361 169309 7395
rect 169343 7392 169355 7395
rect 169754 7392 169760 7404
rect 169343 7364 169760 7392
rect 169343 7361 169355 7364
rect 169297 7355 169355 7361
rect 169754 7352 169760 7364
rect 169812 7352 169818 7404
rect 214101 7395 214159 7401
rect 214101 7361 214113 7395
rect 214147 7392 214159 7395
rect 214147 7364 214328 7392
rect 214147 7361 214159 7364
rect 214101 7355 214159 7361
rect 165154 7324 165160 7336
rect 163240 7296 165160 7324
rect 165154 7284 165160 7296
rect 165212 7284 165218 7336
rect 172514 7284 172520 7336
rect 172572 7324 172578 7336
rect 214190 7324 214196 7336
rect 172572 7296 214196 7324
rect 172572 7284 172578 7296
rect 214190 7284 214196 7296
rect 214248 7284 214254 7336
rect 181162 7256 181168 7268
rect 157306 7228 181168 7256
rect 181162 7216 181168 7228
rect 181220 7216 181226 7268
rect 213914 7216 213920 7268
rect 213972 7256 213978 7268
rect 214300 7256 214328 7364
rect 214466 7352 214472 7404
rect 214524 7352 214530 7404
rect 215570 7401 215576 7404
rect 215527 7395 215576 7401
rect 215527 7361 215539 7395
rect 215573 7361 215576 7395
rect 215527 7355 215576 7361
rect 215570 7352 215576 7355
rect 215628 7352 215634 7404
rect 216398 7352 216404 7404
rect 216456 7352 216462 7404
rect 216674 7352 216680 7404
rect 216732 7392 216738 7404
rect 217781 7395 217839 7401
rect 217781 7392 217793 7395
rect 216732 7364 217793 7392
rect 216732 7352 216738 7364
rect 217781 7361 217793 7364
rect 217827 7361 217839 7395
rect 217781 7355 217839 7361
rect 218698 7352 218704 7404
rect 218756 7352 218762 7404
rect 218974 7352 218980 7404
rect 219032 7352 219038 7404
rect 220354 7352 220360 7404
rect 220412 7392 220418 7404
rect 220541 7395 220599 7401
rect 220541 7392 220553 7395
rect 220412 7364 220553 7392
rect 220412 7352 220418 7364
rect 220541 7361 220553 7364
rect 220587 7361 220599 7395
rect 220541 7355 220599 7361
rect 221458 7352 221464 7404
rect 221516 7352 221522 7404
rect 221550 7352 221556 7404
rect 221608 7401 221614 7404
rect 221608 7395 221636 7401
rect 221624 7361 221636 7395
rect 221608 7355 221636 7361
rect 221608 7352 221614 7355
rect 221734 7352 221740 7404
rect 221792 7352 221798 7404
rect 222838 7352 222844 7404
rect 222896 7392 222902 7404
rect 222933 7395 222991 7401
rect 222933 7392 222945 7395
rect 222896 7364 222945 7392
rect 222896 7352 222902 7364
rect 222933 7361 222945 7364
rect 222979 7361 222991 7395
rect 222933 7355 222991 7361
rect 223850 7352 223856 7404
rect 223908 7352 223914 7404
rect 229741 7395 229799 7401
rect 229741 7361 229753 7395
rect 229787 7392 229799 7395
rect 230106 7392 230112 7404
rect 229787 7364 230112 7392
rect 229787 7361 229799 7364
rect 229741 7355 229799 7361
rect 230106 7352 230112 7364
rect 230164 7352 230170 7404
rect 230290 7352 230296 7404
rect 230348 7352 230354 7404
rect 231210 7352 231216 7404
rect 231268 7352 231274 7404
rect 231302 7352 231308 7404
rect 231360 7392 231366 7404
rect 232409 7395 232467 7401
rect 232409 7392 232421 7395
rect 231360 7364 232421 7392
rect 231360 7352 231366 7364
rect 232409 7361 232421 7364
rect 232455 7361 232467 7395
rect 232409 7355 232467 7361
rect 232593 7395 232651 7401
rect 232593 7361 232605 7395
rect 232639 7392 232651 7395
rect 235258 7392 235264 7404
rect 232639 7364 235264 7392
rect 232639 7361 232651 7364
rect 232593 7355 232651 7361
rect 235258 7352 235264 7364
rect 235316 7352 235322 7404
rect 235350 7352 235356 7404
rect 235408 7352 235414 7404
rect 235445 7395 235503 7401
rect 235445 7361 235457 7395
rect 235491 7392 235503 7395
rect 235994 7392 236000 7404
rect 235491 7364 236000 7392
rect 235491 7361 235503 7364
rect 235445 7355 235503 7361
rect 235994 7352 236000 7364
rect 236052 7352 236058 7404
rect 236178 7352 236184 7404
rect 236236 7352 236242 7404
rect 237282 7352 237288 7404
rect 237340 7352 237346 7404
rect 237374 7352 237380 7404
rect 237432 7392 237438 7404
rect 237469 7395 237527 7401
rect 237469 7392 237481 7395
rect 237432 7364 237481 7392
rect 237432 7352 237438 7364
rect 237469 7361 237481 7364
rect 237515 7392 237527 7395
rect 238018 7392 238024 7404
rect 237515 7364 238024 7392
rect 237515 7361 237527 7364
rect 237469 7355 237527 7361
rect 238018 7352 238024 7364
rect 238076 7392 238082 7404
rect 238573 7395 238631 7401
rect 238573 7392 238585 7395
rect 238076 7364 238585 7392
rect 238076 7352 238082 7364
rect 238573 7361 238585 7364
rect 238619 7392 238631 7395
rect 238662 7392 238668 7404
rect 238619 7364 238668 7392
rect 238619 7361 238631 7364
rect 238573 7355 238631 7361
rect 238662 7352 238668 7364
rect 238720 7352 238726 7404
rect 261128 7401 261156 7432
rect 268010 7420 268016 7432
rect 268068 7420 268074 7472
rect 268749 7463 268807 7469
rect 268749 7460 268761 7463
rect 268120 7432 268761 7460
rect 259825 7395 259883 7401
rect 259825 7361 259837 7395
rect 259871 7361 259883 7395
rect 259825 7355 259883 7361
rect 260469 7395 260527 7401
rect 260469 7361 260481 7395
rect 260515 7361 260527 7395
rect 260469 7355 260527 7361
rect 261113 7395 261171 7401
rect 261113 7361 261125 7395
rect 261159 7361 261171 7395
rect 261113 7355 261171 7361
rect 214653 7327 214711 7333
rect 214653 7293 214665 7327
rect 214699 7324 214711 7327
rect 215018 7324 215024 7336
rect 214699 7296 215024 7324
rect 214699 7293 214711 7296
rect 214653 7287 214711 7293
rect 215018 7284 215024 7296
rect 215076 7284 215082 7336
rect 215110 7284 215116 7336
rect 215168 7284 215174 7336
rect 215389 7327 215447 7333
rect 215389 7324 215401 7327
rect 215220 7296 215401 7324
rect 214834 7256 214840 7268
rect 213972 7228 214236 7256
rect 214300 7228 214840 7256
rect 213972 7216 213978 7228
rect 153381 7191 153439 7197
rect 153381 7188 153393 7191
rect 150952 7160 153393 7188
rect 150952 7148 150958 7160
rect 153381 7157 153393 7160
rect 153427 7188 153439 7191
rect 156046 7188 156052 7200
rect 153427 7160 156052 7188
rect 153427 7157 153439 7160
rect 153381 7151 153439 7157
rect 156046 7148 156052 7160
rect 156104 7148 156110 7200
rect 159266 7148 159272 7200
rect 159324 7188 159330 7200
rect 165614 7188 165620 7200
rect 159324 7160 165620 7188
rect 159324 7148 159330 7160
rect 165614 7148 165620 7160
rect 165672 7148 165678 7200
rect 169110 7148 169116 7200
rect 169168 7148 169174 7200
rect 206922 7148 206928 7200
rect 206980 7188 206986 7200
rect 212350 7188 212356 7200
rect 206980 7160 212356 7188
rect 206980 7148 206986 7160
rect 212350 7148 212356 7160
rect 212408 7148 212414 7200
rect 214208 7188 214236 7228
rect 214834 7216 214840 7228
rect 214892 7256 214898 7268
rect 215220 7256 215248 7296
rect 215389 7293 215401 7296
rect 215435 7293 215447 7327
rect 215389 7287 215447 7293
rect 215665 7327 215723 7333
rect 215665 7293 215677 7327
rect 215711 7324 215723 7327
rect 215711 7296 216444 7324
rect 215711 7293 215723 7296
rect 215665 7287 215723 7293
rect 216416 7268 216444 7296
rect 216582 7284 216588 7336
rect 216640 7284 216646 7336
rect 216950 7284 216956 7336
rect 217008 7324 217014 7336
rect 217965 7327 218023 7333
rect 217965 7324 217977 7327
rect 217008 7296 217977 7324
rect 217008 7284 217014 7296
rect 217965 7293 217977 7296
rect 218011 7293 218023 7327
rect 218716 7324 218744 7352
rect 217965 7287 218023 7293
rect 218348 7296 218744 7324
rect 218839 7327 218897 7333
rect 214892 7228 215248 7256
rect 214892 7216 214898 7228
rect 216398 7216 216404 7268
rect 216456 7216 216462 7268
rect 217229 7259 217287 7265
rect 217229 7225 217241 7259
rect 217275 7256 217287 7259
rect 218348 7256 218376 7296
rect 218839 7293 218851 7327
rect 218885 7324 218897 7327
rect 218885 7296 220032 7324
rect 218885 7293 218897 7296
rect 218839 7287 218897 7293
rect 220004 7268 220032 7296
rect 220722 7284 220728 7336
rect 220780 7284 220786 7336
rect 221200 7296 223068 7324
rect 217275 7228 218376 7256
rect 217275 7225 217287 7228
rect 217229 7219 217287 7225
rect 218422 7216 218428 7268
rect 218480 7216 218486 7268
rect 219986 7216 219992 7268
rect 220044 7216 220050 7268
rect 220538 7216 220544 7268
rect 220596 7256 220602 7268
rect 221200 7265 221228 7296
rect 221185 7259 221243 7265
rect 221185 7256 221197 7259
rect 220596 7228 221197 7256
rect 220596 7216 220602 7228
rect 221185 7225 221197 7228
rect 221231 7225 221243 7259
rect 223040 7256 223068 7296
rect 223114 7284 223120 7336
rect 223172 7284 223178 7336
rect 223942 7284 223948 7336
rect 224000 7333 224006 7336
rect 224000 7327 224028 7333
rect 224016 7293 224028 7327
rect 224000 7287 224028 7293
rect 224000 7284 224006 7287
rect 224126 7284 224132 7336
rect 224184 7284 224190 7336
rect 224954 7284 224960 7336
rect 225012 7324 225018 7336
rect 225141 7327 225199 7333
rect 225141 7324 225153 7327
rect 225012 7296 225153 7324
rect 225012 7284 225018 7296
rect 225141 7293 225153 7296
rect 225187 7324 225199 7327
rect 230308 7324 230336 7352
rect 231489 7327 231547 7333
rect 231489 7324 231501 7327
rect 225187 7296 226932 7324
rect 230308 7296 231501 7324
rect 225187 7293 225199 7296
rect 225141 7287 225199 7293
rect 223298 7256 223304 7268
rect 221185 7219 221243 7225
rect 222166 7228 222516 7256
rect 223040 7228 223304 7256
rect 216309 7191 216367 7197
rect 216309 7188 216321 7191
rect 214208 7160 216321 7188
rect 216309 7157 216321 7160
rect 216355 7157 216367 7191
rect 216309 7151 216367 7157
rect 218054 7148 218060 7200
rect 218112 7188 218118 7200
rect 219621 7191 219679 7197
rect 219621 7188 219633 7191
rect 218112 7160 219633 7188
rect 218112 7148 218118 7160
rect 219621 7157 219633 7160
rect 219667 7157 219679 7191
rect 219621 7151 219679 7157
rect 219710 7148 219716 7200
rect 219768 7188 219774 7200
rect 222166 7188 222194 7228
rect 219768 7160 222194 7188
rect 219768 7148 219774 7160
rect 222378 7148 222384 7200
rect 222436 7148 222442 7200
rect 222488 7188 222516 7228
rect 223298 7216 223304 7228
rect 223356 7256 223362 7268
rect 223577 7259 223635 7265
rect 223577 7256 223589 7259
rect 223356 7228 223589 7256
rect 223356 7216 223362 7228
rect 223577 7225 223589 7228
rect 223623 7225 223635 7259
rect 223577 7219 223635 7225
rect 224773 7259 224831 7265
rect 224773 7225 224785 7259
rect 224819 7256 224831 7259
rect 225506 7256 225512 7268
rect 224819 7228 225512 7256
rect 224819 7225 224831 7228
rect 224773 7219 224831 7225
rect 225506 7216 225512 7228
rect 225564 7216 225570 7268
rect 226904 7256 226932 7296
rect 231489 7293 231501 7296
rect 231535 7293 231547 7327
rect 231489 7287 231547 7293
rect 236086 7284 236092 7336
rect 236144 7324 236150 7336
rect 236457 7327 236515 7333
rect 236457 7324 236469 7327
rect 236144 7296 236469 7324
rect 236144 7284 236150 7296
rect 236457 7293 236469 7296
rect 236503 7293 236515 7327
rect 236457 7287 236515 7293
rect 238389 7327 238447 7333
rect 238389 7293 238401 7327
rect 238435 7324 238447 7327
rect 239122 7324 239128 7336
rect 238435 7296 239128 7324
rect 238435 7293 238447 7296
rect 238389 7287 238447 7293
rect 239122 7284 239128 7296
rect 239180 7284 239186 7336
rect 256786 7324 256792 7336
rect 248386 7296 256792 7324
rect 248386 7256 248414 7296
rect 256786 7284 256792 7296
rect 256844 7284 256850 7336
rect 226904 7228 248414 7256
rect 259840 7256 259868 7355
rect 260484 7324 260512 7355
rect 261570 7352 261576 7404
rect 261628 7352 261634 7404
rect 262306 7352 262312 7404
rect 262364 7352 262370 7404
rect 263042 7352 263048 7404
rect 263100 7352 263106 7404
rect 264146 7352 264152 7404
rect 264204 7352 264210 7404
rect 264238 7352 264244 7404
rect 264296 7392 264302 7404
rect 265069 7395 265127 7401
rect 265069 7392 265081 7395
rect 264296 7364 265081 7392
rect 264296 7352 264302 7364
rect 265069 7361 265081 7364
rect 265115 7361 265127 7395
rect 265069 7355 265127 7361
rect 265250 7352 265256 7404
rect 265308 7392 265314 7404
rect 265713 7395 265771 7401
rect 265713 7392 265725 7395
rect 265308 7364 265725 7392
rect 265308 7352 265314 7364
rect 265713 7361 265725 7364
rect 265759 7392 265771 7395
rect 266541 7395 266599 7401
rect 266541 7392 266553 7395
rect 265759 7364 266553 7392
rect 265759 7361 265771 7364
rect 265713 7355 265771 7361
rect 266541 7361 266553 7364
rect 266587 7392 266599 7395
rect 267366 7392 267372 7404
rect 266587 7364 267372 7392
rect 266587 7361 266599 7364
rect 266541 7355 266599 7361
rect 267366 7352 267372 7364
rect 267424 7352 267430 7404
rect 267642 7352 267648 7404
rect 267700 7392 267706 7404
rect 268120 7392 268148 7432
rect 268749 7429 268761 7432
rect 268795 7460 268807 7463
rect 270034 7460 270040 7472
rect 268795 7432 270040 7460
rect 268795 7429 268807 7432
rect 268749 7423 268807 7429
rect 270034 7420 270040 7432
rect 270092 7420 270098 7472
rect 267700 7364 268148 7392
rect 267700 7352 267706 7364
rect 268378 7352 268384 7404
rect 268436 7352 268442 7404
rect 269482 7352 269488 7404
rect 269540 7352 269546 7404
rect 270129 7395 270187 7401
rect 270129 7361 270141 7395
rect 270175 7392 270187 7395
rect 270494 7392 270500 7404
rect 270175 7364 270500 7392
rect 270175 7361 270187 7364
rect 270129 7355 270187 7361
rect 270494 7352 270500 7364
rect 270552 7352 270558 7404
rect 265529 7327 265587 7333
rect 260484 7296 265480 7324
rect 263870 7256 263876 7268
rect 259840 7228 263876 7256
rect 263870 7216 263876 7228
rect 263928 7216 263934 7268
rect 265452 7256 265480 7296
rect 265529 7293 265541 7327
rect 265575 7324 265587 7327
rect 265802 7324 265808 7336
rect 265575 7296 265808 7324
rect 265575 7293 265587 7296
rect 265529 7287 265587 7293
rect 265802 7284 265808 7296
rect 265860 7284 265866 7336
rect 266357 7327 266415 7333
rect 266357 7293 266369 7327
rect 266403 7324 266415 7327
rect 266630 7324 266636 7336
rect 266403 7296 266636 7324
rect 266403 7293 266415 7296
rect 266357 7287 266415 7293
rect 266630 7284 266636 7296
rect 266688 7284 266694 7336
rect 266998 7284 267004 7336
rect 267056 7324 267062 7336
rect 267185 7327 267243 7333
rect 267185 7324 267197 7327
rect 267056 7296 267197 7324
rect 267056 7284 267062 7296
rect 267185 7293 267197 7296
rect 267231 7324 267243 7327
rect 267274 7324 267280 7336
rect 267231 7296 267280 7324
rect 267231 7293 267243 7296
rect 267185 7287 267243 7293
rect 267274 7284 267280 7296
rect 267332 7284 267338 7336
rect 268010 7324 268016 7336
rect 267660 7296 268016 7324
rect 267660 7256 267688 7296
rect 268010 7284 268016 7296
rect 268068 7284 268074 7336
rect 268194 7284 268200 7336
rect 268252 7324 268258 7336
rect 269301 7327 269359 7333
rect 269301 7324 269313 7327
rect 268252 7296 269313 7324
rect 268252 7284 268258 7296
rect 269301 7293 269313 7296
rect 269347 7293 269359 7327
rect 269301 7287 269359 7293
rect 270405 7327 270463 7333
rect 270405 7293 270417 7327
rect 270451 7293 270463 7327
rect 270405 7287 270463 7293
rect 265452 7228 267688 7256
rect 267734 7216 267740 7268
rect 267792 7256 267798 7268
rect 270420 7256 270448 7287
rect 271138 7284 271144 7336
rect 271196 7324 271202 7336
rect 271966 7324 271972 7336
rect 271196 7296 271972 7324
rect 271196 7284 271202 7296
rect 271966 7284 271972 7296
rect 272024 7284 272030 7336
rect 267792 7228 270448 7256
rect 267792 7216 267798 7228
rect 226978 7188 226984 7200
rect 222488 7160 226984 7188
rect 226978 7148 226984 7160
rect 227036 7148 227042 7200
rect 229557 7191 229615 7197
rect 229557 7157 229569 7191
rect 229603 7188 229615 7191
rect 230198 7188 230204 7200
rect 229603 7160 230204 7188
rect 229603 7157 229615 7160
rect 229557 7151 229615 7157
rect 230198 7148 230204 7160
rect 230256 7148 230262 7200
rect 230290 7148 230296 7200
rect 230348 7188 230354 7200
rect 230385 7191 230443 7197
rect 230385 7188 230397 7191
rect 230348 7160 230397 7188
rect 230348 7148 230354 7160
rect 230385 7157 230397 7160
rect 230431 7157 230443 7191
rect 230385 7151 230443 7157
rect 235626 7148 235632 7200
rect 235684 7148 235690 7200
rect 235994 7148 236000 7200
rect 236052 7188 236058 7200
rect 237282 7188 237288 7200
rect 236052 7160 237288 7188
rect 236052 7148 236058 7160
rect 237282 7148 237288 7160
rect 237340 7148 237346 7200
rect 237374 7148 237380 7200
rect 237432 7188 237438 7200
rect 237653 7191 237711 7197
rect 237653 7188 237665 7191
rect 237432 7160 237665 7188
rect 237432 7148 237438 7160
rect 237653 7157 237665 7160
rect 237699 7157 237711 7191
rect 237653 7151 237711 7157
rect 238754 7148 238760 7200
rect 238812 7148 238818 7200
rect 239122 7148 239128 7200
rect 239180 7148 239186 7200
rect 260929 7191 260987 7197
rect 260929 7157 260941 7191
rect 260975 7188 260987 7191
rect 262674 7188 262680 7200
rect 260975 7160 262680 7188
rect 260975 7157 260987 7160
rect 260929 7151 260987 7157
rect 262674 7148 262680 7160
rect 262732 7148 262738 7200
rect 264882 7148 264888 7200
rect 264940 7148 264946 7200
rect 266725 7191 266783 7197
rect 266725 7157 266737 7191
rect 266771 7188 266783 7191
rect 267458 7188 267464 7200
rect 266771 7160 267464 7188
rect 266771 7157 266783 7160
rect 266725 7151 266783 7157
rect 267458 7148 267464 7160
rect 267516 7148 267522 7200
rect 267553 7191 267611 7197
rect 267553 7157 267565 7191
rect 267599 7188 267611 7191
rect 267642 7188 267648 7200
rect 267599 7160 267648 7188
rect 267599 7157 267611 7160
rect 267553 7151 267611 7157
rect 267642 7148 267648 7160
rect 267700 7148 267706 7200
rect 269390 7148 269396 7200
rect 269448 7188 269454 7200
rect 269669 7191 269727 7197
rect 269669 7188 269681 7191
rect 269448 7160 269681 7188
rect 269448 7148 269454 7160
rect 269669 7157 269681 7160
rect 269715 7157 269727 7191
rect 269669 7151 269727 7157
rect 1104 7098 271492 7120
rect 1104 7046 34748 7098
rect 34800 7046 34812 7098
rect 34864 7046 34876 7098
rect 34928 7046 34940 7098
rect 34992 7046 35004 7098
rect 35056 7046 102345 7098
rect 102397 7046 102409 7098
rect 102461 7046 102473 7098
rect 102525 7046 102537 7098
rect 102589 7046 102601 7098
rect 102653 7046 169942 7098
rect 169994 7046 170006 7098
rect 170058 7046 170070 7098
rect 170122 7046 170134 7098
rect 170186 7046 170198 7098
rect 170250 7046 237539 7098
rect 237591 7046 237603 7098
rect 237655 7046 237667 7098
rect 237719 7046 237731 7098
rect 237783 7046 237795 7098
rect 237847 7046 271492 7098
rect 1104 7024 271492 7046
rect 79042 6944 79048 6996
rect 79100 6984 79106 6996
rect 79229 6987 79287 6993
rect 79229 6984 79241 6987
rect 79100 6956 79241 6984
rect 79100 6944 79106 6956
rect 79229 6953 79241 6956
rect 79275 6953 79287 6987
rect 79229 6947 79287 6953
rect 79410 6944 79416 6996
rect 79468 6944 79474 6996
rect 100938 6944 100944 6996
rect 100996 6984 101002 6996
rect 150250 6984 150256 6996
rect 100996 6956 150256 6984
rect 100996 6944 101002 6956
rect 150250 6944 150256 6956
rect 150308 6944 150314 6996
rect 165154 6944 165160 6996
rect 165212 6984 165218 6996
rect 169110 6984 169116 6996
rect 165212 6956 169116 6984
rect 165212 6944 165218 6956
rect 169110 6944 169116 6956
rect 169168 6944 169174 6996
rect 169573 6987 169631 6993
rect 169573 6953 169585 6987
rect 169619 6984 169631 6987
rect 169619 6956 171134 6984
rect 169619 6953 169631 6956
rect 169573 6947 169631 6953
rect 26970 6916 26976 6928
rect 19306 6888 26976 6916
rect 19306 6656 19334 6888
rect 26970 6876 26976 6888
rect 27028 6876 27034 6928
rect 99834 6876 99840 6928
rect 99892 6916 99898 6928
rect 100021 6919 100079 6925
rect 100021 6916 100033 6919
rect 99892 6888 100033 6916
rect 99892 6876 99898 6888
rect 100021 6885 100033 6888
rect 100067 6885 100079 6919
rect 100021 6879 100079 6885
rect 107102 6876 107108 6928
rect 107160 6916 107166 6928
rect 107746 6916 107752 6928
rect 107160 6888 107752 6916
rect 107160 6876 107166 6888
rect 107746 6876 107752 6888
rect 107804 6876 107810 6928
rect 108684 6888 108896 6916
rect 26142 6848 26148 6860
rect 22066 6820 26148 6848
rect 19978 6740 19984 6792
rect 20036 6780 20042 6792
rect 22066 6780 22094 6820
rect 26142 6808 26148 6820
rect 26200 6808 26206 6860
rect 75822 6808 75828 6860
rect 75880 6848 75886 6860
rect 79686 6848 79692 6860
rect 75880 6820 79692 6848
rect 75880 6808 75886 6820
rect 79686 6808 79692 6820
rect 79744 6808 79750 6860
rect 92842 6808 92848 6860
rect 92900 6848 92906 6860
rect 93213 6851 93271 6857
rect 93213 6848 93225 6851
rect 92900 6820 93225 6848
rect 92900 6808 92906 6820
rect 93213 6817 93225 6820
rect 93259 6817 93271 6851
rect 93213 6811 93271 6817
rect 99006 6808 99012 6860
rect 99064 6848 99070 6860
rect 99561 6851 99619 6857
rect 99561 6848 99573 6851
rect 99064 6820 99573 6848
rect 99064 6808 99070 6820
rect 99561 6817 99573 6820
rect 99607 6817 99619 6851
rect 99561 6811 99619 6817
rect 100294 6808 100300 6860
rect 100352 6808 100358 6860
rect 100435 6851 100493 6857
rect 100435 6817 100447 6851
rect 100481 6848 100493 6851
rect 104434 6848 104440 6860
rect 100481 6820 104440 6848
rect 100481 6817 100493 6820
rect 100435 6811 100493 6817
rect 104434 6808 104440 6820
rect 104492 6808 104498 6860
rect 108301 6851 108359 6857
rect 108301 6848 108313 6851
rect 107764 6820 108313 6848
rect 20036 6752 22094 6780
rect 20036 6740 20042 6752
rect 24210 6740 24216 6792
rect 24268 6780 24274 6792
rect 25593 6783 25651 6789
rect 25593 6780 25605 6783
rect 24268 6752 25605 6780
rect 24268 6740 24274 6752
rect 25593 6749 25605 6752
rect 25639 6749 25651 6783
rect 25593 6743 25651 6749
rect 26510 6740 26516 6792
rect 26568 6740 26574 6792
rect 33042 6740 33048 6792
rect 33100 6780 33106 6792
rect 43990 6780 43996 6792
rect 33100 6752 43996 6780
rect 33100 6740 33106 6752
rect 43990 6740 43996 6752
rect 44048 6740 44054 6792
rect 47854 6740 47860 6792
rect 47912 6780 47918 6792
rect 87874 6780 87880 6792
rect 47912 6752 87880 6780
rect 47912 6740 47918 6752
rect 87874 6740 87880 6752
rect 87932 6740 87938 6792
rect 92474 6740 92480 6792
rect 92532 6780 92538 6792
rect 92753 6783 92811 6789
rect 92753 6780 92765 6783
rect 92532 6752 92765 6780
rect 92532 6740 92538 6752
rect 92753 6749 92765 6752
rect 92799 6749 92811 6783
rect 98641 6783 98699 6789
rect 98641 6780 98653 6783
rect 92753 6743 92811 6749
rect 93596 6752 98653 6780
rect 24394 6672 24400 6724
rect 24452 6712 24458 6724
rect 38562 6712 38568 6724
rect 24452 6684 38568 6712
rect 24452 6672 24458 6684
rect 38562 6672 38568 6684
rect 38620 6672 38626 6724
rect 42610 6672 42616 6724
rect 42668 6712 42674 6724
rect 49878 6712 49884 6724
rect 42668 6684 49884 6712
rect 42668 6672 42674 6684
rect 49878 6672 49884 6684
rect 49936 6672 49942 6724
rect 79045 6715 79103 6721
rect 79045 6681 79057 6715
rect 79091 6712 79103 6715
rect 79134 6712 79140 6724
rect 79091 6684 79140 6712
rect 79091 6681 79103 6684
rect 79045 6675 79103 6681
rect 79134 6672 79140 6684
rect 79192 6672 79198 6724
rect 89622 6672 89628 6724
rect 89680 6712 89686 6724
rect 93596 6712 93624 6752
rect 98641 6749 98653 6752
rect 98687 6780 98699 6783
rect 99377 6783 99435 6789
rect 99377 6780 99389 6783
rect 98687 6752 99389 6780
rect 98687 6749 98699 6752
rect 98641 6743 98699 6749
rect 99377 6749 99389 6752
rect 99423 6749 99435 6783
rect 99377 6743 99435 6749
rect 100570 6740 100576 6792
rect 100628 6740 100634 6792
rect 101306 6740 101312 6792
rect 101364 6780 101370 6792
rect 107764 6789 107792 6820
rect 108301 6817 108313 6820
rect 108347 6817 108359 6851
rect 108684 6848 108712 6888
rect 108301 6811 108359 6817
rect 108408 6820 108712 6848
rect 102229 6783 102287 6789
rect 102229 6780 102241 6783
rect 101364 6752 102241 6780
rect 101364 6740 101370 6752
rect 102229 6749 102241 6752
rect 102275 6749 102287 6783
rect 107749 6783 107807 6789
rect 107749 6780 107761 6783
rect 102229 6743 102287 6749
rect 102704 6752 107761 6780
rect 102704 6712 102732 6752
rect 107749 6749 107761 6752
rect 107795 6749 107807 6783
rect 107749 6743 107807 6749
rect 108114 6740 108120 6792
rect 108172 6780 108178 6792
rect 108408 6780 108436 6820
rect 108758 6808 108764 6860
rect 108816 6808 108822 6860
rect 108868 6848 108896 6888
rect 146294 6876 146300 6928
rect 146352 6916 146358 6928
rect 146352 6888 146524 6916
rect 146352 6876 146358 6888
rect 110233 6851 110291 6857
rect 110233 6848 110245 6851
rect 108868 6820 110245 6848
rect 110233 6817 110245 6820
rect 110279 6817 110291 6851
rect 110233 6811 110291 6817
rect 112438 6808 112444 6860
rect 112496 6808 112502 6860
rect 113174 6808 113180 6860
rect 113232 6848 113238 6860
rect 114557 6851 114615 6857
rect 114557 6848 114569 6851
rect 113232 6820 114569 6848
rect 113232 6808 113238 6820
rect 114557 6817 114569 6820
rect 114603 6848 114615 6851
rect 114922 6848 114928 6860
rect 114603 6820 114928 6848
rect 114603 6817 114615 6820
rect 114557 6811 114615 6817
rect 114922 6808 114928 6820
rect 114980 6808 114986 6860
rect 140498 6808 140504 6860
rect 140556 6848 140562 6860
rect 140685 6851 140743 6857
rect 140685 6848 140697 6851
rect 140556 6820 140697 6848
rect 140556 6808 140562 6820
rect 140685 6817 140697 6820
rect 140731 6817 140743 6851
rect 140685 6811 140743 6817
rect 141326 6808 141332 6860
rect 141384 6808 141390 6860
rect 141602 6808 141608 6860
rect 141660 6808 141666 6860
rect 141694 6808 141700 6860
rect 141752 6857 141758 6860
rect 141752 6851 141780 6857
rect 141768 6817 141780 6851
rect 141752 6811 141780 6817
rect 141752 6808 141758 6811
rect 145834 6808 145840 6860
rect 145892 6808 145898 6860
rect 146021 6851 146079 6857
rect 146021 6817 146033 6851
rect 146067 6848 146079 6851
rect 146386 6848 146392 6860
rect 146067 6820 146392 6848
rect 146067 6817 146079 6820
rect 146021 6811 146079 6817
rect 146386 6808 146392 6820
rect 146444 6808 146450 6860
rect 146496 6857 146524 6888
rect 159174 6876 159180 6928
rect 159232 6916 159238 6928
rect 161842 6916 161848 6928
rect 159232 6888 161848 6916
rect 159232 6876 159238 6888
rect 161842 6876 161848 6888
rect 161900 6876 161906 6928
rect 169754 6876 169760 6928
rect 169812 6876 169818 6928
rect 171106 6916 171134 6956
rect 180058 6944 180064 6996
rect 180116 6984 180122 6996
rect 180116 6956 214420 6984
rect 180116 6944 180122 6956
rect 180978 6916 180984 6928
rect 171106 6888 180984 6916
rect 180978 6876 180984 6888
rect 181036 6876 181042 6928
rect 189994 6876 190000 6928
rect 190052 6876 190058 6928
rect 146481 6851 146539 6857
rect 146481 6817 146493 6851
rect 146527 6848 146539 6851
rect 147582 6848 147588 6860
rect 146527 6820 147588 6848
rect 146527 6817 146539 6820
rect 146481 6811 146539 6817
rect 147582 6808 147588 6820
rect 147640 6808 147646 6860
rect 148226 6808 148232 6860
rect 148284 6808 148290 6860
rect 148873 6851 148931 6857
rect 148873 6817 148885 6851
rect 148919 6848 148931 6851
rect 148962 6848 148968 6860
rect 148919 6820 148968 6848
rect 148919 6817 148931 6820
rect 148873 6811 148931 6817
rect 148962 6808 148968 6820
rect 149020 6808 149026 6860
rect 149146 6808 149152 6860
rect 149204 6808 149210 6860
rect 149287 6851 149345 6857
rect 149287 6817 149299 6851
rect 149333 6848 149345 6851
rect 150342 6848 150348 6860
rect 149333 6820 150348 6848
rect 149333 6817 149345 6820
rect 149287 6811 149345 6817
rect 150342 6808 150348 6820
rect 150400 6808 150406 6860
rect 150526 6808 150532 6860
rect 150584 6808 150590 6860
rect 150894 6808 150900 6860
rect 150952 6848 150958 6860
rect 151173 6851 151231 6857
rect 151173 6848 151185 6851
rect 150952 6820 151185 6848
rect 150952 6808 150958 6820
rect 151173 6817 151185 6820
rect 151219 6817 151231 6851
rect 151173 6811 151231 6817
rect 151446 6808 151452 6860
rect 151504 6808 151510 6860
rect 152366 6808 152372 6860
rect 152424 6808 152430 6860
rect 189074 6848 189080 6860
rect 169220 6820 189080 6848
rect 169220 6792 169248 6820
rect 189074 6808 189080 6820
rect 189132 6808 189138 6860
rect 208762 6808 208768 6860
rect 208820 6848 208826 6860
rect 210237 6851 210295 6857
rect 210237 6848 210249 6851
rect 208820 6820 210249 6848
rect 208820 6808 208826 6820
rect 210237 6817 210249 6820
rect 210283 6817 210295 6851
rect 210237 6811 210295 6817
rect 210786 6808 210792 6860
rect 210844 6848 210850 6860
rect 210881 6851 210939 6857
rect 210881 6848 210893 6851
rect 210844 6820 210893 6848
rect 210844 6808 210850 6820
rect 210881 6817 210893 6820
rect 210927 6817 210939 6851
rect 210881 6811 210939 6817
rect 212537 6851 212595 6857
rect 212537 6817 212549 6851
rect 212583 6848 212595 6851
rect 213914 6848 213920 6860
rect 212583 6820 213920 6848
rect 212583 6817 212595 6820
rect 212537 6811 212595 6817
rect 213914 6808 213920 6820
rect 213972 6808 213978 6860
rect 214392 6857 214420 6956
rect 215110 6944 215116 6996
rect 215168 6944 215174 6996
rect 215478 6944 215484 6996
rect 215536 6984 215542 6996
rect 215536 6956 220768 6984
rect 215536 6944 215542 6956
rect 215128 6916 215156 6944
rect 215938 6916 215944 6928
rect 215128 6888 215944 6916
rect 215938 6876 215944 6888
rect 215996 6916 216002 6928
rect 216582 6916 216588 6928
rect 215996 6888 216588 6916
rect 215996 6876 216002 6888
rect 216582 6876 216588 6888
rect 216640 6916 216646 6928
rect 216640 6888 218192 6916
rect 216640 6876 216646 6888
rect 214377 6851 214435 6857
rect 214377 6848 214389 6851
rect 214335 6820 214389 6848
rect 214377 6817 214389 6820
rect 214423 6848 214435 6851
rect 215110 6848 215116 6860
rect 214423 6820 215116 6848
rect 214423 6817 214435 6820
rect 214377 6811 214435 6817
rect 215110 6808 215116 6820
rect 215168 6808 215174 6860
rect 215665 6851 215723 6857
rect 215665 6817 215677 6851
rect 215711 6848 215723 6851
rect 218054 6848 218060 6860
rect 215711 6820 218060 6848
rect 215711 6817 215723 6820
rect 215665 6811 215723 6817
rect 218054 6808 218060 6820
rect 218112 6808 218118 6860
rect 218164 6848 218192 6888
rect 218330 6876 218336 6928
rect 218388 6916 218394 6928
rect 220740 6916 220768 6956
rect 220814 6944 220820 6996
rect 220872 6984 220878 6996
rect 225230 6984 225236 6996
rect 220872 6956 225236 6984
rect 220872 6944 220878 6956
rect 225230 6944 225236 6956
rect 225288 6944 225294 6996
rect 226242 6944 226248 6996
rect 226300 6984 226306 6996
rect 229186 6984 229192 6996
rect 226300 6956 229192 6984
rect 226300 6944 226306 6956
rect 229186 6944 229192 6956
rect 229244 6944 229250 6996
rect 229925 6987 229983 6993
rect 229925 6953 229937 6987
rect 229971 6953 229983 6987
rect 229925 6947 229983 6953
rect 220906 6916 220912 6928
rect 218388 6888 218744 6916
rect 220740 6888 220912 6916
rect 218388 6876 218394 6888
rect 218609 6851 218667 6857
rect 218609 6848 218621 6851
rect 218164 6820 218621 6848
rect 218609 6817 218621 6820
rect 218655 6817 218667 6851
rect 218716 6848 218744 6888
rect 220906 6876 220912 6888
rect 220964 6876 220970 6928
rect 223224 6888 223436 6916
rect 219161 6851 219219 6857
rect 219161 6848 219173 6851
rect 218716 6820 219173 6848
rect 218609 6811 218667 6817
rect 219161 6817 219173 6820
rect 219207 6817 219219 6851
rect 219161 6811 219219 6817
rect 219342 6808 219348 6860
rect 219400 6848 219406 6860
rect 220173 6851 220231 6857
rect 220173 6848 220185 6851
rect 219400 6820 220185 6848
rect 219400 6808 219406 6820
rect 220173 6817 220185 6820
rect 220219 6817 220231 6851
rect 220538 6848 220544 6860
rect 220173 6811 220231 6817
rect 220280 6820 220544 6848
rect 108172 6752 108436 6780
rect 108172 6740 108178 6752
rect 109034 6740 109040 6792
rect 109092 6740 109098 6792
rect 109218 6789 109224 6792
rect 109175 6783 109224 6789
rect 109175 6749 109187 6783
rect 109221 6749 109224 6783
rect 109175 6743 109224 6749
rect 109218 6740 109224 6743
rect 109276 6740 109282 6792
rect 109310 6740 109316 6792
rect 109368 6740 109374 6792
rect 140866 6740 140872 6792
rect 140924 6740 140930 6792
rect 141878 6740 141884 6792
rect 141936 6740 141942 6792
rect 146754 6740 146760 6792
rect 146812 6740 146818 6792
rect 146938 6789 146944 6792
rect 146895 6783 146944 6789
rect 146895 6749 146907 6783
rect 146941 6749 146944 6783
rect 146895 6743 146944 6749
rect 146938 6740 146944 6743
rect 146996 6740 147002 6792
rect 147030 6740 147036 6792
rect 147088 6740 147094 6792
rect 148318 6740 148324 6792
rect 148376 6780 148382 6792
rect 148413 6783 148471 6789
rect 148413 6780 148425 6783
rect 148376 6752 148425 6780
rect 148376 6740 148382 6752
rect 148413 6749 148425 6752
rect 148459 6749 148471 6783
rect 148413 6743 148471 6749
rect 149422 6740 149428 6792
rect 149480 6740 149486 6792
rect 150618 6740 150624 6792
rect 150676 6780 150682 6792
rect 150713 6783 150771 6789
rect 150713 6780 150725 6783
rect 150676 6752 150725 6780
rect 150676 6740 150682 6752
rect 150713 6749 150725 6752
rect 150759 6749 150771 6783
rect 150713 6743 150771 6749
rect 151538 6740 151544 6792
rect 151596 6789 151602 6792
rect 151596 6783 151624 6789
rect 151612 6749 151624 6783
rect 151596 6743 151624 6749
rect 151596 6740 151602 6743
rect 151722 6740 151728 6792
rect 151780 6740 151786 6792
rect 169202 6740 169208 6792
rect 169260 6740 169266 6792
rect 170309 6783 170367 6789
rect 170309 6749 170321 6783
rect 170355 6780 170367 6783
rect 172514 6780 172520 6792
rect 170355 6752 172520 6780
rect 170355 6749 170367 6752
rect 170309 6743 170367 6749
rect 172514 6740 172520 6752
rect 172572 6740 172578 6792
rect 189350 6740 189356 6792
rect 189408 6780 189414 6792
rect 190181 6783 190239 6789
rect 190181 6780 190193 6783
rect 189408 6752 190193 6780
rect 189408 6740 189414 6752
rect 190181 6749 190193 6752
rect 190227 6749 190239 6783
rect 190181 6743 190239 6749
rect 209866 6740 209872 6792
rect 209924 6780 209930 6792
rect 210421 6783 210479 6789
rect 210421 6780 210433 6783
rect 209924 6752 210433 6780
rect 209924 6740 209930 6752
rect 210421 6749 210433 6752
rect 210467 6749 210479 6783
rect 210421 6743 210479 6749
rect 211154 6740 211160 6792
rect 211212 6740 211218 6792
rect 211338 6789 211344 6792
rect 211295 6783 211344 6789
rect 211295 6749 211307 6783
rect 211341 6749 211344 6783
rect 211295 6743 211344 6749
rect 211338 6740 211344 6743
rect 211396 6740 211402 6792
rect 211430 6740 211436 6792
rect 211488 6740 211494 6792
rect 213932 6752 215294 6780
rect 89680 6684 93624 6712
rect 94332 6684 99374 6712
rect 89680 6672 89686 6684
rect 19242 6604 19248 6656
rect 19300 6616 19334 6656
rect 19300 6604 19306 6616
rect 24762 6604 24768 6656
rect 24820 6644 24826 6656
rect 25777 6647 25835 6653
rect 25777 6644 25789 6647
rect 24820 6616 25789 6644
rect 24820 6604 24826 6616
rect 25777 6613 25789 6616
rect 25823 6613 25835 6647
rect 25777 6607 25835 6613
rect 26694 6604 26700 6656
rect 26752 6604 26758 6656
rect 43898 6604 43904 6656
rect 43956 6644 43962 6656
rect 44453 6647 44511 6653
rect 44453 6644 44465 6647
rect 43956 6616 44465 6644
rect 43956 6604 43962 6616
rect 44453 6613 44465 6616
rect 44499 6613 44511 6647
rect 44453 6607 44511 6613
rect 79255 6647 79313 6653
rect 79255 6613 79267 6647
rect 79301 6644 79313 6647
rect 79410 6644 79416 6656
rect 79301 6616 79416 6644
rect 79301 6613 79313 6616
rect 79255 6607 79313 6613
rect 79410 6604 79416 6616
rect 79468 6604 79474 6656
rect 80054 6604 80060 6656
rect 80112 6644 80118 6656
rect 94332 6644 94360 6684
rect 80112 6616 94360 6644
rect 80112 6604 80118 6616
rect 99006 6604 99012 6656
rect 99064 6604 99070 6656
rect 99346 6644 99374 6684
rect 101140 6684 102732 6712
rect 101140 6644 101168 6684
rect 102778 6672 102784 6724
rect 102836 6672 102842 6724
rect 103330 6672 103336 6724
rect 103388 6712 103394 6724
rect 106734 6712 106740 6724
rect 103388 6684 106740 6712
rect 103388 6672 103394 6684
rect 106734 6672 106740 6684
rect 106792 6672 106798 6724
rect 109788 6684 110092 6712
rect 99346 6616 101168 6644
rect 101217 6647 101275 6653
rect 101217 6613 101229 6647
rect 101263 6644 101275 6647
rect 101766 6644 101772 6656
rect 101263 6616 101772 6644
rect 101263 6613 101275 6616
rect 101217 6607 101275 6613
rect 101766 6604 101772 6616
rect 101824 6604 101830 6656
rect 109034 6604 109040 6656
rect 109092 6644 109098 6656
rect 109788 6644 109816 6684
rect 109092 6616 109816 6644
rect 109092 6604 109098 6616
rect 109954 6604 109960 6656
rect 110012 6604 110018 6656
rect 110064 6644 110092 6684
rect 112622 6672 112628 6724
rect 112680 6672 112686 6724
rect 114370 6672 114376 6724
rect 114428 6712 114434 6724
rect 125594 6712 125600 6724
rect 114428 6684 125600 6712
rect 114428 6672 114434 6684
rect 125594 6672 125600 6684
rect 125652 6672 125658 6724
rect 147508 6684 148456 6712
rect 113358 6644 113364 6656
rect 110064 6616 113364 6644
rect 113358 6604 113364 6616
rect 113416 6604 113422 6656
rect 115750 6604 115756 6656
rect 115808 6644 115814 6656
rect 123478 6644 123484 6656
rect 115808 6616 123484 6644
rect 115808 6604 115814 6616
rect 123478 6604 123484 6616
rect 123536 6604 123542 6656
rect 140409 6647 140467 6653
rect 140409 6613 140421 6647
rect 140455 6644 140467 6647
rect 141694 6644 141700 6656
rect 140455 6616 141700 6644
rect 140455 6613 140467 6616
rect 140409 6607 140467 6613
rect 141694 6604 141700 6616
rect 141752 6604 141758 6656
rect 142525 6647 142583 6653
rect 142525 6613 142537 6647
rect 142571 6644 142583 6647
rect 143074 6644 143080 6656
rect 142571 6616 143080 6644
rect 142571 6613 142583 6616
rect 142525 6607 142583 6613
rect 143074 6604 143080 6616
rect 143132 6604 143138 6656
rect 146846 6604 146852 6656
rect 146904 6644 146910 6656
rect 147030 6644 147036 6656
rect 146904 6616 147036 6644
rect 146904 6604 146910 6616
rect 147030 6604 147036 6616
rect 147088 6644 147094 6656
rect 147508 6644 147536 6684
rect 147088 6616 147536 6644
rect 147677 6647 147735 6653
rect 147088 6604 147094 6616
rect 147677 6613 147689 6647
rect 147723 6644 147735 6647
rect 148226 6644 148232 6656
rect 147723 6616 148232 6644
rect 147723 6613 147735 6616
rect 147677 6607 147735 6613
rect 148226 6604 148232 6616
rect 148284 6604 148290 6656
rect 148428 6644 148456 6684
rect 149992 6684 150756 6712
rect 149422 6644 149428 6656
rect 148428 6616 149428 6644
rect 149422 6604 149428 6616
rect 149480 6644 149486 6656
rect 149992 6644 150020 6684
rect 149480 6616 150020 6644
rect 149480 6604 149486 6616
rect 150066 6604 150072 6656
rect 150124 6604 150130 6656
rect 150728 6644 150756 6684
rect 155586 6672 155592 6724
rect 155644 6712 155650 6724
rect 163498 6712 163504 6724
rect 155644 6684 163504 6712
rect 155644 6672 155650 6684
rect 163498 6672 163504 6684
rect 163556 6672 163562 6724
rect 212721 6715 212779 6721
rect 212000 6684 212212 6712
rect 151078 6644 151084 6656
rect 150728 6616 151084 6644
rect 151078 6604 151084 6616
rect 151136 6644 151142 6656
rect 151722 6644 151728 6656
rect 151136 6616 151728 6644
rect 151136 6604 151142 6616
rect 151722 6604 151728 6616
rect 151780 6604 151786 6656
rect 152366 6604 152372 6656
rect 152424 6644 152430 6656
rect 161106 6644 161112 6656
rect 152424 6616 161112 6644
rect 152424 6604 152430 6616
rect 161106 6604 161112 6616
rect 161164 6604 161170 6656
rect 162670 6604 162676 6656
rect 162728 6644 162734 6656
rect 169573 6647 169631 6653
rect 169573 6644 169585 6647
rect 162728 6616 169585 6644
rect 162728 6604 162734 6616
rect 169573 6613 169585 6616
rect 169619 6644 169631 6647
rect 170401 6647 170459 6653
rect 170401 6644 170413 6647
rect 169619 6616 170413 6644
rect 169619 6613 169631 6616
rect 169573 6607 169631 6613
rect 170401 6613 170413 6616
rect 170447 6613 170459 6647
rect 170401 6607 170459 6613
rect 198826 6604 198832 6656
rect 198884 6644 198890 6656
rect 212000 6644 212028 6684
rect 198884 6616 212028 6644
rect 198884 6604 198890 6616
rect 212074 6604 212080 6656
rect 212132 6604 212138 6656
rect 212184 6644 212212 6684
rect 212721 6681 212733 6715
rect 212767 6712 212779 6715
rect 212994 6712 213000 6724
rect 212767 6684 213000 6712
rect 212767 6681 212779 6684
rect 212721 6675 212779 6681
rect 212994 6672 213000 6684
rect 213052 6712 213058 6724
rect 213932 6712 213960 6752
rect 213052 6684 213960 6712
rect 215266 6712 215294 6752
rect 217686 6740 217692 6792
rect 217744 6780 217750 6792
rect 217965 6783 218023 6789
rect 217965 6780 217977 6783
rect 217744 6752 217977 6780
rect 217744 6740 217750 6752
rect 217965 6749 217977 6752
rect 218011 6749 218023 6783
rect 217965 6743 218023 6749
rect 218149 6783 218207 6789
rect 218149 6749 218161 6783
rect 218195 6749 218207 6783
rect 218149 6743 218207 6749
rect 215849 6715 215907 6721
rect 215849 6712 215861 6715
rect 215266 6684 215861 6712
rect 213052 6672 213058 6684
rect 215849 6681 215861 6684
rect 215895 6712 215907 6715
rect 216306 6712 216312 6724
rect 215895 6684 216312 6712
rect 215895 6681 215907 6684
rect 215849 6675 215907 6681
rect 216306 6672 216312 6684
rect 216364 6672 216370 6724
rect 217505 6715 217563 6721
rect 217505 6681 217517 6715
rect 217551 6681 217563 6715
rect 217505 6675 217563 6681
rect 214282 6644 214288 6656
rect 212184 6616 214288 6644
rect 214282 6604 214288 6616
rect 214340 6604 214346 6656
rect 215389 6647 215447 6653
rect 215389 6613 215401 6647
rect 215435 6644 215447 6647
rect 215570 6644 215576 6656
rect 215435 6616 215576 6644
rect 215435 6613 215447 6616
rect 215389 6607 215447 6613
rect 215570 6604 215576 6616
rect 215628 6644 215634 6656
rect 217520 6644 217548 6675
rect 217594 6672 217600 6724
rect 217652 6712 217658 6724
rect 218164 6712 218192 6743
rect 218882 6740 218888 6792
rect 218940 6740 218946 6792
rect 219066 6789 219072 6792
rect 219023 6783 219072 6789
rect 219023 6749 219035 6783
rect 219069 6749 219072 6783
rect 219023 6743 219072 6749
rect 219066 6740 219072 6743
rect 219124 6740 219130 6792
rect 219894 6740 219900 6792
rect 219952 6780 219958 6792
rect 220280 6780 220308 6820
rect 220538 6808 220544 6820
rect 220596 6848 220602 6860
rect 220817 6851 220875 6857
rect 220817 6848 220829 6851
rect 220596 6820 220829 6848
rect 220596 6808 220602 6820
rect 220817 6817 220829 6820
rect 220863 6817 220875 6851
rect 220817 6811 220875 6817
rect 221090 6808 221096 6860
rect 221148 6808 221154 6860
rect 221379 6851 221437 6857
rect 221379 6817 221391 6851
rect 221425 6848 221437 6851
rect 221734 6848 221740 6860
rect 221425 6820 221740 6848
rect 221425 6817 221437 6820
rect 221379 6811 221437 6817
rect 221734 6808 221740 6820
rect 221792 6808 221798 6860
rect 221918 6808 221924 6860
rect 221976 6808 221982 6860
rect 222102 6808 222108 6860
rect 222160 6848 222166 6860
rect 222657 6851 222715 6857
rect 222657 6848 222669 6851
rect 222160 6820 222669 6848
rect 222160 6808 222166 6820
rect 222657 6817 222669 6820
rect 222703 6817 222715 6851
rect 223224 6848 223252 6888
rect 222657 6811 222715 6817
rect 222764 6820 223252 6848
rect 221274 6789 221280 6792
rect 219952 6752 220308 6780
rect 220357 6783 220415 6789
rect 219952 6740 219958 6752
rect 220357 6749 220369 6783
rect 220403 6749 220415 6783
rect 220357 6743 220415 6749
rect 221231 6783 221280 6789
rect 221231 6749 221243 6783
rect 221277 6749 221280 6783
rect 221231 6743 221280 6749
rect 217652 6684 218192 6712
rect 217652 6672 217658 6684
rect 217686 6644 217692 6656
rect 215628 6616 217692 6644
rect 215628 6604 215634 6616
rect 217686 6604 217692 6616
rect 217744 6644 217750 6656
rect 217781 6647 217839 6653
rect 217781 6644 217793 6647
rect 217744 6616 217793 6644
rect 217744 6604 217750 6616
rect 217781 6613 217793 6616
rect 217827 6613 217839 6647
rect 217781 6607 217839 6613
rect 217870 6604 217876 6656
rect 217928 6644 217934 6656
rect 219805 6647 219863 6653
rect 219805 6644 219817 6647
rect 217928 6616 219817 6644
rect 217928 6604 217934 6616
rect 219805 6613 219817 6616
rect 219851 6613 219863 6647
rect 220372 6644 220400 6743
rect 221274 6740 221280 6743
rect 221332 6740 221338 6792
rect 221936 6780 221964 6808
rect 222286 6780 222292 6792
rect 221936 6752 222292 6780
rect 222286 6740 222292 6752
rect 222344 6740 222350 6792
rect 222381 6783 222439 6789
rect 222381 6749 222393 6783
rect 222427 6780 222439 6783
rect 222764 6780 222792 6820
rect 223298 6808 223304 6860
rect 223356 6808 223362 6860
rect 223408 6848 223436 6888
rect 224954 6876 224960 6928
rect 225012 6916 225018 6928
rect 226334 6916 226340 6928
rect 225012 6888 226340 6916
rect 225012 6876 225018 6888
rect 226334 6876 226340 6888
rect 226392 6876 226398 6928
rect 229940 6916 229968 6947
rect 230106 6944 230112 6996
rect 230164 6944 230170 6996
rect 230474 6944 230480 6996
rect 230532 6984 230538 6996
rect 236914 6984 236920 6996
rect 230532 6956 236920 6984
rect 230532 6944 230538 6956
rect 236914 6944 236920 6956
rect 236972 6944 236978 6996
rect 244246 6956 265020 6984
rect 230842 6916 230848 6928
rect 229940 6888 230848 6916
rect 230842 6876 230848 6888
rect 230900 6876 230906 6928
rect 235718 6876 235724 6928
rect 235776 6916 235782 6928
rect 236546 6916 236552 6928
rect 235776 6888 236552 6916
rect 235776 6876 235782 6888
rect 236546 6876 236552 6888
rect 236604 6916 236610 6928
rect 244246 6916 244274 6956
rect 236604 6888 244274 6916
rect 236604 6876 236610 6888
rect 262674 6876 262680 6928
rect 262732 6876 262738 6928
rect 263686 6916 263692 6928
rect 262784 6888 263692 6916
rect 223577 6851 223635 6857
rect 223577 6848 223589 6851
rect 223408 6820 223589 6848
rect 223577 6817 223589 6820
rect 223623 6848 223635 6851
rect 224862 6848 224868 6860
rect 223623 6820 224868 6848
rect 223623 6817 223635 6820
rect 223577 6811 223635 6817
rect 224862 6808 224868 6820
rect 224920 6808 224926 6860
rect 225506 6808 225512 6860
rect 225564 6808 225570 6860
rect 229554 6808 229560 6860
rect 229612 6808 229618 6860
rect 235997 6851 236055 6857
rect 235997 6848 236009 6851
rect 229664 6820 236009 6848
rect 223758 6789 223764 6792
rect 222427 6752 222792 6780
rect 222841 6783 222899 6789
rect 222427 6749 222439 6752
rect 222381 6743 222439 6749
rect 222841 6749 222853 6783
rect 222887 6749 222899 6783
rect 222841 6743 222899 6749
rect 223715 6783 223764 6789
rect 223715 6749 223727 6783
rect 223761 6749 223764 6783
rect 223715 6743 223764 6749
rect 222102 6672 222108 6724
rect 222160 6712 222166 6724
rect 222856 6712 222884 6743
rect 223758 6740 223764 6743
rect 223816 6740 223822 6792
rect 223850 6740 223856 6792
rect 223908 6740 223914 6792
rect 224696 6752 225460 6780
rect 222160 6684 222884 6712
rect 222160 6672 222166 6684
rect 220906 6644 220912 6656
rect 220372 6616 220912 6644
rect 219805 6607 219863 6613
rect 220906 6604 220912 6616
rect 220964 6604 220970 6656
rect 222010 6604 222016 6656
rect 222068 6604 222074 6656
rect 223666 6604 223672 6656
rect 223724 6644 223730 6656
rect 224497 6647 224555 6653
rect 224497 6644 224509 6647
rect 223724 6616 224509 6644
rect 223724 6604 223730 6616
rect 224497 6613 224509 6616
rect 224543 6613 224555 6647
rect 224497 6607 224555 6613
rect 224586 6604 224592 6656
rect 224644 6644 224650 6656
rect 224696 6644 224724 6752
rect 224957 6647 225015 6653
rect 224957 6644 224969 6647
rect 224644 6616 224969 6644
rect 224644 6604 224650 6616
rect 224957 6613 224969 6616
rect 225003 6613 225015 6647
rect 225432 6644 225460 6752
rect 227622 6740 227628 6792
rect 227680 6780 227686 6792
rect 229664 6780 229692 6820
rect 235997 6817 236009 6820
rect 236043 6817 236055 6851
rect 237374 6848 237380 6860
rect 235997 6811 236055 6817
rect 236472 6820 237380 6848
rect 227680 6752 229692 6780
rect 227680 6740 227686 6752
rect 230474 6740 230480 6792
rect 230532 6740 230538 6792
rect 231118 6740 231124 6792
rect 231176 6740 231182 6792
rect 235721 6783 235779 6789
rect 235721 6749 235733 6783
rect 235767 6780 235779 6783
rect 236472 6780 236500 6820
rect 237374 6808 237380 6820
rect 237432 6808 237438 6860
rect 262784 6848 262812 6888
rect 263686 6876 263692 6888
rect 263744 6876 263750 6928
rect 264992 6916 265020 6956
rect 265066 6944 265072 6996
rect 265124 6984 265130 6996
rect 270954 6984 270960 6996
rect 265124 6956 270960 6984
rect 265124 6944 265130 6956
rect 270954 6944 270960 6956
rect 271012 6944 271018 6996
rect 266170 6916 266176 6928
rect 264992 6888 266176 6916
rect 266170 6876 266176 6888
rect 266228 6876 266234 6928
rect 268010 6848 268016 6860
rect 244246 6820 262812 6848
rect 262876 6820 268016 6848
rect 235767 6752 236500 6780
rect 236733 6783 236791 6789
rect 235767 6749 235779 6752
rect 235721 6743 235779 6749
rect 236733 6749 236745 6783
rect 236779 6780 236791 6783
rect 237101 6783 237159 6789
rect 237101 6780 237113 6783
rect 236779 6752 237113 6780
rect 236779 6749 236791 6752
rect 236733 6743 236791 6749
rect 237101 6749 237113 6752
rect 237147 6749 237159 6783
rect 237101 6743 237159 6749
rect 225693 6715 225751 6721
rect 225693 6681 225705 6715
rect 225739 6712 225751 6715
rect 225966 6712 225972 6724
rect 225739 6684 225972 6712
rect 225739 6681 225751 6684
rect 225693 6675 225751 6681
rect 225966 6672 225972 6684
rect 226024 6672 226030 6724
rect 227349 6715 227407 6721
rect 227349 6681 227361 6715
rect 227395 6712 227407 6715
rect 227395 6684 227760 6712
rect 227395 6681 227407 6684
rect 227349 6675 227407 6681
rect 227364 6644 227392 6675
rect 227732 6653 227760 6684
rect 229002 6672 229008 6724
rect 229060 6712 229066 6724
rect 230492 6712 230520 6740
rect 229060 6684 230520 6712
rect 229060 6672 229066 6684
rect 231762 6672 231768 6724
rect 231820 6672 231826 6724
rect 237116 6712 237144 6743
rect 237190 6740 237196 6792
rect 237248 6740 237254 6792
rect 244246 6780 244274 6820
rect 237300 6752 244274 6780
rect 237300 6712 237328 6752
rect 261018 6740 261024 6792
rect 261076 6740 261082 6792
rect 262217 6783 262275 6789
rect 262217 6749 262229 6783
rect 262263 6780 262275 6783
rect 262490 6780 262496 6792
rect 262263 6752 262496 6780
rect 262263 6749 262275 6752
rect 262217 6743 262275 6749
rect 262490 6740 262496 6752
rect 262548 6740 262554 6792
rect 262876 6789 262904 6820
rect 268010 6808 268016 6820
rect 268068 6808 268074 6860
rect 270865 6851 270923 6857
rect 270865 6848 270877 6851
rect 268120 6820 270877 6848
rect 262861 6783 262919 6789
rect 262861 6749 262873 6783
rect 262907 6749 262919 6783
rect 262861 6743 262919 6749
rect 263321 6783 263379 6789
rect 263321 6749 263333 6783
rect 263367 6780 263379 6783
rect 263502 6780 263508 6792
rect 263367 6752 263508 6780
rect 263367 6749 263379 6752
rect 263321 6743 263379 6749
rect 263502 6740 263508 6752
rect 263560 6740 263566 6792
rect 264054 6740 264060 6792
rect 264112 6740 264118 6792
rect 264238 6740 264244 6792
rect 264296 6780 264302 6792
rect 264793 6783 264851 6789
rect 264793 6780 264805 6783
rect 264296 6752 264805 6780
rect 264296 6740 264302 6752
rect 264793 6749 264805 6752
rect 264839 6749 264851 6783
rect 264793 6743 264851 6749
rect 265526 6740 265532 6792
rect 265584 6740 265590 6792
rect 266998 6740 267004 6792
rect 267056 6780 267062 6792
rect 267185 6783 267243 6789
rect 267185 6780 267197 6783
rect 267056 6752 267197 6780
rect 267056 6740 267062 6752
rect 267185 6749 267197 6752
rect 267231 6749 267243 6783
rect 267185 6743 267243 6749
rect 267369 6783 267427 6789
rect 267369 6749 267381 6783
rect 267415 6780 267427 6783
rect 267415 6752 267780 6780
rect 267415 6749 267427 6752
rect 267369 6743 267427 6749
rect 237116 6684 237328 6712
rect 237466 6672 237472 6724
rect 237524 6712 237530 6724
rect 262122 6712 262128 6724
rect 237524 6684 262128 6712
rect 237524 6672 237530 6684
rect 262122 6672 262128 6684
rect 262180 6672 262186 6724
rect 225432 6616 227392 6644
rect 227717 6647 227775 6653
rect 224957 6607 225015 6613
rect 227717 6613 227729 6647
rect 227763 6644 227775 6647
rect 228085 6647 228143 6653
rect 228085 6644 228097 6647
rect 227763 6616 228097 6644
rect 227763 6613 227775 6616
rect 227717 6607 227775 6613
rect 228085 6613 228097 6616
rect 228131 6644 228143 6647
rect 228174 6644 228180 6656
rect 228131 6616 228180 6644
rect 228131 6613 228143 6616
rect 228085 6607 228143 6613
rect 228174 6604 228180 6616
rect 228232 6604 228238 6656
rect 229925 6647 229983 6653
rect 229925 6613 229937 6647
rect 229971 6644 229983 6647
rect 230474 6644 230480 6656
rect 229971 6616 230480 6644
rect 229971 6613 229983 6616
rect 229925 6607 229983 6613
rect 230474 6604 230480 6616
rect 230532 6604 230538 6656
rect 237374 6604 237380 6656
rect 237432 6604 237438 6656
rect 239122 6604 239128 6656
rect 239180 6644 239186 6656
rect 258626 6644 258632 6656
rect 239180 6616 258632 6644
rect 239180 6604 239186 6616
rect 258626 6604 258632 6616
rect 258684 6604 258690 6656
rect 260190 6604 260196 6656
rect 260248 6604 260254 6656
rect 262033 6647 262091 6653
rect 262033 6613 262045 6647
rect 262079 6644 262091 6647
rect 263410 6644 263416 6656
rect 262079 6616 263416 6644
rect 262079 6613 262091 6616
rect 262033 6607 262091 6613
rect 263410 6604 263416 6616
rect 263468 6604 263474 6656
rect 263505 6647 263563 6653
rect 263505 6613 263517 6647
rect 263551 6644 263563 6647
rect 264146 6644 264152 6656
rect 263551 6616 264152 6644
rect 263551 6613 263563 6616
rect 263505 6607 263563 6613
rect 264146 6604 264152 6616
rect 264204 6604 264210 6656
rect 264241 6647 264299 6653
rect 264241 6613 264253 6647
rect 264287 6644 264299 6647
rect 264422 6644 264428 6656
rect 264287 6616 264428 6644
rect 264287 6613 264299 6616
rect 264241 6607 264299 6613
rect 264422 6604 264428 6616
rect 264480 6604 264486 6656
rect 264698 6604 264704 6656
rect 264756 6644 264762 6656
rect 264977 6647 265035 6653
rect 264977 6644 264989 6647
rect 264756 6616 264989 6644
rect 264756 6604 264762 6616
rect 264977 6613 264989 6616
rect 265023 6613 265035 6647
rect 264977 6607 265035 6613
rect 265710 6604 265716 6656
rect 265768 6604 265774 6656
rect 265802 6604 265808 6656
rect 265860 6644 265866 6656
rect 267553 6647 267611 6653
rect 267553 6644 267565 6647
rect 265860 6616 267565 6644
rect 265860 6604 265866 6616
rect 267553 6613 267565 6616
rect 267599 6613 267611 6647
rect 267752 6644 267780 6752
rect 267826 6740 267832 6792
rect 267884 6780 267890 6792
rect 268120 6789 268148 6820
rect 270865 6817 270877 6820
rect 270911 6817 270923 6851
rect 270865 6811 270923 6817
rect 268105 6783 268163 6789
rect 267884 6752 268056 6780
rect 267884 6740 267890 6752
rect 268028 6712 268056 6752
rect 268105 6749 268117 6783
rect 268151 6749 268163 6783
rect 268105 6743 268163 6749
rect 269206 6740 269212 6792
rect 269264 6740 269270 6792
rect 269482 6740 269488 6792
rect 269540 6740 269546 6792
rect 270494 6740 270500 6792
rect 270552 6740 270558 6792
rect 270681 6783 270739 6789
rect 270681 6749 270693 6783
rect 270727 6749 270739 6783
rect 270681 6743 270739 6749
rect 268473 6715 268531 6721
rect 268473 6712 268485 6715
rect 268028 6684 268485 6712
rect 268473 6681 268485 6684
rect 268519 6681 268531 6715
rect 268473 6675 268531 6681
rect 269500 6712 269528 6740
rect 270402 6712 270408 6724
rect 269500 6684 270408 6712
rect 269500 6644 269528 6684
rect 270402 6672 270408 6684
rect 270460 6712 270466 6724
rect 270696 6712 270724 6743
rect 270460 6684 270724 6712
rect 270460 6672 270466 6684
rect 267752 6616 269528 6644
rect 267553 6607 267611 6613
rect 1104 6554 271651 6576
rect 1104 6502 68546 6554
rect 68598 6502 68610 6554
rect 68662 6502 68674 6554
rect 68726 6502 68738 6554
rect 68790 6502 68802 6554
rect 68854 6502 136143 6554
rect 136195 6502 136207 6554
rect 136259 6502 136271 6554
rect 136323 6502 136335 6554
rect 136387 6502 136399 6554
rect 136451 6502 203740 6554
rect 203792 6502 203804 6554
rect 203856 6502 203868 6554
rect 203920 6502 203932 6554
rect 203984 6502 203996 6554
rect 204048 6502 271337 6554
rect 271389 6502 271401 6554
rect 271453 6502 271465 6554
rect 271517 6502 271529 6554
rect 271581 6502 271593 6554
rect 271645 6502 271651 6554
rect 1104 6480 271651 6502
rect 15562 6400 15568 6452
rect 15620 6440 15626 6452
rect 42610 6440 42616 6452
rect 15620 6412 42616 6440
rect 15620 6400 15626 6412
rect 42610 6400 42616 6412
rect 42668 6400 42674 6452
rect 42720 6412 43576 6440
rect 13722 6332 13728 6384
rect 13780 6372 13786 6384
rect 36538 6372 36544 6384
rect 13780 6344 36544 6372
rect 13780 6332 13786 6344
rect 36538 6332 36544 6344
rect 36596 6332 36602 6384
rect 9950 6264 9956 6316
rect 10008 6304 10014 6316
rect 42720 6304 42748 6412
rect 42797 6375 42855 6381
rect 42797 6341 42809 6375
rect 42843 6372 42855 6375
rect 42978 6372 42984 6384
rect 42843 6344 42984 6372
rect 42843 6341 42855 6344
rect 42797 6335 42855 6341
rect 42978 6332 42984 6344
rect 43036 6332 43042 6384
rect 43073 6375 43131 6381
rect 43073 6341 43085 6375
rect 43119 6372 43131 6375
rect 43346 6372 43352 6384
rect 43119 6344 43352 6372
rect 43119 6341 43131 6344
rect 43073 6335 43131 6341
rect 43346 6332 43352 6344
rect 43404 6332 43410 6384
rect 43548 6372 43576 6412
rect 46014 6400 46020 6452
rect 46072 6440 46078 6452
rect 46109 6443 46167 6449
rect 46109 6440 46121 6443
rect 46072 6412 46121 6440
rect 46072 6400 46078 6412
rect 46109 6409 46121 6412
rect 46155 6440 46167 6443
rect 46661 6443 46719 6449
rect 46661 6440 46673 6443
rect 46155 6412 46673 6440
rect 46155 6409 46167 6412
rect 46109 6403 46167 6409
rect 46661 6409 46673 6412
rect 46707 6409 46719 6443
rect 46661 6403 46719 6409
rect 72326 6400 72332 6452
rect 72384 6440 72390 6452
rect 72384 6412 79548 6440
rect 72384 6400 72390 6412
rect 43548 6344 43852 6372
rect 10008 6276 42748 6304
rect 10008 6264 10014 6276
rect 43162 6264 43168 6316
rect 43220 6264 43226 6316
rect 43548 6313 43576 6344
rect 43533 6307 43591 6313
rect 43533 6273 43545 6307
rect 43579 6273 43591 6307
rect 43824 6304 43852 6344
rect 43898 6332 43904 6384
rect 43956 6332 43962 6384
rect 45002 6332 45008 6384
rect 45060 6332 45066 6384
rect 45281 6375 45339 6381
rect 45281 6341 45293 6375
rect 45327 6372 45339 6375
rect 45554 6372 45560 6384
rect 45327 6344 45560 6372
rect 45327 6341 45339 6344
rect 45281 6335 45339 6341
rect 45554 6332 45560 6344
rect 45612 6332 45618 6384
rect 45738 6332 45744 6384
rect 45796 6332 45802 6384
rect 79318 6332 79324 6384
rect 79376 6372 79382 6384
rect 79413 6375 79471 6381
rect 79413 6372 79425 6375
rect 79376 6344 79425 6372
rect 79376 6332 79382 6344
rect 79413 6341 79425 6344
rect 79459 6341 79471 6375
rect 79520 6372 79548 6412
rect 79594 6400 79600 6452
rect 79652 6400 79658 6452
rect 99006 6440 99012 6452
rect 79704 6412 99012 6440
rect 79704 6372 79732 6412
rect 99006 6400 99012 6412
rect 99064 6400 99070 6452
rect 100110 6400 100116 6452
rect 100168 6400 100174 6452
rect 100202 6400 100208 6452
rect 100260 6440 100266 6452
rect 100297 6443 100355 6449
rect 100297 6440 100309 6443
rect 100260 6412 100309 6440
rect 100260 6400 100266 6412
rect 100297 6409 100309 6412
rect 100343 6409 100355 6443
rect 100297 6403 100355 6409
rect 100754 6400 100760 6452
rect 100812 6440 100818 6452
rect 104710 6440 104716 6452
rect 100812 6412 104716 6440
rect 100812 6400 100818 6412
rect 104710 6400 104716 6412
rect 104768 6400 104774 6452
rect 107286 6400 107292 6452
rect 107344 6440 107350 6452
rect 108574 6440 108580 6452
rect 107344 6412 108580 6440
rect 107344 6400 107350 6412
rect 108574 6400 108580 6412
rect 108632 6440 108638 6452
rect 109310 6440 109316 6452
rect 108632 6412 109316 6440
rect 108632 6400 108638 6412
rect 109310 6400 109316 6412
rect 109368 6400 109374 6452
rect 111242 6400 111248 6452
rect 111300 6440 111306 6452
rect 144454 6440 144460 6452
rect 111300 6412 144460 6440
rect 111300 6400 111306 6412
rect 144454 6400 144460 6412
rect 144512 6400 144518 6452
rect 148042 6400 148048 6452
rect 148100 6440 148106 6452
rect 162486 6440 162492 6452
rect 148100 6412 162492 6440
rect 148100 6400 148106 6412
rect 162486 6400 162492 6412
rect 162544 6400 162550 6452
rect 162578 6400 162584 6452
rect 162636 6440 162642 6452
rect 168282 6440 168288 6452
rect 162636 6412 168288 6440
rect 162636 6400 162642 6412
rect 168282 6400 168288 6412
rect 168340 6400 168346 6452
rect 181806 6400 181812 6452
rect 181864 6400 181870 6452
rect 189166 6440 189172 6452
rect 189224 6449 189230 6452
rect 189224 6443 189243 6449
rect 181916 6412 189172 6440
rect 79520 6344 79732 6372
rect 79413 6335 79471 6341
rect 81342 6332 81348 6384
rect 81400 6372 81406 6384
rect 91462 6372 91468 6384
rect 81400 6344 91468 6372
rect 81400 6332 81406 6344
rect 91462 6332 91468 6344
rect 91520 6332 91526 6384
rect 100662 6372 100668 6384
rect 91572 6344 100668 6372
rect 44453 6307 44511 6313
rect 44453 6304 44465 6307
rect 43824 6276 44465 6304
rect 43533 6267 43591 6273
rect 44453 6273 44465 6276
rect 44499 6273 44511 6307
rect 44453 6267 44511 6273
rect 45370 6264 45376 6316
rect 45428 6264 45434 6316
rect 87690 6304 87696 6316
rect 79520 6276 87696 6304
rect 46020 6248 46072 6254
rect 23658 6196 23664 6248
rect 23716 6236 23722 6248
rect 40494 6236 40500 6248
rect 23716 6208 40500 6236
rect 23716 6196 23722 6208
rect 40494 6196 40500 6208
rect 40552 6196 40558 6248
rect 44726 6236 44732 6248
rect 43838 6208 44732 6236
rect 44726 6196 44732 6208
rect 44784 6196 44790 6248
rect 47578 6236 47584 6248
rect 46072 6208 47584 6236
rect 47578 6196 47584 6208
rect 47636 6196 47642 6248
rect 71590 6196 71596 6248
rect 71648 6236 71654 6248
rect 79520 6236 79548 6276
rect 87690 6264 87696 6276
rect 87748 6264 87754 6316
rect 91572 6304 91600 6344
rect 100662 6332 100668 6344
rect 100720 6332 100726 6384
rect 108114 6372 108120 6384
rect 101692 6344 108120 6372
rect 87800 6276 91600 6304
rect 87800 6236 87828 6276
rect 99926 6264 99932 6316
rect 99984 6304 99990 6316
rect 101692 6304 101720 6344
rect 108114 6332 108120 6344
rect 108172 6332 108178 6384
rect 112070 6372 112076 6384
rect 109006 6344 112076 6372
rect 99984 6276 101720 6304
rect 99984 6264 99990 6276
rect 101766 6264 101772 6316
rect 101824 6264 101830 6316
rect 106366 6264 106372 6316
rect 106424 6304 106430 6316
rect 106921 6307 106979 6313
rect 106921 6304 106933 6307
rect 106424 6276 106933 6304
rect 106424 6264 106430 6276
rect 106921 6273 106933 6276
rect 106967 6273 106979 6307
rect 106921 6267 106979 6273
rect 108666 6264 108672 6316
rect 108724 6304 108730 6316
rect 108761 6307 108819 6313
rect 108761 6304 108773 6307
rect 108724 6276 108773 6304
rect 108724 6264 108730 6276
rect 108761 6273 108773 6276
rect 108807 6273 108819 6307
rect 108761 6267 108819 6273
rect 91557 6239 91615 6245
rect 91557 6236 91569 6239
rect 71648 6208 79548 6236
rect 84166 6208 87828 6236
rect 89686 6208 91569 6236
rect 71648 6196 71654 6208
rect 46020 6190 46072 6196
rect 17218 6128 17224 6180
rect 17276 6168 17282 6180
rect 42518 6168 42524 6180
rect 17276 6140 42524 6168
rect 17276 6128 17282 6140
rect 42518 6128 42524 6140
rect 42576 6128 42582 6180
rect 44082 6128 44088 6180
rect 44140 6128 44146 6180
rect 46293 6171 46351 6177
rect 46293 6137 46305 6171
rect 46339 6168 46351 6171
rect 46339 6140 51074 6168
rect 46339 6137 46351 6140
rect 46293 6131 46351 6137
rect 51046 6100 51074 6140
rect 79042 6128 79048 6180
rect 79100 6128 79106 6180
rect 79336 6140 79548 6168
rect 79336 6100 79364 6140
rect 51046 6072 79364 6100
rect 79410 6060 79416 6112
rect 79468 6060 79474 6112
rect 79520 6100 79548 6140
rect 79686 6128 79692 6180
rect 79744 6168 79750 6180
rect 84166 6168 84194 6208
rect 89686 6168 89714 6208
rect 91557 6205 91569 6208
rect 91603 6205 91615 6239
rect 91557 6199 91615 6205
rect 91741 6239 91799 6245
rect 91741 6205 91753 6239
rect 91787 6236 91799 6239
rect 92750 6236 92756 6248
rect 91787 6208 92756 6236
rect 91787 6205 91799 6208
rect 91741 6199 91799 6205
rect 92750 6196 92756 6208
rect 92808 6196 92814 6248
rect 93394 6196 93400 6248
rect 93452 6196 93458 6248
rect 101953 6239 102011 6245
rect 101953 6205 101965 6239
rect 101999 6205 102011 6239
rect 101953 6199 102011 6205
rect 79744 6140 84194 6168
rect 87984 6140 89714 6168
rect 90913 6171 90971 6177
rect 79744 6128 79750 6140
rect 87984 6100 88012 6140
rect 90913 6137 90925 6171
rect 90959 6168 90971 6171
rect 91281 6171 91339 6177
rect 91281 6168 91293 6171
rect 90959 6140 91293 6168
rect 90959 6137 90971 6140
rect 90913 6131 90971 6137
rect 91281 6137 91293 6140
rect 91327 6168 91339 6171
rect 93412 6168 93440 6196
rect 91327 6140 93440 6168
rect 91327 6137 91339 6140
rect 91281 6131 91339 6137
rect 99742 6128 99748 6180
rect 99800 6128 99806 6180
rect 79520 6072 88012 6100
rect 90266 6060 90272 6112
rect 90324 6100 90330 6112
rect 96798 6100 96804 6112
rect 90324 6072 96804 6100
rect 90324 6060 90330 6072
rect 96798 6060 96804 6072
rect 96856 6060 96862 6112
rect 100110 6060 100116 6112
rect 100168 6060 100174 6112
rect 101968 6100 101996 6199
rect 102226 6196 102232 6248
rect 102284 6196 102290 6248
rect 104710 6196 104716 6248
rect 104768 6236 104774 6248
rect 107105 6239 107163 6245
rect 107105 6236 107117 6239
rect 104768 6208 107117 6236
rect 104768 6196 104774 6208
rect 107105 6205 107117 6208
rect 107151 6236 107163 6239
rect 109006 6236 109034 6344
rect 112070 6332 112076 6344
rect 112128 6332 112134 6384
rect 115934 6332 115940 6384
rect 115992 6372 115998 6384
rect 119893 6375 119951 6381
rect 119893 6372 119905 6375
rect 115992 6344 119905 6372
rect 115992 6332 115998 6344
rect 119893 6341 119905 6344
rect 119939 6341 119951 6375
rect 119893 6335 119951 6341
rect 109954 6264 109960 6316
rect 110012 6304 110018 6316
rect 110877 6307 110935 6313
rect 110877 6304 110889 6307
rect 110012 6276 110889 6304
rect 110012 6264 110018 6276
rect 110877 6273 110889 6276
rect 110923 6273 110935 6307
rect 110877 6267 110935 6273
rect 112714 6264 112720 6316
rect 112772 6264 112778 6316
rect 119908 6304 119936 6335
rect 119982 6332 119988 6384
rect 120040 6372 120046 6384
rect 120093 6375 120151 6381
rect 120093 6372 120105 6375
rect 120040 6344 120105 6372
rect 120040 6332 120046 6344
rect 120093 6341 120105 6344
rect 120139 6372 120151 6375
rect 121089 6375 121147 6381
rect 121089 6372 121101 6375
rect 120139 6344 121101 6372
rect 120139 6341 120151 6344
rect 120093 6335 120151 6341
rect 121089 6341 121101 6344
rect 121135 6341 121147 6375
rect 130194 6372 130200 6384
rect 121089 6335 121147 6341
rect 121932 6344 130200 6372
rect 120721 6307 120779 6313
rect 120721 6304 120733 6307
rect 119908 6276 120733 6304
rect 120721 6273 120733 6276
rect 120767 6304 120779 6307
rect 121932 6304 121960 6344
rect 130194 6332 130200 6344
rect 130252 6332 130258 6384
rect 130286 6332 130292 6384
rect 130344 6332 130350 6384
rect 141326 6332 141332 6384
rect 141384 6372 141390 6384
rect 143442 6372 143448 6384
rect 141384 6344 143448 6372
rect 141384 6332 141390 6344
rect 143442 6332 143448 6344
rect 143500 6332 143506 6384
rect 147490 6372 147496 6384
rect 146496 6344 147496 6372
rect 120767 6276 121960 6304
rect 120767 6273 120779 6276
rect 120721 6267 120779 6273
rect 122098 6264 122104 6316
rect 122156 6304 122162 6316
rect 122156 6276 122328 6304
rect 122156 6264 122162 6276
rect 109310 6236 109316 6248
rect 107151 6208 109316 6236
rect 107151 6205 107163 6208
rect 107105 6199 107163 6205
rect 109310 6196 109316 6208
rect 109368 6196 109374 6248
rect 111061 6239 111119 6245
rect 111061 6205 111073 6239
rect 111107 6236 111119 6239
rect 112622 6236 112628 6248
rect 111107 6208 112628 6236
rect 111107 6205 111119 6208
rect 111061 6199 111119 6205
rect 112622 6196 112628 6208
rect 112680 6196 112686 6248
rect 119062 6196 119068 6248
rect 119120 6236 119126 6248
rect 119341 6239 119399 6245
rect 119341 6236 119353 6239
rect 119120 6208 119353 6236
rect 119120 6196 119126 6208
rect 119341 6205 119353 6208
rect 119387 6236 119399 6239
rect 122006 6236 122012 6248
rect 119387 6208 122012 6236
rect 119387 6205 119399 6208
rect 119341 6199 119399 6205
rect 122006 6196 122012 6208
rect 122064 6196 122070 6248
rect 122300 6236 122328 6276
rect 125134 6264 125140 6316
rect 125192 6264 125198 6316
rect 129918 6264 129924 6316
rect 129976 6304 129982 6316
rect 146496 6313 146524 6344
rect 147490 6332 147496 6344
rect 147548 6332 147554 6384
rect 147674 6332 147680 6384
rect 147732 6372 147738 6384
rect 148778 6372 148784 6384
rect 147732 6344 148784 6372
rect 147732 6332 147738 6344
rect 148778 6332 148784 6344
rect 148836 6372 148842 6384
rect 148962 6372 148968 6384
rect 148836 6344 148968 6372
rect 148836 6332 148842 6344
rect 148962 6332 148968 6344
rect 149020 6372 149026 6384
rect 150710 6372 150716 6384
rect 149020 6344 150716 6372
rect 149020 6332 149026 6344
rect 150710 6332 150716 6344
rect 150768 6332 150774 6384
rect 152642 6332 152648 6384
rect 152700 6332 152706 6384
rect 152734 6332 152740 6384
rect 152792 6372 152798 6384
rect 162854 6372 162860 6384
rect 152792 6344 162860 6372
rect 152792 6332 152798 6344
rect 162854 6332 162860 6344
rect 162912 6332 162918 6384
rect 177850 6372 177856 6384
rect 171106 6344 177856 6372
rect 130657 6307 130715 6313
rect 130657 6304 130669 6307
rect 129976 6276 130669 6304
rect 129976 6264 129982 6276
rect 130657 6273 130669 6276
rect 130703 6273 130715 6307
rect 146481 6307 146539 6313
rect 130657 6267 130715 6273
rect 137986 6276 142844 6304
rect 125413 6239 125471 6245
rect 125413 6236 125425 6239
rect 122300 6208 125425 6236
rect 125413 6205 125425 6208
rect 125459 6236 125471 6239
rect 137986 6236 138014 6276
rect 125459 6208 138014 6236
rect 125459 6205 125471 6208
rect 125413 6199 125471 6205
rect 102244 6168 102272 6196
rect 114370 6168 114376 6180
rect 102244 6140 114376 6168
rect 114370 6128 114376 6140
rect 114428 6128 114434 6180
rect 120258 6128 120264 6180
rect 120316 6128 120322 6180
rect 122098 6168 122104 6180
rect 121104 6140 122104 6168
rect 103146 6100 103152 6112
rect 101968 6072 103152 6100
rect 103146 6060 103152 6072
rect 103204 6060 103210 6112
rect 107654 6060 107660 6112
rect 107712 6100 107718 6112
rect 108758 6100 108764 6112
rect 107712 6072 108764 6100
rect 107712 6060 107718 6072
rect 108758 6060 108764 6072
rect 108816 6060 108822 6112
rect 112070 6060 112076 6112
rect 112128 6100 112134 6112
rect 115842 6100 115848 6112
rect 112128 6072 115848 6100
rect 112128 6060 112134 6072
rect 115842 6060 115848 6072
rect 115900 6060 115906 6112
rect 120074 6060 120080 6112
rect 120132 6100 120138 6112
rect 121104 6109 121132 6140
rect 122098 6128 122104 6140
rect 122156 6128 122162 6180
rect 122190 6128 122196 6180
rect 122248 6168 122254 6180
rect 122248 6140 122696 6168
rect 122248 6128 122254 6140
rect 121089 6103 121147 6109
rect 121089 6100 121101 6103
rect 120132 6072 121101 6100
rect 120132 6060 120138 6072
rect 121089 6069 121101 6072
rect 121135 6069 121147 6103
rect 121089 6063 121147 6069
rect 121273 6103 121331 6109
rect 121273 6069 121285 6103
rect 121319 6100 121331 6103
rect 122558 6100 122564 6112
rect 121319 6072 122564 6100
rect 121319 6069 121331 6072
rect 121273 6063 121331 6069
rect 122558 6060 122564 6072
rect 122616 6060 122622 6112
rect 122668 6100 122696 6140
rect 125594 6128 125600 6180
rect 125652 6168 125658 6180
rect 142614 6168 142620 6180
rect 125652 6140 142620 6168
rect 125652 6128 125658 6140
rect 142614 6128 142620 6140
rect 142672 6128 142678 6180
rect 142816 6168 142844 6276
rect 146481 6273 146493 6307
rect 146527 6273 146539 6307
rect 146481 6267 146539 6273
rect 148060 6276 148456 6304
rect 143350 6196 143356 6248
rect 143408 6236 143414 6248
rect 146665 6239 146723 6245
rect 146665 6236 146677 6239
rect 143408 6208 146677 6236
rect 143408 6196 143414 6208
rect 146665 6205 146677 6208
rect 146711 6236 146723 6239
rect 148060 6236 148088 6276
rect 148428 6248 148456 6276
rect 148870 6264 148876 6316
rect 148928 6264 148934 6316
rect 150066 6264 150072 6316
rect 150124 6304 150130 6316
rect 150805 6307 150863 6313
rect 150805 6304 150817 6307
rect 150124 6276 150817 6304
rect 150124 6264 150130 6276
rect 150805 6273 150817 6276
rect 150851 6273 150863 6307
rect 150805 6267 150863 6273
rect 156049 6307 156107 6313
rect 156049 6273 156061 6307
rect 156095 6304 156107 6307
rect 156138 6304 156144 6316
rect 156095 6276 156144 6304
rect 156095 6273 156107 6276
rect 156049 6267 156107 6273
rect 156138 6264 156144 6276
rect 156196 6264 156202 6316
rect 156782 6264 156788 6316
rect 156840 6304 156846 6316
rect 156877 6307 156935 6313
rect 156877 6304 156889 6307
rect 156840 6276 156889 6304
rect 156840 6264 156846 6276
rect 156877 6273 156889 6276
rect 156923 6273 156935 6307
rect 156877 6267 156935 6273
rect 156966 6264 156972 6316
rect 157024 6304 157030 6316
rect 158162 6304 158168 6316
rect 157024 6276 158168 6304
rect 157024 6264 157030 6276
rect 158162 6264 158168 6276
rect 158220 6264 158226 6316
rect 171106 6304 171134 6344
rect 177850 6332 177856 6344
rect 177908 6332 177914 6384
rect 180978 6332 180984 6384
rect 181036 6372 181042 6384
rect 181916 6372 181944 6412
rect 189166 6400 189172 6412
rect 189231 6409 189243 6443
rect 189224 6403 189243 6409
rect 189224 6400 189230 6403
rect 189350 6400 189356 6452
rect 189408 6400 189414 6452
rect 216766 6440 216772 6452
rect 190426 6412 216772 6440
rect 182174 6372 182180 6384
rect 181036 6344 181944 6372
rect 182008 6344 182180 6372
rect 181036 6332 181042 6344
rect 182008 6313 182036 6344
rect 182174 6332 182180 6344
rect 182232 6372 182238 6384
rect 182232 6344 186314 6372
rect 182232 6332 182238 6344
rect 158272 6276 171134 6304
rect 181809 6307 181867 6313
rect 146711 6208 148088 6236
rect 146711 6205 146723 6208
rect 146665 6199 146723 6205
rect 148134 6196 148140 6248
rect 148192 6196 148198 6248
rect 148410 6196 148416 6248
rect 148468 6236 148474 6248
rect 149241 6239 149299 6245
rect 149241 6236 149253 6239
rect 148468 6208 149253 6236
rect 148468 6196 148474 6208
rect 149241 6205 149253 6208
rect 149287 6205 149299 6239
rect 149241 6199 149299 6205
rect 150986 6196 150992 6248
rect 151044 6236 151050 6248
rect 153286 6236 153292 6248
rect 151044 6208 153292 6236
rect 151044 6196 151050 6208
rect 153286 6196 153292 6208
rect 153344 6196 153350 6248
rect 157058 6196 157064 6248
rect 157116 6196 157122 6248
rect 157242 6196 157248 6248
rect 157300 6236 157306 6248
rect 158272 6236 158300 6276
rect 181809 6273 181821 6307
rect 181855 6273 181867 6307
rect 181809 6267 181867 6273
rect 181993 6307 182051 6313
rect 181993 6273 182005 6307
rect 182039 6273 182051 6307
rect 181993 6267 182051 6273
rect 157300 6208 158300 6236
rect 157300 6196 157306 6208
rect 161566 6196 161572 6248
rect 161624 6236 161630 6248
rect 162578 6236 162584 6248
rect 161624 6208 162584 6236
rect 161624 6196 161630 6208
rect 162578 6196 162584 6208
rect 162636 6196 162642 6248
rect 162854 6196 162860 6248
rect 162912 6236 162918 6248
rect 181824 6236 181852 6267
rect 182542 6264 182548 6316
rect 182600 6264 182606 6316
rect 186286 6304 186314 6344
rect 188430 6332 188436 6384
rect 188488 6372 188494 6384
rect 188985 6375 189043 6381
rect 188985 6372 188997 6375
rect 188488 6344 188997 6372
rect 188488 6332 188494 6344
rect 188985 6341 188997 6344
rect 189031 6341 189043 6375
rect 190426 6372 190454 6412
rect 216766 6400 216772 6412
rect 216824 6400 216830 6452
rect 218330 6400 218336 6452
rect 218388 6440 218394 6452
rect 219894 6440 219900 6452
rect 218388 6412 219900 6440
rect 218388 6400 218394 6412
rect 219894 6400 219900 6412
rect 219952 6400 219958 6452
rect 219989 6443 220047 6449
rect 219989 6409 220001 6443
rect 220035 6440 220047 6443
rect 221182 6440 221188 6452
rect 220035 6412 221188 6440
rect 220035 6409 220047 6412
rect 219989 6403 220047 6409
rect 221182 6400 221188 6412
rect 221240 6440 221246 6452
rect 221240 6412 225552 6440
rect 221240 6400 221246 6412
rect 212074 6372 212080 6384
rect 188985 6335 189043 6341
rect 189092 6344 190454 6372
rect 207584 6344 212080 6372
rect 189092 6304 189120 6344
rect 200758 6304 200764 6316
rect 186286 6276 189120 6304
rect 190426 6276 200764 6304
rect 182082 6236 182088 6248
rect 162912 6208 176654 6236
rect 181824 6208 182088 6236
rect 162912 6196 162918 6208
rect 169202 6168 169208 6180
rect 142816 6140 169208 6168
rect 169202 6128 169208 6140
rect 169260 6128 169266 6180
rect 176626 6168 176654 6208
rect 182082 6196 182088 6208
rect 182140 6196 182146 6248
rect 190426 6168 190454 6276
rect 200758 6264 200764 6276
rect 200816 6264 200822 6316
rect 207584 6313 207612 6344
rect 212074 6332 212080 6344
rect 212132 6332 212138 6384
rect 217870 6372 217876 6384
rect 214208 6344 217876 6372
rect 214208 6313 214236 6344
rect 217870 6332 217876 6344
rect 217928 6332 217934 6384
rect 222102 6332 222108 6384
rect 222160 6372 222166 6384
rect 223850 6372 223856 6384
rect 222160 6344 223856 6372
rect 222160 6332 222166 6344
rect 223850 6332 223856 6344
rect 223908 6372 223914 6384
rect 224126 6372 224132 6384
rect 223908 6344 224132 6372
rect 223908 6332 223914 6344
rect 224126 6332 224132 6344
rect 224184 6372 224190 6384
rect 225322 6372 225328 6384
rect 224184 6344 225328 6372
rect 224184 6332 224190 6344
rect 225322 6332 225328 6344
rect 225380 6332 225386 6384
rect 225524 6372 225552 6412
rect 225598 6400 225604 6452
rect 225656 6440 225662 6452
rect 254762 6440 254768 6452
rect 225656 6412 254768 6440
rect 225656 6400 225662 6412
rect 254762 6400 254768 6412
rect 254820 6400 254826 6452
rect 258626 6400 258632 6452
rect 258684 6440 258690 6452
rect 262950 6440 262956 6452
rect 258684 6412 262956 6440
rect 258684 6400 258690 6412
rect 262950 6400 262956 6412
rect 263008 6400 263014 6452
rect 263410 6400 263416 6452
rect 263468 6400 263474 6452
rect 263502 6400 263508 6452
rect 263560 6440 263566 6452
rect 265618 6440 265624 6452
rect 263560 6412 265624 6440
rect 263560 6400 263566 6412
rect 265618 6400 265624 6412
rect 265676 6400 265682 6452
rect 266170 6400 266176 6452
rect 266228 6440 266234 6452
rect 269206 6440 269212 6452
rect 266228 6412 269212 6440
rect 266228 6400 266234 6412
rect 269206 6400 269212 6412
rect 269264 6400 269270 6452
rect 226978 6372 226984 6384
rect 225524 6344 226984 6372
rect 226978 6332 226984 6344
rect 227036 6332 227042 6384
rect 227714 6332 227720 6384
rect 227772 6372 227778 6384
rect 244274 6372 244280 6384
rect 227772 6344 244280 6372
rect 227772 6332 227778 6344
rect 244274 6332 244280 6344
rect 244332 6332 244338 6384
rect 264698 6372 264704 6384
rect 262508 6344 264704 6372
rect 262508 6316 262536 6344
rect 264698 6332 264704 6344
rect 264756 6332 264762 6384
rect 270865 6375 270923 6381
rect 270865 6372 270877 6375
rect 266648 6344 270877 6372
rect 207569 6307 207627 6313
rect 207569 6273 207581 6307
rect 207615 6273 207627 6307
rect 207569 6267 207627 6273
rect 214193 6307 214251 6313
rect 214193 6273 214205 6307
rect 214239 6273 214251 6307
rect 214193 6267 214251 6273
rect 217778 6264 217784 6316
rect 217836 6264 217842 6316
rect 221182 6264 221188 6316
rect 221240 6264 221246 6316
rect 221366 6313 221372 6316
rect 221323 6307 221372 6313
rect 221323 6273 221335 6307
rect 221369 6273 221372 6307
rect 221323 6267 221372 6273
rect 221366 6264 221372 6267
rect 221424 6264 221430 6316
rect 221458 6264 221464 6316
rect 221516 6264 221522 6316
rect 223025 6307 223083 6313
rect 223025 6273 223037 6307
rect 223071 6304 223083 6307
rect 223390 6304 223396 6316
rect 223071 6276 223396 6304
rect 223071 6273 223083 6276
rect 223025 6267 223083 6273
rect 223390 6264 223396 6276
rect 223448 6264 223454 6316
rect 223666 6264 223672 6316
rect 223724 6264 223730 6316
rect 225509 6307 225567 6313
rect 225509 6304 225521 6307
rect 225248 6276 225521 6304
rect 207750 6196 207756 6248
rect 207808 6196 207814 6248
rect 208394 6196 208400 6248
rect 208452 6236 208458 6248
rect 208452 6208 209774 6236
rect 208452 6196 208458 6208
rect 176626 6140 190454 6168
rect 209746 6168 209774 6208
rect 214098 6196 214104 6248
rect 214156 6236 214162 6248
rect 214377 6239 214435 6245
rect 214377 6236 214389 6239
rect 214156 6208 214389 6236
rect 214156 6196 214162 6208
rect 214377 6205 214389 6208
rect 214423 6236 214435 6239
rect 214650 6236 214656 6248
rect 214423 6208 214656 6236
rect 214423 6205 214435 6208
rect 214377 6199 214435 6205
rect 214650 6196 214656 6208
rect 214708 6196 214714 6248
rect 215294 6196 215300 6248
rect 215352 6236 215358 6248
rect 216033 6239 216091 6245
rect 216033 6236 216045 6239
rect 215352 6208 216045 6236
rect 215352 6196 215358 6208
rect 216033 6205 216045 6208
rect 216079 6236 216091 6239
rect 217134 6236 217140 6248
rect 216079 6208 217140 6236
rect 216079 6205 216091 6208
rect 216033 6199 216091 6205
rect 217134 6196 217140 6208
rect 217192 6196 217198 6248
rect 217962 6196 217968 6248
rect 218020 6196 218026 6248
rect 218330 6196 218336 6248
rect 218388 6236 218394 6248
rect 218425 6239 218483 6245
rect 218425 6236 218437 6239
rect 218388 6208 218437 6236
rect 218388 6196 218394 6208
rect 218425 6205 218437 6208
rect 218471 6205 218483 6239
rect 218701 6239 218759 6245
rect 218701 6236 218713 6239
rect 218425 6199 218483 6205
rect 218532 6208 218713 6236
rect 218054 6168 218060 6180
rect 209746 6140 218060 6168
rect 218054 6128 218060 6140
rect 218112 6128 218118 6180
rect 155034 6100 155040 6112
rect 122668 6072 155040 6100
rect 155034 6060 155040 6072
rect 155092 6060 155098 6112
rect 156322 6060 156328 6112
rect 156380 6060 156386 6112
rect 158806 6060 158812 6112
rect 158864 6100 158870 6112
rect 169294 6100 169300 6112
rect 158864 6072 169300 6100
rect 158864 6060 158870 6072
rect 169294 6060 169300 6072
rect 169352 6060 169358 6112
rect 189074 6060 189080 6112
rect 189132 6100 189138 6112
rect 189169 6103 189227 6109
rect 189169 6100 189181 6103
rect 189132 6072 189181 6100
rect 189132 6060 189138 6072
rect 189169 6069 189181 6072
rect 189215 6100 189227 6103
rect 206922 6100 206928 6112
rect 189215 6072 206928 6100
rect 189215 6069 189227 6072
rect 189169 6063 189227 6069
rect 206922 6060 206928 6072
rect 206980 6060 206986 6112
rect 218532 6100 218560 6208
rect 218701 6205 218713 6208
rect 218747 6205 218759 6239
rect 218701 6199 218759 6205
rect 218790 6196 218796 6248
rect 218848 6245 218854 6248
rect 218848 6239 218876 6245
rect 218864 6205 218876 6239
rect 218848 6199 218876 6205
rect 218848 6196 218854 6199
rect 218974 6196 218980 6248
rect 219032 6196 219038 6248
rect 219158 6196 219164 6248
rect 219216 6236 219222 6248
rect 220265 6239 220323 6245
rect 220265 6236 220277 6239
rect 219216 6208 220277 6236
rect 219216 6196 219222 6208
rect 220265 6205 220277 6208
rect 220311 6205 220323 6239
rect 220265 6199 220323 6205
rect 220354 6196 220360 6248
rect 220412 6236 220418 6248
rect 220449 6239 220507 6245
rect 220449 6236 220461 6239
rect 220412 6208 220461 6236
rect 220412 6196 220418 6208
rect 220449 6205 220461 6208
rect 220495 6205 220507 6239
rect 220449 6199 220507 6205
rect 220538 6196 220544 6248
rect 220596 6236 220602 6248
rect 220596 6208 223436 6236
rect 220596 6196 220602 6208
rect 219894 6128 219900 6180
rect 219952 6168 219958 6180
rect 220909 6171 220967 6177
rect 220909 6168 220921 6171
rect 219952 6140 220921 6168
rect 219952 6128 219958 6140
rect 220909 6137 220921 6140
rect 220955 6137 220967 6171
rect 220909 6131 220967 6137
rect 219158 6100 219164 6112
rect 218532 6072 219164 6100
rect 219158 6060 219164 6072
rect 219216 6060 219222 6112
rect 219434 6060 219440 6112
rect 219492 6100 219498 6112
rect 219621 6103 219679 6109
rect 219621 6100 219633 6103
rect 219492 6072 219633 6100
rect 219492 6060 219498 6072
rect 219621 6069 219633 6072
rect 219667 6069 219679 6103
rect 219621 6063 219679 6069
rect 220630 6060 220636 6112
rect 220688 6100 220694 6112
rect 222105 6103 222163 6109
rect 222105 6100 222117 6103
rect 220688 6072 222117 6100
rect 220688 6060 220694 6072
rect 222105 6069 222117 6072
rect 222151 6069 222163 6103
rect 223408 6100 223436 6208
rect 223850 6196 223856 6248
rect 223908 6196 223914 6248
rect 224126 6196 224132 6248
rect 224184 6236 224190 6248
rect 225248 6236 225276 6276
rect 225509 6273 225521 6276
rect 225555 6304 225567 6307
rect 225874 6304 225880 6316
rect 225555 6276 225880 6304
rect 225555 6273 225567 6276
rect 225509 6267 225567 6273
rect 225874 6264 225880 6276
rect 225932 6264 225938 6316
rect 226058 6264 226064 6316
rect 226116 6304 226122 6316
rect 230201 6307 230259 6313
rect 230201 6304 230213 6307
rect 226116 6276 226840 6304
rect 226116 6264 226122 6276
rect 224184 6208 225276 6236
rect 224184 6196 224190 6208
rect 225322 6196 225328 6248
rect 225380 6236 225386 6248
rect 226702 6236 226708 6248
rect 225380 6208 226708 6236
rect 225380 6196 225386 6208
rect 226702 6196 226708 6208
rect 226760 6196 226766 6248
rect 226812 6236 226840 6276
rect 227272 6276 230213 6304
rect 227272 6236 227300 6276
rect 230201 6273 230213 6276
rect 230247 6304 230259 6307
rect 230290 6304 230296 6316
rect 230247 6276 230296 6304
rect 230247 6273 230259 6276
rect 230201 6267 230259 6273
rect 230290 6264 230296 6276
rect 230348 6264 230354 6316
rect 231305 6307 231363 6313
rect 231305 6273 231317 6307
rect 231351 6304 231363 6307
rect 235626 6304 235632 6316
rect 231351 6276 235632 6304
rect 231351 6273 231363 6276
rect 231305 6267 231363 6273
rect 235626 6264 235632 6276
rect 235684 6264 235690 6316
rect 236181 6307 236239 6313
rect 236181 6273 236193 6307
rect 236227 6304 236239 6307
rect 237374 6304 237380 6316
rect 236227 6276 237380 6304
rect 236227 6273 236239 6276
rect 236181 6267 236239 6273
rect 237374 6264 237380 6276
rect 237432 6264 237438 6316
rect 261202 6264 261208 6316
rect 261260 6264 261266 6316
rect 262398 6264 262404 6316
rect 262456 6264 262462 6316
rect 262490 6264 262496 6316
rect 262548 6264 262554 6316
rect 263597 6307 263655 6313
rect 263597 6273 263609 6307
rect 263643 6273 263655 6307
rect 263597 6267 263655 6273
rect 226812 6208 227300 6236
rect 228450 6196 228456 6248
rect 228508 6236 228514 6248
rect 231578 6236 231584 6248
rect 228508 6208 231584 6236
rect 228508 6196 228514 6208
rect 231578 6196 231584 6208
rect 231636 6196 231642 6248
rect 231670 6196 231676 6248
rect 231728 6196 231734 6248
rect 231762 6196 231768 6248
rect 231820 6236 231826 6248
rect 236457 6239 236515 6245
rect 236457 6236 236469 6239
rect 231820 6208 236469 6236
rect 231820 6196 231826 6208
rect 236457 6205 236469 6208
rect 236503 6205 236515 6239
rect 236457 6199 236515 6205
rect 261478 6196 261484 6248
rect 261536 6196 261542 6248
rect 224218 6128 224224 6180
rect 224276 6168 224282 6180
rect 226242 6168 226248 6180
rect 224276 6140 226248 6168
rect 224276 6128 224282 6140
rect 226242 6128 226248 6140
rect 226300 6128 226306 6180
rect 226978 6128 226984 6180
rect 227036 6168 227042 6180
rect 252830 6168 252836 6180
rect 227036 6140 252836 6168
rect 227036 6128 227042 6140
rect 252830 6128 252836 6140
rect 252888 6128 252894 6180
rect 260190 6128 260196 6180
rect 260248 6168 260254 6180
rect 263612 6168 263640 6267
rect 264238 6264 264244 6316
rect 264296 6264 264302 6316
rect 264606 6264 264612 6316
rect 264664 6264 264670 6316
rect 265437 6307 265495 6313
rect 265437 6273 265449 6307
rect 265483 6304 265495 6307
rect 265802 6304 265808 6316
rect 265483 6276 265808 6304
rect 265483 6273 265495 6276
rect 265437 6267 265495 6273
rect 265802 6264 265808 6276
rect 265860 6264 265866 6316
rect 266648 6313 266676 6344
rect 270865 6341 270877 6344
rect 270911 6341 270923 6375
rect 270865 6335 270923 6341
rect 266633 6307 266691 6313
rect 266633 6273 266645 6307
rect 266679 6273 266691 6307
rect 266633 6267 266691 6273
rect 267826 6264 267832 6316
rect 267884 6264 267890 6316
rect 268381 6307 268439 6313
rect 268381 6273 268393 6307
rect 268427 6304 268439 6307
rect 268470 6304 268476 6316
rect 268427 6276 268476 6304
rect 268427 6273 268439 6276
rect 268381 6267 268439 6273
rect 268470 6264 268476 6276
rect 268528 6264 268534 6316
rect 269390 6264 269396 6316
rect 269448 6264 269454 6316
rect 270402 6264 270408 6316
rect 270460 6304 270466 6316
rect 270681 6307 270739 6313
rect 270681 6304 270693 6307
rect 270460 6276 270693 6304
rect 270460 6264 270466 6276
rect 270681 6273 270693 6276
rect 270727 6273 270739 6307
rect 270681 6267 270739 6273
rect 265158 6196 265164 6248
rect 265216 6236 265222 6248
rect 265713 6239 265771 6245
rect 265713 6236 265725 6239
rect 265216 6208 265725 6236
rect 265216 6196 265222 6208
rect 265713 6205 265725 6208
rect 265759 6205 265771 6239
rect 265713 6199 265771 6205
rect 266906 6196 266912 6248
rect 266964 6196 266970 6248
rect 269114 6196 269120 6248
rect 269172 6236 269178 6248
rect 269669 6239 269727 6245
rect 269669 6236 269681 6239
rect 269172 6208 269681 6236
rect 269172 6196 269178 6208
rect 269669 6205 269681 6208
rect 269715 6205 269727 6239
rect 269669 6199 269727 6205
rect 270034 6196 270040 6248
rect 270092 6236 270098 6248
rect 270497 6239 270555 6245
rect 270497 6236 270509 6239
rect 270092 6208 270509 6236
rect 270092 6196 270098 6208
rect 270497 6205 270509 6208
rect 270543 6205 270555 6239
rect 270497 6199 270555 6205
rect 268102 6168 268108 6180
rect 260248 6140 262812 6168
rect 263612 6140 268108 6168
rect 260248 6128 260254 6140
rect 226426 6100 226432 6112
rect 223408 6072 226432 6100
rect 222105 6063 222163 6069
rect 226426 6060 226432 6072
rect 226484 6060 226490 6112
rect 226518 6060 226524 6112
rect 226576 6100 226582 6112
rect 227714 6100 227720 6112
rect 226576 6072 227720 6100
rect 226576 6060 226582 6072
rect 227714 6060 227720 6072
rect 227772 6060 227778 6112
rect 229830 6060 229836 6112
rect 229888 6100 229894 6112
rect 230106 6100 230112 6112
rect 229888 6072 230112 6100
rect 229888 6060 229894 6072
rect 230106 6060 230112 6072
rect 230164 6060 230170 6112
rect 230474 6060 230480 6112
rect 230532 6100 230538 6112
rect 230750 6100 230756 6112
rect 230532 6072 230756 6100
rect 230532 6060 230538 6072
rect 230750 6060 230756 6072
rect 230808 6060 230814 6112
rect 231118 6060 231124 6112
rect 231176 6100 231182 6112
rect 238754 6100 238760 6112
rect 231176 6072 238760 6100
rect 231176 6060 231182 6072
rect 238754 6060 238760 6072
rect 238812 6060 238818 6112
rect 261662 6060 261668 6112
rect 261720 6100 261726 6112
rect 262677 6103 262735 6109
rect 262677 6100 262689 6103
rect 261720 6072 262689 6100
rect 261720 6060 261726 6072
rect 262677 6069 262689 6072
rect 262723 6069 262735 6103
rect 262784 6100 262812 6140
rect 268102 6128 268108 6140
rect 268160 6128 268166 6180
rect 266722 6100 266728 6112
rect 262784 6072 266728 6100
rect 262677 6063 262735 6069
rect 266722 6060 266728 6072
rect 266780 6060 266786 6112
rect 267090 6060 267096 6112
rect 267148 6100 267154 6112
rect 269022 6100 269028 6112
rect 267148 6072 269028 6100
rect 267148 6060 267154 6072
rect 269022 6060 269028 6072
rect 269080 6060 269086 6112
rect 270310 6060 270316 6112
rect 270368 6100 270374 6112
rect 271966 6100 271972 6112
rect 270368 6072 271972 6100
rect 270368 6060 270374 6072
rect 271966 6060 271972 6072
rect 272024 6060 272030 6112
rect 1104 6010 271492 6032
rect 1104 5958 34748 6010
rect 34800 5958 34812 6010
rect 34864 5958 34876 6010
rect 34928 5958 34940 6010
rect 34992 5958 35004 6010
rect 35056 5958 102345 6010
rect 102397 5958 102409 6010
rect 102461 5958 102473 6010
rect 102525 5958 102537 6010
rect 102589 5958 102601 6010
rect 102653 5958 169942 6010
rect 169994 5958 170006 6010
rect 170058 5958 170070 6010
rect 170122 5958 170134 6010
rect 170186 5958 170198 6010
rect 170250 5958 237539 6010
rect 237591 5958 237603 6010
rect 237655 5958 237667 6010
rect 237719 5958 237731 6010
rect 237783 5958 237795 6010
rect 237847 5958 271492 6010
rect 1104 5936 271492 5958
rect 36538 5856 36544 5908
rect 36596 5896 36602 5908
rect 42794 5896 42800 5908
rect 36596 5868 42800 5896
rect 36596 5856 36602 5868
rect 42794 5856 42800 5868
rect 42852 5856 42858 5908
rect 47854 5856 47860 5908
rect 47912 5856 47918 5908
rect 79042 5856 79048 5908
rect 79100 5896 79106 5908
rect 79321 5899 79379 5905
rect 79321 5896 79333 5899
rect 79100 5868 79333 5896
rect 79100 5856 79106 5868
rect 79321 5865 79333 5868
rect 79367 5896 79379 5899
rect 99742 5896 99748 5908
rect 79367 5868 99748 5896
rect 79367 5865 79379 5868
rect 79321 5859 79379 5865
rect 99742 5856 99748 5868
rect 99800 5896 99806 5908
rect 120074 5896 120080 5908
rect 99800 5868 120080 5896
rect 99800 5856 99806 5868
rect 120074 5856 120080 5868
rect 120132 5856 120138 5908
rect 162762 5896 162768 5908
rect 128648 5868 162768 5896
rect 77294 5788 77300 5840
rect 77352 5828 77358 5840
rect 79505 5831 79563 5837
rect 79505 5828 79517 5831
rect 77352 5800 79517 5828
rect 77352 5788 77358 5800
rect 79505 5797 79517 5800
rect 79551 5797 79563 5831
rect 79505 5791 79563 5797
rect 84194 5788 84200 5840
rect 84252 5828 84258 5840
rect 84252 5800 89714 5828
rect 84252 5788 84258 5800
rect 47584 5772 47636 5778
rect 33226 5720 33232 5772
rect 33284 5760 33290 5772
rect 44726 5760 44732 5772
rect 33284 5732 43024 5760
rect 44298 5732 44732 5760
rect 33284 5720 33290 5732
rect 42702 5692 42708 5704
rect 22066 5664 42708 5692
rect 11330 5584 11336 5636
rect 11388 5624 11394 5636
rect 22066 5624 22094 5664
rect 42702 5652 42708 5664
rect 42760 5652 42766 5704
rect 11388 5596 22094 5624
rect 11388 5584 11394 5596
rect 42058 5584 42064 5636
rect 42116 5584 42122 5636
rect 42996 5624 43024 5732
rect 44726 5720 44732 5732
rect 44784 5760 44790 5772
rect 46014 5760 46020 5772
rect 44784 5732 46020 5760
rect 44784 5720 44790 5732
rect 46014 5720 46020 5732
rect 46072 5720 46078 5772
rect 48038 5760 48044 5772
rect 47636 5732 48044 5760
rect 48038 5720 48044 5732
rect 48096 5720 48102 5772
rect 51626 5760 51632 5772
rect 51566 5732 51632 5760
rect 51626 5720 51632 5732
rect 51684 5760 51690 5772
rect 53098 5760 53104 5772
rect 51684 5732 53104 5760
rect 51684 5720 51690 5732
rect 53098 5720 53104 5732
rect 53156 5720 53162 5772
rect 78953 5763 79011 5769
rect 78953 5729 78965 5763
rect 78999 5760 79011 5763
rect 79318 5760 79324 5772
rect 78999 5732 79324 5760
rect 78999 5729 79011 5732
rect 78953 5723 79011 5729
rect 79318 5720 79324 5732
rect 79376 5720 79382 5772
rect 80790 5720 80796 5772
rect 80848 5760 80854 5772
rect 81253 5763 81311 5769
rect 81253 5760 81265 5763
rect 80848 5732 81265 5760
rect 80848 5720 80854 5732
rect 81253 5729 81265 5732
rect 81299 5760 81311 5763
rect 81986 5760 81992 5772
rect 81299 5732 81992 5760
rect 81299 5729 81311 5732
rect 81253 5723 81311 5729
rect 81986 5720 81992 5732
rect 82044 5720 82050 5772
rect 84930 5720 84936 5772
rect 84988 5760 84994 5772
rect 87141 5763 87199 5769
rect 87141 5760 87153 5763
rect 84988 5732 87153 5760
rect 84988 5720 84994 5732
rect 87141 5729 87153 5732
rect 87187 5729 87199 5763
rect 89686 5760 89714 5800
rect 93854 5788 93860 5840
rect 93912 5828 93918 5840
rect 93912 5800 100064 5828
rect 93912 5788 93918 5800
rect 99926 5760 99932 5772
rect 89686 5732 99932 5760
rect 87141 5723 87199 5729
rect 99926 5720 99932 5732
rect 99984 5720 99990 5772
rect 100036 5760 100064 5800
rect 100110 5788 100116 5840
rect 100168 5828 100174 5840
rect 101033 5831 101091 5837
rect 101033 5828 101045 5831
rect 100168 5800 101045 5828
rect 100168 5788 100174 5800
rect 101033 5797 101045 5800
rect 101079 5828 101091 5831
rect 101079 5800 109356 5828
rect 101079 5797 101091 5800
rect 101033 5791 101091 5797
rect 108850 5760 108856 5772
rect 100036 5732 108856 5760
rect 108850 5720 108856 5732
rect 108908 5720 108914 5772
rect 109034 5720 109040 5772
rect 109092 5720 109098 5772
rect 109328 5760 109356 5800
rect 111242 5788 111248 5840
rect 111300 5788 111306 5840
rect 111518 5788 111524 5840
rect 111576 5828 111582 5840
rect 112441 5831 112499 5837
rect 112441 5828 112453 5831
rect 111576 5800 112453 5828
rect 111576 5788 111582 5800
rect 112441 5797 112453 5800
rect 112487 5828 112499 5831
rect 112809 5831 112867 5837
rect 112809 5828 112821 5831
rect 112487 5800 112821 5828
rect 112487 5797 112499 5800
rect 112441 5791 112499 5797
rect 112809 5797 112821 5800
rect 112855 5828 112867 5831
rect 115106 5828 115112 5840
rect 112855 5800 115112 5828
rect 112855 5797 112867 5800
rect 112809 5791 112867 5797
rect 115106 5788 115112 5800
rect 115164 5828 115170 5840
rect 115293 5831 115351 5837
rect 115293 5828 115305 5831
rect 115164 5800 115305 5828
rect 115164 5788 115170 5800
rect 115293 5797 115305 5800
rect 115339 5828 115351 5831
rect 115661 5831 115719 5837
rect 115661 5828 115673 5831
rect 115339 5800 115673 5828
rect 115339 5797 115351 5800
rect 115293 5791 115351 5797
rect 115661 5797 115673 5800
rect 115707 5828 115719 5831
rect 115750 5828 115756 5840
rect 115707 5800 115756 5828
rect 115707 5797 115719 5800
rect 115661 5791 115719 5797
rect 115750 5788 115756 5800
rect 115808 5788 115814 5840
rect 115842 5788 115848 5840
rect 115900 5828 115906 5840
rect 115900 5800 120304 5828
rect 115900 5788 115906 5800
rect 119982 5760 119988 5772
rect 109328 5732 119988 5760
rect 119982 5720 119988 5732
rect 120040 5720 120046 5772
rect 120276 5769 120304 5800
rect 120261 5763 120319 5769
rect 120261 5729 120273 5763
rect 120307 5729 120319 5763
rect 128648 5760 128676 5868
rect 162762 5856 162768 5868
rect 162820 5856 162826 5908
rect 163038 5856 163044 5908
rect 163096 5896 163102 5908
rect 163096 5868 171134 5896
rect 163096 5856 163102 5868
rect 156966 5828 156972 5840
rect 120261 5723 120319 5729
rect 125060 5732 128676 5760
rect 128832 5800 156972 5828
rect 47584 5714 47636 5720
rect 43438 5652 43444 5704
rect 43496 5692 43502 5704
rect 43533 5695 43591 5701
rect 43533 5692 43545 5695
rect 43496 5664 43545 5692
rect 43496 5652 43502 5664
rect 43533 5661 43545 5664
rect 43579 5661 43591 5695
rect 43533 5655 43591 5661
rect 43622 5652 43628 5704
rect 43680 5652 43686 5704
rect 43714 5652 43720 5704
rect 43772 5692 43778 5704
rect 43993 5695 44051 5701
rect 43993 5692 44005 5695
rect 43772 5664 44005 5692
rect 43772 5652 43778 5664
rect 43993 5661 44005 5664
rect 44039 5661 44051 5695
rect 43993 5655 44051 5661
rect 44358 5652 44364 5704
rect 44416 5701 44422 5704
rect 44416 5695 44433 5701
rect 44421 5661 44433 5695
rect 44416 5655 44433 5661
rect 44416 5652 44422 5655
rect 46842 5652 46848 5704
rect 46900 5652 46906 5704
rect 46934 5652 46940 5704
rect 46992 5652 46998 5704
rect 47302 5652 47308 5704
rect 47360 5652 47366 5704
rect 50430 5652 50436 5704
rect 50488 5692 50494 5704
rect 50801 5695 50859 5701
rect 50801 5692 50813 5695
rect 50488 5664 50813 5692
rect 50488 5652 50494 5664
rect 50801 5661 50813 5664
rect 50847 5661 50859 5695
rect 50801 5655 50859 5661
rect 51074 5652 51080 5704
rect 51132 5692 51138 5704
rect 51261 5695 51319 5701
rect 51261 5692 51273 5695
rect 51132 5664 51273 5692
rect 51132 5652 51138 5664
rect 51261 5661 51273 5664
rect 51307 5661 51319 5695
rect 51261 5655 51319 5661
rect 81434 5652 81440 5704
rect 81492 5652 81498 5704
rect 83369 5695 83427 5701
rect 83369 5661 83381 5695
rect 83415 5661 83427 5695
rect 83369 5655 83427 5661
rect 50893 5627 50951 5633
rect 42996 5596 50660 5624
rect 41322 5516 41328 5568
rect 41380 5556 41386 5568
rect 42153 5559 42211 5565
rect 42153 5556 42165 5559
rect 41380 5528 42165 5556
rect 41380 5516 41386 5528
rect 42153 5525 42165 5528
rect 42199 5525 42211 5559
rect 42153 5519 42211 5525
rect 43257 5559 43315 5565
rect 43257 5525 43269 5559
rect 43303 5556 43315 5559
rect 44450 5556 44456 5568
rect 43303 5528 44456 5556
rect 43303 5525 43315 5528
rect 43257 5519 43315 5525
rect 44450 5516 44456 5528
rect 44508 5516 44514 5568
rect 44542 5516 44548 5568
rect 44600 5516 44606 5568
rect 46569 5559 46627 5565
rect 46569 5525 46581 5559
rect 46615 5556 46627 5559
rect 46658 5556 46664 5568
rect 46615 5528 46664 5556
rect 46615 5525 46627 5528
rect 46569 5519 46627 5525
rect 46658 5516 46664 5528
rect 46716 5516 46722 5568
rect 47670 5516 47676 5568
rect 47728 5516 47734 5568
rect 50522 5516 50528 5568
rect 50580 5516 50586 5568
rect 50632 5556 50660 5596
rect 50893 5593 50905 5627
rect 50939 5624 50951 5627
rect 50982 5624 50988 5636
rect 50939 5596 50988 5624
rect 50939 5593 50951 5596
rect 50893 5587 50951 5593
rect 50982 5584 50988 5596
rect 51040 5584 51046 5636
rect 83384 5624 83412 5655
rect 86770 5652 86776 5704
rect 86828 5692 86834 5704
rect 86865 5695 86923 5701
rect 86865 5692 86877 5695
rect 86828 5664 86877 5692
rect 86828 5652 86834 5664
rect 86865 5661 86877 5664
rect 86911 5692 86923 5695
rect 86911 5664 88104 5692
rect 86911 5661 86923 5664
rect 86865 5655 86923 5661
rect 60706 5596 83412 5624
rect 83553 5627 83611 5633
rect 51629 5559 51687 5565
rect 51629 5556 51641 5559
rect 50632 5528 51641 5556
rect 51629 5525 51641 5528
rect 51675 5525 51687 5559
rect 51629 5519 51687 5525
rect 51813 5559 51871 5565
rect 51813 5525 51825 5559
rect 51859 5556 51871 5559
rect 60706 5556 60734 5596
rect 83553 5593 83565 5627
rect 83599 5624 83611 5627
rect 84930 5624 84936 5636
rect 83599 5596 84936 5624
rect 83599 5593 83611 5596
rect 83553 5587 83611 5593
rect 84930 5584 84936 5596
rect 84988 5584 84994 5636
rect 85209 5627 85267 5633
rect 85209 5593 85221 5627
rect 85255 5624 85267 5627
rect 85574 5624 85580 5636
rect 85255 5596 85580 5624
rect 85255 5593 85267 5596
rect 85209 5587 85267 5593
rect 51859 5528 60734 5556
rect 79321 5559 79379 5565
rect 51859 5525 51871 5528
rect 51813 5519 51871 5525
rect 79321 5525 79333 5559
rect 79367 5556 79379 5559
rect 79410 5556 79416 5568
rect 79367 5528 79416 5556
rect 79367 5525 79379 5528
rect 79321 5519 79379 5525
rect 79410 5516 79416 5528
rect 79468 5556 79474 5568
rect 81621 5559 81679 5565
rect 81621 5556 81633 5559
rect 79468 5528 81633 5556
rect 79468 5516 79474 5528
rect 81621 5525 81633 5528
rect 81667 5525 81679 5559
rect 81621 5519 81679 5525
rect 82725 5559 82783 5565
rect 82725 5525 82737 5559
rect 82771 5556 82783 5559
rect 83093 5559 83151 5565
rect 83093 5556 83105 5559
rect 82771 5528 83105 5556
rect 82771 5525 82783 5528
rect 82725 5519 82783 5525
rect 83093 5525 83105 5528
rect 83139 5556 83151 5559
rect 85224 5556 85252 5587
rect 85574 5584 85580 5596
rect 85632 5584 85638 5636
rect 88076 5568 88104 5664
rect 92658 5652 92664 5704
rect 92716 5652 92722 5704
rect 94498 5652 94504 5704
rect 94556 5652 94562 5704
rect 100389 5695 100447 5701
rect 100389 5661 100401 5695
rect 100435 5692 100447 5695
rect 100570 5692 100576 5704
rect 100435 5664 100576 5692
rect 100435 5661 100447 5664
rect 100389 5655 100447 5661
rect 100570 5652 100576 5664
rect 100628 5692 100634 5704
rect 100665 5695 100723 5701
rect 100665 5692 100677 5695
rect 100628 5664 100677 5692
rect 100628 5652 100634 5664
rect 100665 5661 100677 5664
rect 100711 5661 100723 5695
rect 100665 5655 100723 5661
rect 100849 5695 100907 5701
rect 100849 5661 100861 5695
rect 100895 5692 100907 5695
rect 100938 5692 100944 5704
rect 100895 5664 100944 5692
rect 100895 5661 100907 5664
rect 100849 5655 100907 5661
rect 100938 5652 100944 5664
rect 100996 5652 101002 5704
rect 102137 5695 102195 5701
rect 102137 5661 102149 5695
rect 102183 5692 102195 5695
rect 102778 5692 102784 5704
rect 102183 5664 102784 5692
rect 102183 5661 102195 5664
rect 102137 5655 102195 5661
rect 102778 5652 102784 5664
rect 102836 5692 102842 5704
rect 110877 5695 110935 5701
rect 102836 5664 104664 5692
rect 102836 5652 102842 5664
rect 92842 5584 92848 5636
rect 92900 5584 92906 5636
rect 93394 5584 93400 5636
rect 93452 5624 93458 5636
rect 101858 5624 101864 5636
rect 93452 5596 101864 5624
rect 93452 5584 93458 5596
rect 101858 5584 101864 5596
rect 101916 5584 101922 5636
rect 103146 5584 103152 5636
rect 103204 5584 103210 5636
rect 104636 5624 104664 5664
rect 110877 5661 110889 5695
rect 110923 5692 110935 5695
rect 111242 5692 111248 5704
rect 110923 5664 111248 5692
rect 110923 5661 110935 5664
rect 110877 5655 110935 5661
rect 104710 5624 104716 5636
rect 104636 5596 104716 5624
rect 104710 5584 104716 5596
rect 104768 5584 104774 5636
rect 108393 5627 108451 5633
rect 108393 5624 108405 5627
rect 106246 5596 108405 5624
rect 83139 5528 85252 5556
rect 83139 5525 83151 5528
rect 83093 5519 83151 5525
rect 88058 5516 88064 5568
rect 88116 5556 88122 5568
rect 92474 5556 92480 5568
rect 88116 5528 92480 5556
rect 88116 5516 88122 5528
rect 92474 5516 92480 5528
rect 92532 5556 92538 5568
rect 95050 5556 95056 5568
rect 92532 5528 95056 5556
rect 92532 5516 92538 5528
rect 95050 5516 95056 5528
rect 95108 5516 95114 5568
rect 102042 5516 102048 5568
rect 102100 5556 102106 5568
rect 106246 5556 106274 5596
rect 108393 5593 108405 5596
rect 108439 5624 108451 5627
rect 108761 5627 108819 5633
rect 108761 5624 108773 5627
rect 108439 5596 108773 5624
rect 108439 5593 108451 5596
rect 108393 5587 108451 5593
rect 108761 5593 108773 5596
rect 108807 5624 108819 5627
rect 109221 5627 109279 5633
rect 108807 5596 109172 5624
rect 108807 5593 108819 5596
rect 108761 5587 108819 5593
rect 102100 5528 106274 5556
rect 109144 5556 109172 5596
rect 109221 5593 109233 5627
rect 109267 5624 109279 5627
rect 109310 5624 109316 5636
rect 109267 5596 109316 5624
rect 109267 5593 109279 5596
rect 109221 5587 109279 5593
rect 109310 5584 109316 5596
rect 109368 5584 109374 5636
rect 110892 5556 110920 5655
rect 111242 5652 111248 5664
rect 111300 5652 111306 5704
rect 111794 5652 111800 5704
rect 111852 5692 111858 5704
rect 113177 5695 113235 5701
rect 113177 5692 113189 5695
rect 111852 5664 113189 5692
rect 111852 5652 111858 5664
rect 113177 5661 113189 5664
rect 113223 5661 113235 5695
rect 113177 5655 113235 5661
rect 115017 5695 115075 5701
rect 115017 5661 115029 5695
rect 115063 5692 115075 5695
rect 115106 5692 115112 5704
rect 115063 5664 115112 5692
rect 115063 5661 115075 5664
rect 115017 5655 115075 5661
rect 115106 5652 115112 5664
rect 115164 5652 115170 5704
rect 116762 5652 116768 5704
rect 116820 5692 116826 5704
rect 119062 5692 119068 5704
rect 116820 5664 119068 5692
rect 116820 5652 116826 5664
rect 119062 5652 119068 5664
rect 119120 5652 119126 5704
rect 120074 5652 120080 5704
rect 120132 5652 120138 5704
rect 125060 5701 125088 5732
rect 125045 5695 125103 5701
rect 125045 5661 125057 5695
rect 125091 5661 125103 5695
rect 128832 5692 128860 5800
rect 156966 5788 156972 5800
rect 157024 5788 157030 5840
rect 163056 5828 163084 5856
rect 161032 5800 163084 5828
rect 171106 5828 171134 5868
rect 180978 5856 180984 5908
rect 181036 5856 181042 5908
rect 182910 5856 182916 5908
rect 182968 5856 182974 5908
rect 216030 5896 216036 5908
rect 190426 5868 216036 5896
rect 181806 5828 181812 5840
rect 171106 5800 181812 5828
rect 130194 5720 130200 5772
rect 130252 5720 130258 5772
rect 143074 5720 143080 5772
rect 143132 5720 143138 5772
rect 143261 5763 143319 5769
rect 143261 5729 143273 5763
rect 143307 5760 143319 5763
rect 143350 5760 143356 5772
rect 143307 5732 143356 5760
rect 143307 5729 143319 5732
rect 143261 5723 143319 5729
rect 143350 5720 143356 5732
rect 143408 5720 143414 5772
rect 143534 5720 143540 5772
rect 143592 5720 143598 5772
rect 144454 5720 144460 5772
rect 144512 5760 144518 5772
rect 147582 5760 147588 5772
rect 144512 5732 147588 5760
rect 144512 5720 144518 5732
rect 147582 5720 147588 5732
rect 147640 5760 147646 5772
rect 147677 5763 147735 5769
rect 147677 5760 147689 5763
rect 147640 5732 147689 5760
rect 147640 5720 147646 5732
rect 147677 5729 147689 5732
rect 147723 5729 147735 5763
rect 147677 5723 147735 5729
rect 148226 5720 148232 5772
rect 148284 5720 148290 5772
rect 150069 5763 150127 5769
rect 150069 5729 150081 5763
rect 150115 5760 150127 5763
rect 150437 5763 150495 5769
rect 150437 5760 150449 5763
rect 150115 5732 150449 5760
rect 150115 5729 150127 5732
rect 150069 5723 150127 5729
rect 150437 5729 150449 5732
rect 150483 5760 150495 5763
rect 150805 5763 150863 5769
rect 150805 5760 150817 5763
rect 150483 5732 150817 5760
rect 150483 5729 150495 5732
rect 150437 5723 150495 5729
rect 150805 5729 150817 5732
rect 150851 5760 150863 5763
rect 152734 5760 152740 5772
rect 150851 5732 152740 5760
rect 150851 5729 150863 5732
rect 150805 5723 150863 5729
rect 125045 5655 125103 5661
rect 128326 5664 128860 5692
rect 112622 5584 112628 5636
rect 112680 5624 112686 5636
rect 113361 5627 113419 5633
rect 113361 5624 113373 5627
rect 112680 5596 113373 5624
rect 112680 5584 112686 5596
rect 113361 5593 113373 5596
rect 113407 5624 113419 5627
rect 114370 5624 114376 5636
rect 113407 5596 114376 5624
rect 113407 5593 113419 5596
rect 113361 5587 113419 5593
rect 114370 5584 114376 5596
rect 114428 5584 114434 5636
rect 119430 5584 119436 5636
rect 119488 5624 119494 5636
rect 119801 5627 119859 5633
rect 119801 5624 119813 5627
rect 119488 5596 119813 5624
rect 119488 5584 119494 5596
rect 119801 5593 119813 5596
rect 119847 5624 119859 5627
rect 121917 5627 121975 5633
rect 121917 5624 121929 5627
rect 119847 5596 121929 5624
rect 119847 5593 119859 5596
rect 119801 5587 119859 5593
rect 121917 5593 121929 5596
rect 121963 5624 121975 5627
rect 122561 5627 122619 5633
rect 122561 5624 122573 5627
rect 121963 5596 122573 5624
rect 121963 5593 121975 5596
rect 121917 5587 121975 5593
rect 122561 5593 122573 5596
rect 122607 5624 122619 5627
rect 128326 5624 128354 5664
rect 129918 5652 129924 5704
rect 129976 5652 129982 5704
rect 145190 5652 145196 5704
rect 145248 5692 145254 5704
rect 148042 5692 148048 5704
rect 145248 5664 148048 5692
rect 145248 5652 145254 5664
rect 148042 5652 148048 5664
rect 148100 5652 148106 5704
rect 122607 5596 128354 5624
rect 122607 5593 122619 5596
rect 122561 5587 122619 5593
rect 142614 5584 142620 5636
rect 142672 5624 142678 5636
rect 143534 5624 143540 5636
rect 142672 5596 143540 5624
rect 142672 5584 142678 5596
rect 143534 5584 143540 5596
rect 143592 5584 143598 5636
rect 148134 5584 148140 5636
rect 148192 5624 148198 5636
rect 148410 5624 148416 5636
rect 148192 5596 148416 5624
rect 148192 5584 148198 5596
rect 148410 5584 148416 5596
rect 148468 5584 148474 5636
rect 109144 5528 110920 5556
rect 102100 5516 102106 5528
rect 122190 5516 122196 5568
rect 122248 5556 122254 5568
rect 125134 5556 125140 5568
rect 122248 5528 125140 5556
rect 122248 5516 122254 5528
rect 125134 5516 125140 5528
rect 125192 5516 125198 5568
rect 147582 5516 147588 5568
rect 147640 5556 147646 5568
rect 150084 5556 150112 5723
rect 152734 5720 152740 5732
rect 152792 5720 152798 5772
rect 153841 5763 153899 5769
rect 153841 5760 153853 5763
rect 152936 5732 153853 5760
rect 152936 5692 152964 5732
rect 153841 5729 153853 5732
rect 153887 5729 153899 5763
rect 153841 5723 153899 5729
rect 155034 5720 155040 5772
rect 155092 5760 155098 5772
rect 155092 5732 157564 5760
rect 155092 5720 155098 5732
rect 152752 5664 152964 5692
rect 147640 5528 150112 5556
rect 147640 5516 147646 5528
rect 151998 5516 152004 5568
rect 152056 5556 152062 5568
rect 152752 5565 152780 5664
rect 153378 5652 153384 5704
rect 153436 5652 153442 5704
rect 155678 5652 155684 5704
rect 155736 5652 155742 5704
rect 157536 5701 157564 5732
rect 157521 5695 157579 5701
rect 157521 5661 157533 5695
rect 157567 5692 157579 5695
rect 157889 5695 157947 5701
rect 157889 5692 157901 5695
rect 157567 5664 157901 5692
rect 157567 5661 157579 5664
rect 157521 5655 157579 5661
rect 157889 5661 157901 5664
rect 157935 5692 157947 5695
rect 158625 5695 158683 5701
rect 158625 5692 158637 5695
rect 157935 5664 158637 5692
rect 157935 5661 157947 5664
rect 157889 5655 157947 5661
rect 158625 5661 158637 5664
rect 158671 5692 158683 5695
rect 158993 5695 159051 5701
rect 158993 5692 159005 5695
rect 158671 5664 159005 5692
rect 158671 5661 158683 5664
rect 158625 5655 158683 5661
rect 158993 5661 159005 5664
rect 159039 5692 159051 5695
rect 159361 5695 159419 5701
rect 159361 5692 159373 5695
rect 159039 5664 159373 5692
rect 159039 5661 159051 5664
rect 158993 5655 159051 5661
rect 159361 5661 159373 5664
rect 159407 5692 159419 5695
rect 160646 5692 160652 5704
rect 159407 5664 160652 5692
rect 159407 5661 159419 5664
rect 159361 5655 159419 5661
rect 160646 5652 160652 5664
rect 160704 5652 160710 5704
rect 161032 5692 161060 5800
rect 161290 5720 161296 5772
rect 161348 5760 161354 5772
rect 161348 5732 180748 5760
rect 161348 5720 161354 5732
rect 161109 5695 161167 5701
rect 161109 5692 161121 5695
rect 161032 5664 161121 5692
rect 161109 5661 161121 5664
rect 161155 5661 161167 5695
rect 161109 5655 161167 5661
rect 161201 5695 161259 5701
rect 161201 5661 161213 5695
rect 161247 5692 161259 5695
rect 161753 5695 161811 5701
rect 161753 5692 161765 5695
rect 161247 5664 161765 5692
rect 161247 5661 161259 5664
rect 161201 5655 161259 5661
rect 161753 5661 161765 5664
rect 161799 5661 161811 5695
rect 180613 5695 180671 5701
rect 180613 5692 180625 5695
rect 161753 5655 161811 5661
rect 161860 5664 171134 5692
rect 153286 5584 153292 5636
rect 153344 5624 153350 5636
rect 153565 5627 153623 5633
rect 153565 5624 153577 5627
rect 153344 5596 153577 5624
rect 153344 5584 153350 5596
rect 153565 5593 153577 5596
rect 153611 5624 153623 5627
rect 155862 5624 155868 5636
rect 153611 5596 155868 5624
rect 153611 5593 153623 5596
rect 153565 5587 153623 5593
rect 155862 5584 155868 5596
rect 155920 5584 155926 5636
rect 161860 5624 161888 5664
rect 157306 5596 161888 5624
rect 152369 5559 152427 5565
rect 152369 5556 152381 5559
rect 152056 5528 152381 5556
rect 152056 5516 152062 5528
rect 152369 5525 152381 5528
rect 152415 5556 152427 5559
rect 152737 5559 152795 5565
rect 152737 5556 152749 5559
rect 152415 5528 152749 5556
rect 152415 5525 152427 5528
rect 152369 5519 152427 5525
rect 152737 5525 152749 5528
rect 152783 5556 152795 5559
rect 157306 5556 157334 5596
rect 162026 5584 162032 5636
rect 162084 5624 162090 5636
rect 162121 5627 162179 5633
rect 162121 5624 162133 5627
rect 162084 5596 162133 5624
rect 162084 5584 162090 5596
rect 162121 5593 162133 5596
rect 162167 5593 162179 5627
rect 162121 5587 162179 5593
rect 162762 5584 162768 5636
rect 162820 5584 162826 5636
rect 152783 5528 157334 5556
rect 152783 5525 152795 5528
rect 152737 5519 152795 5525
rect 158070 5516 158076 5568
rect 158128 5556 158134 5568
rect 160189 5559 160247 5565
rect 160189 5556 160201 5559
rect 158128 5528 160201 5556
rect 158128 5516 158134 5528
rect 160189 5525 160201 5528
rect 160235 5556 160247 5559
rect 160554 5556 160560 5568
rect 160235 5528 160560 5556
rect 160235 5525 160247 5528
rect 160189 5519 160247 5525
rect 160554 5516 160560 5528
rect 160612 5516 160618 5568
rect 160646 5516 160652 5568
rect 160704 5556 160710 5568
rect 161290 5556 161296 5568
rect 160704 5528 161296 5556
rect 160704 5516 160710 5528
rect 161290 5516 161296 5528
rect 161348 5516 161354 5568
rect 162578 5516 162584 5568
rect 162636 5556 162642 5568
rect 162857 5559 162915 5565
rect 162857 5556 162869 5559
rect 162636 5528 162869 5556
rect 162636 5516 162642 5528
rect 162857 5525 162869 5528
rect 162903 5525 162915 5559
rect 171106 5556 171134 5664
rect 180536 5664 180625 5692
rect 177022 5556 177028 5568
rect 171106 5528 177028 5556
rect 162857 5519 162915 5525
rect 177022 5516 177028 5528
rect 177080 5516 177086 5568
rect 177942 5516 177948 5568
rect 178000 5556 178006 5568
rect 180337 5559 180395 5565
rect 180337 5556 180349 5559
rect 178000 5528 180349 5556
rect 178000 5516 178006 5528
rect 180337 5525 180349 5528
rect 180383 5556 180395 5559
rect 180536 5556 180564 5664
rect 180613 5661 180625 5664
rect 180659 5661 180671 5695
rect 180613 5655 180671 5661
rect 180720 5624 180748 5732
rect 180812 5701 180840 5800
rect 181806 5788 181812 5800
rect 181864 5788 181870 5840
rect 190426 5828 190454 5868
rect 216030 5856 216036 5868
rect 216088 5856 216094 5908
rect 217229 5899 217287 5905
rect 217229 5896 217241 5899
rect 216140 5868 217241 5896
rect 186286 5800 190454 5828
rect 182174 5760 182180 5772
rect 181640 5732 182180 5760
rect 181640 5701 181668 5732
rect 182174 5720 182180 5732
rect 182232 5720 182238 5772
rect 180797 5695 180855 5701
rect 180797 5661 180809 5695
rect 180843 5661 180855 5695
rect 180797 5655 180855 5661
rect 181625 5695 181683 5701
rect 181625 5661 181637 5695
rect 181671 5661 181683 5695
rect 181625 5655 181683 5661
rect 182082 5652 182088 5704
rect 182140 5652 182146 5704
rect 182361 5695 182419 5701
rect 182361 5661 182373 5695
rect 182407 5692 182419 5695
rect 182542 5692 182548 5704
rect 182407 5664 182548 5692
rect 182407 5661 182419 5664
rect 182361 5655 182419 5661
rect 182542 5652 182548 5664
rect 182600 5692 182606 5704
rect 186286 5692 186314 5800
rect 200758 5788 200764 5840
rect 200816 5828 200822 5840
rect 216140 5828 216168 5868
rect 217229 5865 217241 5868
rect 217275 5865 217287 5899
rect 217229 5859 217287 5865
rect 220998 5856 221004 5908
rect 221056 5896 221062 5908
rect 221093 5899 221151 5905
rect 221093 5896 221105 5899
rect 221056 5868 221105 5896
rect 221056 5856 221062 5868
rect 221093 5865 221105 5868
rect 221139 5896 221151 5899
rect 221461 5899 221519 5905
rect 221461 5896 221473 5899
rect 221139 5868 221473 5896
rect 221139 5865 221151 5868
rect 221093 5859 221151 5865
rect 221461 5865 221473 5868
rect 221507 5865 221519 5899
rect 221461 5859 221519 5865
rect 200816 5800 212212 5828
rect 200816 5788 200822 5800
rect 182600 5664 186314 5692
rect 190426 5732 195974 5760
rect 182600 5652 182606 5664
rect 190426 5624 190454 5732
rect 180720 5596 190454 5624
rect 186314 5556 186320 5568
rect 180383 5528 186320 5556
rect 180383 5525 180395 5528
rect 180337 5519 180395 5525
rect 186314 5516 186320 5528
rect 186372 5516 186378 5568
rect 195946 5556 195974 5732
rect 212184 5701 212212 5800
rect 212920 5800 216168 5828
rect 221476 5828 221504 5859
rect 223758 5856 223764 5908
rect 223816 5896 223822 5908
rect 224218 5896 224224 5908
rect 223816 5868 224224 5896
rect 223816 5856 223822 5868
rect 224218 5856 224224 5868
rect 224276 5856 224282 5908
rect 226150 5896 226156 5908
rect 224696 5868 226156 5896
rect 221476 5800 222332 5828
rect 212920 5776 212948 5800
rect 212828 5769 212948 5776
rect 212813 5763 212948 5769
rect 212813 5729 212825 5763
rect 212859 5748 212948 5763
rect 212859 5729 212871 5748
rect 212813 5723 212871 5729
rect 215386 5720 215392 5772
rect 215444 5720 215450 5772
rect 215938 5720 215944 5772
rect 215996 5760 216002 5772
rect 216033 5763 216091 5769
rect 216033 5760 216045 5763
rect 215996 5732 216045 5760
rect 215996 5720 216002 5732
rect 216033 5729 216045 5732
rect 216079 5729 216091 5763
rect 216033 5723 216091 5729
rect 216122 5720 216128 5772
rect 216180 5760 216186 5772
rect 216585 5763 216643 5769
rect 216585 5760 216597 5763
rect 216180 5732 216597 5760
rect 216180 5720 216186 5732
rect 216585 5729 216597 5732
rect 216631 5760 216643 5763
rect 218882 5760 218888 5772
rect 216631 5732 218888 5760
rect 216631 5729 216643 5732
rect 216585 5723 216643 5729
rect 218882 5720 218888 5732
rect 218940 5720 218946 5772
rect 221829 5763 221887 5769
rect 221829 5729 221841 5763
rect 221875 5760 221887 5763
rect 222010 5760 222016 5772
rect 221875 5732 222016 5760
rect 221875 5729 221887 5732
rect 221829 5723 221887 5729
rect 222010 5720 222016 5732
rect 222068 5720 222074 5772
rect 222304 5769 222332 5800
rect 223390 5788 223396 5840
rect 223448 5828 223454 5840
rect 224586 5828 224592 5840
rect 223448 5800 224592 5828
rect 223448 5788 223454 5800
rect 224586 5788 224592 5800
rect 224644 5788 224650 5840
rect 222289 5763 222347 5769
rect 222289 5729 222301 5763
rect 222335 5760 222347 5763
rect 223945 5763 224003 5769
rect 223945 5760 223957 5763
rect 222335 5732 223957 5760
rect 222335 5729 222347 5732
rect 222289 5723 222347 5729
rect 223945 5729 223957 5732
rect 223991 5760 224003 5763
rect 224313 5763 224371 5769
rect 224313 5760 224325 5763
rect 223991 5732 224325 5760
rect 223991 5729 224003 5732
rect 223945 5723 224003 5729
rect 224313 5729 224325 5732
rect 224359 5760 224371 5763
rect 224696 5760 224724 5868
rect 226150 5856 226156 5868
rect 226208 5856 226214 5908
rect 226242 5856 226248 5908
rect 226300 5896 226306 5908
rect 226300 5868 227116 5896
rect 226300 5856 226306 5868
rect 224957 5831 225015 5837
rect 224957 5797 224969 5831
rect 225003 5828 225015 5831
rect 227088 5828 227116 5868
rect 227622 5856 227628 5908
rect 227680 5896 227686 5908
rect 228453 5899 228511 5905
rect 228453 5896 228465 5899
rect 227680 5868 228465 5896
rect 227680 5856 227686 5868
rect 228453 5865 228465 5868
rect 228499 5865 228511 5899
rect 228453 5859 228511 5865
rect 228560 5868 229232 5896
rect 228560 5828 228588 5868
rect 225003 5800 226288 5828
rect 227088 5800 228588 5828
rect 228637 5831 228695 5837
rect 225003 5797 225015 5800
rect 224957 5791 225015 5797
rect 225509 5763 225567 5769
rect 225509 5760 225521 5763
rect 224359 5732 224724 5760
rect 224926 5732 225521 5760
rect 224359 5729 224371 5732
rect 224313 5723 224371 5729
rect 212169 5695 212227 5701
rect 212169 5661 212181 5695
rect 212215 5692 212227 5695
rect 212534 5692 212540 5704
rect 212215 5664 212540 5692
rect 212215 5661 212227 5664
rect 212169 5655 212227 5661
rect 212534 5652 212540 5664
rect 212592 5652 212598 5704
rect 214650 5652 214656 5704
rect 214708 5652 214714 5704
rect 215570 5652 215576 5704
rect 215628 5652 215634 5704
rect 216306 5652 216312 5704
rect 216364 5652 216370 5704
rect 216490 5701 216496 5704
rect 216447 5695 216496 5701
rect 216447 5661 216459 5695
rect 216493 5661 216496 5695
rect 216447 5655 216496 5661
rect 216490 5652 216496 5655
rect 216548 5652 216554 5704
rect 223574 5652 223580 5704
rect 223632 5692 223638 5704
rect 224926 5692 224954 5732
rect 225509 5729 225521 5732
rect 225555 5729 225567 5763
rect 225509 5723 225567 5729
rect 226058 5720 226064 5772
rect 226116 5760 226122 5772
rect 226153 5763 226211 5769
rect 226153 5760 226165 5763
rect 226116 5732 226165 5760
rect 226116 5720 226122 5732
rect 226153 5729 226165 5732
rect 226199 5729 226211 5763
rect 226260 5760 226288 5800
rect 228637 5797 228649 5831
rect 228683 5828 228695 5831
rect 229204 5828 229232 5868
rect 229554 5856 229560 5908
rect 229612 5896 229618 5908
rect 230845 5899 230903 5905
rect 230845 5896 230857 5899
rect 229612 5868 230857 5896
rect 229612 5856 229618 5868
rect 230845 5865 230857 5868
rect 230891 5865 230903 5899
rect 230845 5859 230903 5865
rect 231029 5899 231087 5905
rect 231029 5865 231041 5899
rect 231075 5896 231087 5899
rect 231302 5896 231308 5908
rect 231075 5868 231308 5896
rect 231075 5865 231087 5868
rect 231029 5859 231087 5865
rect 231302 5856 231308 5868
rect 231360 5856 231366 5908
rect 231394 5856 231400 5908
rect 231452 5896 231458 5908
rect 232501 5899 232559 5905
rect 232501 5896 232513 5899
rect 231452 5868 232513 5896
rect 231452 5856 231458 5868
rect 232501 5865 232513 5868
rect 232547 5865 232559 5899
rect 232501 5859 232559 5865
rect 258350 5856 258356 5908
rect 258408 5896 258414 5908
rect 261110 5896 261116 5908
rect 258408 5868 261116 5896
rect 258408 5856 258414 5868
rect 261110 5856 261116 5868
rect 261168 5856 261174 5908
rect 261202 5856 261208 5908
rect 261260 5896 261266 5908
rect 265529 5899 265587 5905
rect 265529 5896 265541 5899
rect 261260 5868 265541 5896
rect 261260 5856 261266 5868
rect 265529 5865 265541 5868
rect 265575 5865 265587 5899
rect 270494 5896 270500 5908
rect 265529 5859 265587 5865
rect 267016 5868 270500 5896
rect 244182 5828 244188 5840
rect 228683 5800 229140 5828
rect 229204 5800 244188 5828
rect 228683 5797 228695 5800
rect 228637 5791 228695 5797
rect 229112 5769 229140 5800
rect 244182 5788 244188 5800
rect 244240 5788 244246 5840
rect 258810 5788 258816 5840
rect 258868 5828 258874 5840
rect 260098 5828 260104 5840
rect 258868 5800 260104 5828
rect 258868 5788 258874 5800
rect 260098 5788 260104 5800
rect 260156 5788 260162 5840
rect 262674 5788 262680 5840
rect 262732 5828 262738 5840
rect 267016 5828 267044 5868
rect 270494 5856 270500 5868
rect 270552 5856 270558 5908
rect 262732 5800 267044 5828
rect 262732 5788 262738 5800
rect 267734 5788 267740 5840
rect 267792 5828 267798 5840
rect 270681 5831 270739 5837
rect 270681 5828 270693 5831
rect 267792 5800 270693 5828
rect 267792 5788 267798 5800
rect 270681 5797 270693 5800
rect 270727 5797 270739 5831
rect 270681 5791 270739 5797
rect 226429 5763 226487 5769
rect 226429 5760 226441 5763
rect 226260 5732 226441 5760
rect 226153 5723 226211 5729
rect 226429 5729 226441 5732
rect 226475 5760 226487 5763
rect 229097 5763 229155 5769
rect 226475 5732 228680 5760
rect 226475 5729 226487 5732
rect 226429 5723 226487 5729
rect 223632 5664 224954 5692
rect 223632 5652 223638 5664
rect 225046 5652 225052 5704
rect 225104 5692 225110 5704
rect 225693 5695 225751 5701
rect 225693 5692 225705 5695
rect 225104 5664 225705 5692
rect 225104 5652 225110 5664
rect 225693 5661 225705 5664
rect 225739 5661 225751 5695
rect 225693 5655 225751 5661
rect 226518 5652 226524 5704
rect 226576 5701 226582 5704
rect 226576 5695 226604 5701
rect 226592 5661 226604 5695
rect 226576 5655 226604 5661
rect 226576 5652 226582 5655
rect 226702 5652 226708 5704
rect 226760 5652 226766 5704
rect 227714 5652 227720 5704
rect 227772 5652 227778 5704
rect 228082 5652 228088 5704
rect 228140 5652 228146 5704
rect 209958 5584 209964 5636
rect 210016 5624 210022 5636
rect 212994 5624 213000 5636
rect 210016 5596 213000 5624
rect 210016 5584 210022 5596
rect 212994 5584 213000 5596
rect 213052 5584 213058 5636
rect 215478 5624 215484 5636
rect 213104 5596 215484 5624
rect 213104 5556 213132 5596
rect 215478 5584 215484 5596
rect 215536 5584 215542 5636
rect 217134 5584 217140 5636
rect 217192 5624 217198 5636
rect 219250 5624 219256 5636
rect 217192 5596 219256 5624
rect 217192 5584 217198 5596
rect 219250 5584 219256 5596
rect 219308 5584 219314 5636
rect 222010 5584 222016 5636
rect 222068 5584 222074 5636
rect 222286 5584 222292 5636
rect 222344 5624 222350 5636
rect 222838 5624 222844 5636
rect 222344 5596 222844 5624
rect 222344 5584 222350 5596
rect 222838 5584 222844 5596
rect 222896 5584 222902 5636
rect 223298 5584 223304 5636
rect 223356 5624 223362 5636
rect 224862 5624 224868 5636
rect 223356 5596 224868 5624
rect 223356 5584 223362 5596
rect 224862 5584 224868 5596
rect 224920 5584 224926 5636
rect 228450 5624 228456 5636
rect 227180 5596 228456 5624
rect 195946 5528 213132 5556
rect 214650 5516 214656 5568
rect 214708 5556 214714 5568
rect 215297 5559 215355 5565
rect 215297 5556 215309 5559
rect 214708 5528 215309 5556
rect 214708 5516 214714 5528
rect 215297 5525 215309 5528
rect 215343 5556 215355 5559
rect 215938 5556 215944 5568
rect 215343 5528 215944 5556
rect 215343 5525 215355 5528
rect 215297 5519 215355 5525
rect 215938 5516 215944 5528
rect 215996 5516 216002 5568
rect 216030 5516 216036 5568
rect 216088 5556 216094 5568
rect 227180 5556 227208 5596
rect 228450 5584 228456 5596
rect 228508 5584 228514 5636
rect 216088 5528 227208 5556
rect 216088 5516 216094 5528
rect 227346 5516 227352 5568
rect 227404 5516 227410 5568
rect 228652 5556 228680 5732
rect 229097 5729 229109 5763
rect 229143 5729 229155 5763
rect 231210 5760 231216 5772
rect 229097 5723 229155 5729
rect 230032 5732 231216 5760
rect 230032 5704 230060 5732
rect 231210 5720 231216 5732
rect 231268 5760 231274 5772
rect 231268 5732 231716 5760
rect 231268 5720 231274 5732
rect 229373 5695 229431 5701
rect 229373 5661 229385 5695
rect 229419 5692 229431 5695
rect 230014 5692 230020 5704
rect 229419 5664 230020 5692
rect 229419 5661 229431 5664
rect 229373 5655 229431 5661
rect 230014 5652 230020 5664
rect 230072 5652 230078 5704
rect 231486 5652 231492 5704
rect 231544 5652 231550 5704
rect 231688 5701 231716 5732
rect 231854 5720 231860 5772
rect 231912 5760 231918 5772
rect 259270 5760 259276 5772
rect 231912 5732 259276 5760
rect 231912 5720 231918 5732
rect 259270 5720 259276 5732
rect 259328 5720 259334 5772
rect 231673 5695 231731 5701
rect 231673 5661 231685 5695
rect 231719 5661 231731 5695
rect 231673 5655 231731 5661
rect 232314 5652 232320 5704
rect 232372 5652 232378 5704
rect 256878 5692 256884 5704
rect 234586 5664 256884 5692
rect 228910 5584 228916 5636
rect 228968 5624 228974 5636
rect 229830 5624 229836 5636
rect 228968 5596 229836 5624
rect 228968 5584 228974 5596
rect 229830 5584 229836 5596
rect 229888 5584 229894 5636
rect 229922 5584 229928 5636
rect 229980 5624 229986 5636
rect 230658 5624 230664 5636
rect 229980 5596 230664 5624
rect 229980 5584 229986 5596
rect 230658 5584 230664 5596
rect 230716 5584 230722 5636
rect 230842 5584 230848 5636
rect 230900 5633 230906 5636
rect 230900 5627 230919 5633
rect 230907 5624 230919 5627
rect 231857 5627 231915 5633
rect 231857 5624 231869 5627
rect 230907 5596 231869 5624
rect 230907 5593 230919 5596
rect 230900 5587 230919 5593
rect 231857 5593 231869 5596
rect 231903 5593 231915 5627
rect 231857 5587 231915 5593
rect 230900 5584 230906 5587
rect 234586 5556 234614 5664
rect 256878 5652 256884 5664
rect 256936 5652 256942 5704
rect 258997 5695 259055 5701
rect 258997 5661 259009 5695
rect 259043 5692 259055 5695
rect 259043 5664 260052 5692
rect 259043 5661 259055 5664
rect 258997 5655 259055 5661
rect 237374 5584 237380 5636
rect 237432 5624 237438 5636
rect 259086 5624 259092 5636
rect 237432 5596 259092 5624
rect 237432 5584 237438 5596
rect 259086 5584 259092 5596
rect 259144 5624 259150 5636
rect 259365 5627 259423 5633
rect 259365 5624 259377 5627
rect 259144 5596 259377 5624
rect 259144 5584 259150 5596
rect 259365 5593 259377 5596
rect 259411 5593 259423 5627
rect 259365 5587 259423 5593
rect 228652 5528 234614 5556
rect 252278 5516 252284 5568
rect 252336 5556 252342 5568
rect 258810 5556 258816 5568
rect 252336 5528 258816 5556
rect 252336 5516 252342 5528
rect 258810 5516 258816 5528
rect 258868 5516 258874 5568
rect 260024 5556 260052 5664
rect 260116 5624 260144 5788
rect 262214 5760 262220 5772
rect 260208 5732 262220 5760
rect 260208 5701 260236 5732
rect 262214 5720 262220 5732
rect 262272 5720 262278 5772
rect 263134 5720 263140 5772
rect 263192 5720 263198 5772
rect 266722 5760 266728 5772
rect 263980 5732 266728 5760
rect 260193 5695 260251 5701
rect 260193 5661 260205 5695
rect 260239 5661 260251 5695
rect 260193 5655 260251 5661
rect 261662 5652 261668 5704
rect 261720 5652 261726 5704
rect 262861 5695 262919 5701
rect 262861 5661 262873 5695
rect 262907 5692 262919 5695
rect 263980 5692 264008 5732
rect 266722 5720 266728 5732
rect 266780 5720 266786 5772
rect 269853 5763 269911 5769
rect 269853 5760 269865 5763
rect 267108 5732 269865 5760
rect 262907 5664 264008 5692
rect 262907 5661 262919 5664
rect 262861 5655 262919 5661
rect 264054 5652 264060 5704
rect 264112 5652 264118 5704
rect 264514 5652 264520 5704
rect 264572 5652 264578 5704
rect 265250 5652 265256 5704
rect 265308 5652 265314 5704
rect 265345 5695 265403 5701
rect 265345 5661 265357 5695
rect 265391 5661 265403 5695
rect 265345 5655 265403 5661
rect 265989 5695 266047 5701
rect 265989 5661 266001 5695
rect 266035 5692 266047 5695
rect 266817 5695 266875 5701
rect 266035 5664 266768 5692
rect 266035 5661 266047 5664
rect 265989 5655 266047 5661
rect 260561 5627 260619 5633
rect 260561 5624 260573 5627
rect 260116 5596 260573 5624
rect 260561 5593 260573 5596
rect 260607 5593 260619 5627
rect 260561 5587 260619 5593
rect 261110 5584 261116 5636
rect 261168 5624 261174 5636
rect 262033 5627 262091 5633
rect 262033 5624 262045 5627
rect 261168 5596 262045 5624
rect 261168 5584 261174 5596
rect 262033 5593 262045 5596
rect 262079 5593 262091 5627
rect 262033 5587 262091 5593
rect 263134 5584 263140 5636
rect 263192 5624 263198 5636
rect 263594 5624 263600 5636
rect 263192 5596 263600 5624
rect 263192 5584 263198 5596
rect 263594 5584 263600 5596
rect 263652 5584 263658 5636
rect 264882 5584 264888 5636
rect 264940 5624 264946 5636
rect 265360 5624 265388 5655
rect 265894 5624 265900 5636
rect 264940 5596 265900 5624
rect 264940 5584 264946 5596
rect 265894 5584 265900 5596
rect 265952 5624 265958 5636
rect 266170 5624 266176 5636
rect 265952 5596 266176 5624
rect 265952 5584 265958 5596
rect 266170 5584 266176 5596
rect 266228 5584 266234 5636
rect 266740 5624 266768 5664
rect 266817 5661 266829 5695
rect 266863 5692 266875 5695
rect 267108 5692 267136 5732
rect 269853 5729 269865 5732
rect 269899 5729 269911 5763
rect 269853 5723 269911 5729
rect 266863 5664 267136 5692
rect 266863 5661 266875 5664
rect 266817 5655 266875 5661
rect 267182 5652 267188 5704
rect 267240 5652 267246 5704
rect 268381 5695 268439 5701
rect 268381 5661 268393 5695
rect 268427 5692 268439 5695
rect 269022 5692 269028 5704
rect 268427 5664 269028 5692
rect 268427 5661 268439 5664
rect 268381 5655 268439 5661
rect 269022 5652 269028 5664
rect 269080 5652 269086 5704
rect 269482 5652 269488 5704
rect 269540 5652 269546 5704
rect 269669 5695 269727 5701
rect 269669 5661 269681 5695
rect 269715 5661 269727 5695
rect 269669 5655 269727 5661
rect 270313 5695 270371 5701
rect 270313 5661 270325 5695
rect 270359 5661 270371 5695
rect 270313 5655 270371 5661
rect 268654 5624 268660 5636
rect 266740 5596 268660 5624
rect 268654 5584 268660 5596
rect 268712 5584 268718 5636
rect 268838 5584 268844 5636
rect 268896 5584 268902 5636
rect 269206 5584 269212 5636
rect 269264 5624 269270 5636
rect 269684 5624 269712 5655
rect 269264 5596 269712 5624
rect 269264 5584 269270 5596
rect 261938 5556 261944 5568
rect 260024 5528 261944 5556
rect 261938 5516 261944 5528
rect 261996 5516 262002 5568
rect 266354 5516 266360 5568
rect 266412 5556 266418 5568
rect 270328 5556 270356 5655
rect 270402 5652 270408 5704
rect 270460 5692 270466 5704
rect 270497 5695 270555 5701
rect 270497 5692 270509 5695
rect 270460 5664 270509 5692
rect 270460 5652 270466 5664
rect 270497 5661 270509 5664
rect 270543 5661 270555 5695
rect 270497 5655 270555 5661
rect 266412 5528 270356 5556
rect 266412 5516 266418 5528
rect 1104 5466 271651 5488
rect 1104 5414 68546 5466
rect 68598 5414 68610 5466
rect 68662 5414 68674 5466
rect 68726 5414 68738 5466
rect 68790 5414 68802 5466
rect 68854 5414 136143 5466
rect 136195 5414 136207 5466
rect 136259 5414 136271 5466
rect 136323 5414 136335 5466
rect 136387 5414 136399 5466
rect 136451 5414 203740 5466
rect 203792 5414 203804 5466
rect 203856 5414 203868 5466
rect 203920 5414 203932 5466
rect 203984 5414 203996 5466
rect 204048 5414 271337 5466
rect 271389 5414 271401 5466
rect 271453 5414 271465 5466
rect 271517 5414 271529 5466
rect 271581 5414 271593 5466
rect 271645 5414 271651 5466
rect 1104 5392 271651 5414
rect 15286 5312 15292 5364
rect 15344 5352 15350 5364
rect 34606 5352 34612 5364
rect 15344 5324 34612 5352
rect 15344 5312 15350 5324
rect 34606 5312 34612 5324
rect 34664 5312 34670 5364
rect 35084 5324 38424 5352
rect 26878 5244 26884 5296
rect 26936 5284 26942 5296
rect 35084 5284 35112 5324
rect 26936 5256 35112 5284
rect 37645 5287 37703 5293
rect 26936 5244 26942 5256
rect 37645 5253 37657 5287
rect 37691 5284 37703 5287
rect 37826 5284 37832 5296
rect 37691 5256 37832 5284
rect 37691 5253 37703 5256
rect 37645 5247 37703 5253
rect 37826 5244 37832 5256
rect 37884 5244 37890 5296
rect 37918 5244 37924 5296
rect 37976 5244 37982 5296
rect 38396 5293 38424 5324
rect 43530 5312 43536 5364
rect 43588 5312 43594 5364
rect 45370 5312 45376 5364
rect 45428 5352 45434 5364
rect 46842 5352 46848 5364
rect 45428 5324 46848 5352
rect 45428 5312 45434 5324
rect 38381 5287 38439 5293
rect 38381 5253 38393 5287
rect 38427 5253 38439 5287
rect 38381 5247 38439 5253
rect 38746 5244 38752 5296
rect 38804 5244 38810 5296
rect 43346 5244 43352 5296
rect 43404 5244 43410 5296
rect 43548 5284 43576 5312
rect 43625 5287 43683 5293
rect 43625 5284 43637 5287
rect 43548 5256 43637 5284
rect 43625 5253 43637 5256
rect 43671 5253 43683 5287
rect 43625 5247 43683 5253
rect 43714 5244 43720 5296
rect 43772 5244 43778 5296
rect 44358 5244 44364 5296
rect 44416 5284 44422 5296
rect 44453 5287 44511 5293
rect 44453 5284 44465 5287
rect 44416 5256 44465 5284
rect 44416 5244 44422 5256
rect 44453 5253 44465 5256
rect 44499 5253 44511 5287
rect 44453 5247 44511 5253
rect 45830 5244 45836 5296
rect 45888 5244 45894 5296
rect 46106 5244 46112 5296
rect 46164 5244 46170 5296
rect 46216 5293 46244 5324
rect 46842 5312 46848 5324
rect 46900 5312 46906 5364
rect 47121 5355 47179 5361
rect 47121 5321 47133 5355
rect 47167 5352 47179 5355
rect 47167 5324 52040 5352
rect 47167 5321 47179 5324
rect 47121 5315 47179 5321
rect 46201 5287 46259 5293
rect 46201 5253 46213 5287
rect 46247 5253 46259 5287
rect 46201 5247 46259 5253
rect 46290 5244 46296 5296
rect 46348 5284 46354 5296
rect 46937 5287 46995 5293
rect 46937 5284 46949 5287
rect 46348 5256 46949 5284
rect 46348 5244 46354 5256
rect 46937 5253 46949 5256
rect 46983 5253 46995 5287
rect 50617 5287 50675 5293
rect 46937 5247 46995 5253
rect 49344 5256 50568 5284
rect 49344 5228 49372 5256
rect 38013 5219 38071 5225
rect 38013 5185 38025 5219
rect 38059 5216 38071 5219
rect 38194 5216 38200 5228
rect 38059 5188 38200 5216
rect 38059 5185 38071 5188
rect 38013 5179 38071 5185
rect 38194 5176 38200 5188
rect 38252 5176 38258 5228
rect 41601 5219 41659 5225
rect 41601 5185 41613 5219
rect 41647 5216 41659 5219
rect 42610 5216 42616 5228
rect 41647 5188 42616 5216
rect 41647 5185 41659 5188
rect 41601 5179 41659 5185
rect 42610 5176 42616 5188
rect 42668 5176 42674 5228
rect 43806 5176 43812 5228
rect 43864 5216 43870 5228
rect 44085 5219 44143 5225
rect 44085 5216 44097 5219
rect 43864 5188 44097 5216
rect 43864 5176 43870 5188
rect 44085 5185 44097 5188
rect 44131 5185 44143 5219
rect 44085 5179 44143 5185
rect 45922 5176 45928 5228
rect 45980 5216 45986 5228
rect 46569 5219 46627 5225
rect 46569 5216 46581 5219
rect 45980 5188 46581 5216
rect 45980 5176 45986 5188
rect 46569 5185 46581 5188
rect 46615 5185 46627 5219
rect 46569 5179 46627 5185
rect 47946 5176 47952 5228
rect 48004 5216 48010 5228
rect 49326 5216 49332 5228
rect 48004 5188 49332 5216
rect 48004 5176 48010 5188
rect 49326 5176 49332 5188
rect 49384 5176 49390 5228
rect 50540 5216 50568 5256
rect 50617 5253 50629 5287
rect 50663 5284 50675 5287
rect 50706 5284 50712 5296
rect 50663 5256 50712 5284
rect 50663 5253 50675 5256
rect 50617 5247 50675 5253
rect 50706 5244 50712 5256
rect 50764 5244 50770 5296
rect 50893 5287 50951 5293
rect 50893 5253 50905 5287
rect 50939 5284 50951 5287
rect 51166 5284 51172 5296
rect 50939 5256 51172 5284
rect 50939 5253 50951 5256
rect 50893 5247 50951 5253
rect 51166 5244 51172 5256
rect 51224 5244 51230 5296
rect 51350 5244 51356 5296
rect 51408 5244 51414 5296
rect 51442 5244 51448 5296
rect 51500 5284 51506 5296
rect 51721 5287 51779 5293
rect 51721 5284 51733 5287
rect 51500 5256 51733 5284
rect 51500 5244 51506 5256
rect 51721 5253 51733 5256
rect 51767 5253 51779 5287
rect 51721 5247 51779 5253
rect 50982 5216 50988 5228
rect 50540 5188 50988 5216
rect 50982 5176 50988 5188
rect 51040 5176 51046 5228
rect 51632 5160 51684 5166
rect 38470 5108 38476 5160
rect 38528 5108 38534 5160
rect 40770 5108 40776 5160
rect 40828 5148 40834 5160
rect 41138 5148 41144 5160
rect 40828 5120 41144 5148
rect 40828 5108 40834 5120
rect 41138 5108 41144 5120
rect 41196 5148 41202 5160
rect 41785 5151 41843 5157
rect 41785 5148 41797 5151
rect 41196 5120 41797 5148
rect 41196 5108 41202 5120
rect 41785 5117 41797 5120
rect 41831 5117 41843 5151
rect 41785 5111 41843 5117
rect 42426 5108 42432 5160
rect 42484 5148 42490 5160
rect 42705 5151 42763 5157
rect 42705 5148 42717 5151
rect 42484 5120 42717 5148
rect 42484 5108 42490 5120
rect 42705 5117 42717 5120
rect 42751 5117 42763 5151
rect 44726 5148 44732 5160
rect 44390 5120 44732 5148
rect 42705 5111 42763 5117
rect 44726 5108 44732 5120
rect 44784 5108 44790 5160
rect 48038 5148 48044 5160
rect 46874 5120 48044 5148
rect 48038 5108 48044 5120
rect 48096 5108 48102 5160
rect 51632 5102 51684 5108
rect 38933 5083 38991 5089
rect 38933 5049 38945 5083
rect 38979 5080 38991 5083
rect 42886 5080 42892 5092
rect 38979 5052 42892 5080
rect 38979 5049 38991 5052
rect 38933 5043 38991 5049
rect 42886 5040 42892 5052
rect 42944 5040 42950 5092
rect 44634 5040 44640 5092
rect 44692 5040 44698 5092
rect 52012 5080 52040 5324
rect 53098 5312 53104 5364
rect 53156 5312 53162 5364
rect 101125 5355 101183 5361
rect 60706 5324 81480 5352
rect 52086 5244 52092 5296
rect 52144 5284 52150 5296
rect 60706 5284 60734 5324
rect 52144 5256 60734 5284
rect 52144 5244 52150 5256
rect 80330 5244 80336 5296
rect 80388 5244 80394 5296
rect 80701 5287 80759 5293
rect 80701 5253 80713 5287
rect 80747 5284 80759 5287
rect 81342 5284 81348 5296
rect 80747 5256 81348 5284
rect 80747 5253 80759 5256
rect 80701 5247 80759 5253
rect 81342 5244 81348 5256
rect 81400 5244 81406 5296
rect 53009 5219 53067 5225
rect 53009 5185 53021 5219
rect 53055 5185 53067 5219
rect 53009 5179 53067 5185
rect 53024 5148 53052 5179
rect 80790 5176 80796 5228
rect 80848 5176 80854 5228
rect 80882 5176 80888 5228
rect 80940 5176 80946 5228
rect 81452 5225 81480 5324
rect 82832 5324 99374 5352
rect 81618 5244 81624 5296
rect 81676 5244 81682 5296
rect 81437 5219 81495 5225
rect 81437 5185 81449 5219
rect 81483 5185 81495 5219
rect 81437 5179 81495 5185
rect 53745 5151 53803 5157
rect 53745 5148 53757 5151
rect 53024 5120 53757 5148
rect 53745 5117 53757 5120
rect 53791 5148 53803 5151
rect 79781 5151 79839 5157
rect 79781 5148 79793 5151
rect 53791 5120 79793 5148
rect 53791 5117 53803 5120
rect 53745 5111 53803 5117
rect 79781 5117 79793 5120
rect 79827 5148 79839 5151
rect 80149 5151 80207 5157
rect 80149 5148 80161 5151
rect 79827 5120 80161 5148
rect 79827 5117 79839 5120
rect 79781 5111 79839 5117
rect 80149 5117 80161 5120
rect 80195 5148 80207 5151
rect 82832 5148 82860 5324
rect 82906 5244 82912 5296
rect 82964 5284 82970 5296
rect 84746 5284 84752 5296
rect 82964 5256 84752 5284
rect 82964 5244 82970 5256
rect 84746 5244 84752 5256
rect 84804 5244 84810 5296
rect 84930 5244 84936 5296
rect 84988 5244 84994 5296
rect 86586 5244 86592 5296
rect 86644 5244 86650 5296
rect 87693 5287 87751 5293
rect 87693 5253 87705 5287
rect 87739 5284 87751 5287
rect 88061 5287 88119 5293
rect 88061 5284 88073 5287
rect 87739 5256 88073 5284
rect 87739 5253 87751 5256
rect 87693 5247 87751 5253
rect 88061 5253 88073 5256
rect 88107 5284 88119 5287
rect 88429 5287 88487 5293
rect 88429 5284 88441 5287
rect 88107 5256 88441 5284
rect 88107 5253 88119 5256
rect 88061 5247 88119 5253
rect 88429 5253 88441 5256
rect 88475 5284 88487 5287
rect 89165 5287 89223 5293
rect 89165 5284 89177 5287
rect 88475 5256 89177 5284
rect 88475 5253 88487 5256
rect 88429 5247 88487 5253
rect 89165 5253 89177 5256
rect 89211 5284 89223 5287
rect 91281 5287 91339 5293
rect 91281 5284 91293 5287
rect 89211 5256 91293 5284
rect 89211 5253 89223 5256
rect 89165 5247 89223 5253
rect 91281 5253 91293 5256
rect 91327 5284 91339 5287
rect 91649 5287 91707 5293
rect 91649 5284 91661 5287
rect 91327 5256 91661 5284
rect 91327 5253 91339 5256
rect 91281 5247 91339 5253
rect 91649 5253 91661 5256
rect 91695 5284 91707 5287
rect 93854 5284 93860 5296
rect 91695 5256 93860 5284
rect 91695 5253 91707 5256
rect 91649 5247 91707 5253
rect 93854 5244 93860 5256
rect 93912 5244 93918 5296
rect 99346 5284 99374 5324
rect 101125 5321 101137 5355
rect 101171 5352 101183 5355
rect 101306 5352 101312 5364
rect 101171 5324 101312 5352
rect 101171 5321 101183 5324
rect 101125 5315 101183 5321
rect 101306 5312 101312 5324
rect 101364 5312 101370 5364
rect 108758 5352 108764 5364
rect 101416 5324 108764 5352
rect 101416 5284 101444 5324
rect 108758 5312 108764 5324
rect 108816 5312 108822 5364
rect 110690 5312 110696 5364
rect 110748 5352 110754 5364
rect 115014 5352 115020 5364
rect 110748 5324 115020 5352
rect 110748 5312 110754 5324
rect 115014 5312 115020 5324
rect 115072 5312 115078 5364
rect 119249 5355 119307 5361
rect 119249 5321 119261 5355
rect 119295 5352 119307 5355
rect 120074 5352 120080 5364
rect 119295 5324 120080 5352
rect 119295 5321 119307 5324
rect 119249 5315 119307 5321
rect 120074 5312 120080 5324
rect 120132 5312 120138 5364
rect 142798 5312 142804 5364
rect 142856 5352 142862 5364
rect 152366 5352 152372 5364
rect 142856 5324 152372 5352
rect 142856 5312 142862 5324
rect 152366 5312 152372 5324
rect 152424 5312 152430 5364
rect 152461 5355 152519 5361
rect 152461 5321 152473 5355
rect 152507 5352 152519 5355
rect 153378 5352 153384 5364
rect 152507 5324 153384 5352
rect 152507 5321 152519 5324
rect 152461 5315 152519 5321
rect 153378 5312 153384 5324
rect 153436 5312 153442 5364
rect 157794 5352 157800 5364
rect 157306 5324 157800 5352
rect 99346 5256 101444 5284
rect 114370 5244 114376 5296
rect 114428 5284 114434 5296
rect 115293 5287 115351 5293
rect 115293 5284 115305 5287
rect 114428 5256 115305 5284
rect 114428 5244 114434 5256
rect 115293 5253 115305 5256
rect 115339 5284 115351 5287
rect 116302 5284 116308 5296
rect 115339 5256 116308 5284
rect 115339 5253 115351 5256
rect 115293 5247 115351 5253
rect 116302 5244 116308 5256
rect 116360 5244 116366 5296
rect 120258 5284 120264 5296
rect 120092 5256 120264 5284
rect 100938 5176 100944 5228
rect 100996 5216 101002 5228
rect 101033 5219 101091 5225
rect 101033 5216 101045 5219
rect 100996 5188 101045 5216
rect 100996 5176 101002 5188
rect 101033 5185 101045 5188
rect 101079 5185 101091 5219
rect 101033 5179 101091 5185
rect 106108 5188 106412 5216
rect 80195 5120 82860 5148
rect 83277 5151 83335 5157
rect 80195 5117 80207 5120
rect 80149 5111 80207 5117
rect 83277 5117 83289 5151
rect 83323 5148 83335 5151
rect 83829 5151 83887 5157
rect 83829 5148 83841 5151
rect 83323 5120 83841 5148
rect 83323 5117 83335 5120
rect 83277 5111 83335 5117
rect 83829 5117 83841 5120
rect 83875 5148 83887 5151
rect 84654 5148 84660 5160
rect 83875 5120 84660 5148
rect 83875 5117 83887 5120
rect 83829 5111 83887 5117
rect 84654 5108 84660 5120
rect 84712 5108 84718 5160
rect 84746 5108 84752 5160
rect 84804 5108 84810 5160
rect 89441 5151 89499 5157
rect 89441 5117 89453 5151
rect 89487 5117 89499 5151
rect 89441 5111 89499 5117
rect 89625 5151 89683 5157
rect 89625 5117 89637 5151
rect 89671 5117 89683 5151
rect 89625 5111 89683 5117
rect 89456 5080 89484 5111
rect 52012 5052 89484 5080
rect 89530 5040 89536 5092
rect 89588 5080 89594 5092
rect 89640 5080 89668 5111
rect 91738 5108 91744 5160
rect 91796 5108 91802 5160
rect 91922 5108 91928 5160
rect 91980 5148 91986 5160
rect 92658 5148 92664 5160
rect 91980 5120 92664 5148
rect 91980 5108 91986 5120
rect 92658 5108 92664 5120
rect 92716 5108 92722 5160
rect 93581 5151 93639 5157
rect 93581 5117 93593 5151
rect 93627 5148 93639 5151
rect 93627 5120 94268 5148
rect 93627 5117 93639 5120
rect 93581 5111 93639 5117
rect 94240 5089 94268 5120
rect 100662 5108 100668 5160
rect 100720 5148 100726 5160
rect 106108 5157 106136 5188
rect 106093 5151 106151 5157
rect 106093 5148 106105 5151
rect 100720 5120 106105 5148
rect 100720 5108 100726 5120
rect 106093 5117 106105 5120
rect 106139 5117 106151 5151
rect 106093 5111 106151 5117
rect 106277 5151 106335 5157
rect 106277 5117 106289 5151
rect 106323 5117 106335 5151
rect 106384 5148 106412 5188
rect 107010 5176 107016 5228
rect 107068 5176 107074 5228
rect 107194 5225 107200 5228
rect 107151 5219 107200 5225
rect 107151 5185 107163 5219
rect 107197 5185 107200 5219
rect 107151 5179 107200 5185
rect 107194 5176 107200 5179
rect 107252 5176 107258 5228
rect 107286 5176 107292 5228
rect 107344 5176 107350 5228
rect 117406 5176 117412 5228
rect 117464 5176 117470 5228
rect 120092 5225 120120 5256
rect 120258 5244 120264 5256
rect 120316 5244 120322 5296
rect 150253 5287 150311 5293
rect 150253 5253 150265 5287
rect 150299 5284 150311 5287
rect 150526 5284 150532 5296
rect 150299 5256 150532 5284
rect 150299 5253 150311 5256
rect 150253 5247 150311 5253
rect 150526 5244 150532 5256
rect 150584 5244 150590 5296
rect 153286 5244 153292 5296
rect 153344 5244 153350 5296
rect 120077 5219 120135 5225
rect 120077 5185 120089 5219
rect 120123 5185 120135 5219
rect 120077 5179 120135 5185
rect 120994 5176 121000 5228
rect 121052 5176 121058 5228
rect 122190 5176 122196 5228
rect 122248 5176 122254 5228
rect 123478 5176 123484 5228
rect 123536 5216 123542 5228
rect 123536 5188 138014 5216
rect 123536 5176 123542 5188
rect 108209 5151 108267 5157
rect 108209 5148 108221 5151
rect 106384 5120 108221 5148
rect 106277 5111 106335 5117
rect 108209 5117 108221 5120
rect 108255 5117 108267 5151
rect 108209 5111 108267 5117
rect 89588 5052 89668 5080
rect 94225 5083 94283 5089
rect 89588 5040 89594 5052
rect 94225 5049 94237 5083
rect 94271 5080 94283 5083
rect 94593 5083 94651 5089
rect 94593 5080 94605 5083
rect 94271 5052 94605 5080
rect 94271 5049 94283 5052
rect 94225 5043 94283 5049
rect 94593 5049 94605 5052
rect 94639 5080 94651 5083
rect 94961 5083 95019 5089
rect 94961 5080 94973 5083
rect 94639 5052 94973 5080
rect 94639 5049 94651 5052
rect 94593 5043 94651 5049
rect 94961 5049 94973 5052
rect 95007 5080 95019 5083
rect 102042 5080 102048 5092
rect 95007 5052 102048 5080
rect 95007 5049 95019 5052
rect 94961 5043 95019 5049
rect 102042 5040 102048 5052
rect 102100 5040 102106 5092
rect 106292 5080 106320 5111
rect 108390 5108 108396 5160
rect 108448 5148 108454 5160
rect 110598 5148 110604 5160
rect 108448 5120 110604 5148
rect 108448 5108 108454 5120
rect 110598 5108 110604 5120
rect 110656 5108 110662 5160
rect 111797 5151 111855 5157
rect 111797 5117 111809 5151
rect 111843 5117 111855 5151
rect 111797 5111 111855 5117
rect 105740 5052 106320 5080
rect 17126 4972 17132 5024
rect 17184 5012 17190 5024
rect 33226 5012 33232 5024
rect 17184 4984 33232 5012
rect 17184 4972 17190 4984
rect 33226 4972 33232 4984
rect 33284 4972 33290 5024
rect 40310 4972 40316 5024
rect 40368 5012 40374 5024
rect 42058 5012 42064 5024
rect 40368 4984 42064 5012
rect 40368 4972 40374 4984
rect 42058 4972 42064 4984
rect 42116 4972 42122 5024
rect 47854 4972 47860 5024
rect 47912 5012 47918 5024
rect 48133 5015 48191 5021
rect 48133 5012 48145 5015
rect 47912 4984 48145 5012
rect 47912 4972 47918 4984
rect 48133 4981 48145 4984
rect 48179 4981 48191 5015
rect 48133 4975 48191 4981
rect 51902 4972 51908 5024
rect 51960 4972 51966 5024
rect 51994 4972 52000 5024
rect 52052 5012 52058 5024
rect 78122 5012 78128 5024
rect 52052 4984 78128 5012
rect 52052 4972 52058 4984
rect 78122 4972 78128 4984
rect 78180 4972 78186 5024
rect 84289 5015 84347 5021
rect 84289 4981 84301 5015
rect 84335 5012 84347 5015
rect 84654 5012 84660 5024
rect 84335 4984 84660 5012
rect 84335 4981 84347 4984
rect 84289 4975 84347 4981
rect 84654 4972 84660 4984
rect 84712 4972 84718 5024
rect 84838 4972 84844 5024
rect 84896 5012 84902 5024
rect 89898 5012 89904 5024
rect 84896 4984 89904 5012
rect 84896 4972 84902 4984
rect 89898 4972 89904 4984
rect 89956 4972 89962 5024
rect 94130 4972 94136 5024
rect 94188 5012 94194 5024
rect 99650 5012 99656 5024
rect 94188 4984 99656 5012
rect 94188 4972 94194 4984
rect 99650 4972 99656 4984
rect 99708 4972 99714 5024
rect 103514 4972 103520 5024
rect 103572 5012 103578 5024
rect 105740 5021 105768 5052
rect 106642 5040 106648 5092
rect 106700 5080 106706 5092
rect 106737 5083 106795 5089
rect 106737 5080 106749 5083
rect 106700 5052 106749 5080
rect 106700 5040 106706 5052
rect 106737 5049 106749 5052
rect 106783 5049 106795 5083
rect 111429 5083 111487 5089
rect 111429 5080 111441 5083
rect 106737 5043 106795 5049
rect 107672 5052 111441 5080
rect 105725 5015 105783 5021
rect 105725 5012 105737 5015
rect 103572 4984 105737 5012
rect 103572 4972 103578 4984
rect 105725 4981 105737 4984
rect 105771 4981 105783 5015
rect 105725 4975 105783 4981
rect 105814 4972 105820 5024
rect 105872 5012 105878 5024
rect 107672 5012 107700 5052
rect 111429 5049 111441 5052
rect 111475 5080 111487 5083
rect 111812 5080 111840 5111
rect 111978 5108 111984 5160
rect 112036 5108 112042 5160
rect 112717 5151 112775 5157
rect 112717 5148 112729 5151
rect 112548 5120 112729 5148
rect 112438 5080 112444 5092
rect 111475 5052 111840 5080
rect 112364 5052 112444 5080
rect 111475 5049 111487 5052
rect 111429 5043 111487 5049
rect 105872 4984 107700 5012
rect 105872 4972 105878 4984
rect 107930 4972 107936 5024
rect 107988 4972 107994 5024
rect 110230 4972 110236 5024
rect 110288 5012 110294 5024
rect 112364 5012 112392 5052
rect 112438 5040 112444 5052
rect 112496 5040 112502 5092
rect 110288 4984 112392 5012
rect 112548 5012 112576 5120
rect 112717 5117 112729 5120
rect 112763 5117 112775 5151
rect 112717 5111 112775 5117
rect 112806 5108 112812 5160
rect 112864 5157 112870 5160
rect 112864 5151 112892 5157
rect 112880 5117 112892 5151
rect 112864 5111 112892 5117
rect 112993 5151 113051 5157
rect 112993 5117 113005 5151
rect 113039 5148 113051 5151
rect 113174 5148 113180 5160
rect 113039 5120 113180 5148
rect 113039 5117 113051 5120
rect 112993 5111 113051 5117
rect 112864 5108 112870 5111
rect 113174 5108 113180 5120
rect 113232 5108 113238 5160
rect 114186 5108 114192 5160
rect 114244 5148 114250 5160
rect 115109 5151 115167 5157
rect 115109 5148 115121 5151
rect 114244 5120 115121 5148
rect 114244 5108 114250 5120
rect 115109 5117 115121 5120
rect 115155 5117 115167 5151
rect 115109 5111 115167 5117
rect 115569 5151 115627 5157
rect 115569 5117 115581 5151
rect 115615 5148 115627 5151
rect 116762 5148 116768 5160
rect 115615 5120 116768 5148
rect 115615 5117 115627 5120
rect 115569 5111 115627 5117
rect 114278 5080 114284 5092
rect 113376 5052 114284 5080
rect 113376 5012 113404 5052
rect 114278 5040 114284 5052
rect 114336 5040 114342 5092
rect 115584 5080 115612 5111
rect 116762 5108 116768 5120
rect 116820 5108 116826 5160
rect 117590 5108 117596 5160
rect 117648 5108 117654 5160
rect 118326 5108 118332 5160
rect 118384 5157 118390 5160
rect 118510 5157 118516 5160
rect 118384 5151 118405 5157
rect 118393 5117 118405 5151
rect 118384 5111 118405 5117
rect 118467 5151 118516 5157
rect 118467 5117 118479 5151
rect 118513 5117 118516 5151
rect 118467 5111 118516 5117
rect 118384 5108 118390 5111
rect 118510 5108 118516 5111
rect 118568 5108 118574 5160
rect 118605 5151 118663 5157
rect 118605 5117 118617 5151
rect 118651 5148 118663 5151
rect 119430 5148 119436 5160
rect 118651 5120 119436 5148
rect 118651 5117 118663 5120
rect 118605 5111 118663 5117
rect 119430 5108 119436 5120
rect 119488 5108 119494 5160
rect 120261 5151 120319 5157
rect 120261 5117 120273 5151
rect 120307 5148 120319 5151
rect 120442 5148 120448 5160
rect 120307 5120 120448 5148
rect 120307 5117 120319 5120
rect 120261 5111 120319 5117
rect 120442 5108 120448 5120
rect 120500 5108 120506 5160
rect 120810 5108 120816 5160
rect 120868 5148 120874 5160
rect 121114 5151 121172 5157
rect 121114 5148 121126 5151
rect 120868 5120 121126 5148
rect 120868 5108 120874 5120
rect 121114 5117 121126 5120
rect 121160 5117 121172 5151
rect 121114 5111 121172 5117
rect 121273 5151 121331 5157
rect 121273 5117 121285 5151
rect 121319 5148 121331 5151
rect 121319 5120 122420 5148
rect 121319 5117 121331 5120
rect 121273 5111 121331 5117
rect 118050 5080 118056 5092
rect 114756 5052 115612 5080
rect 117332 5052 118056 5080
rect 112548 4984 113404 5012
rect 110288 4972 110294 4984
rect 113634 4972 113640 5024
rect 113692 4972 113698 5024
rect 113726 4972 113732 5024
rect 113784 5012 113790 5024
rect 114756 5021 114784 5052
rect 114097 5015 114155 5021
rect 114097 5012 114109 5015
rect 113784 4984 114109 5012
rect 113784 4972 113790 4984
rect 114097 4981 114109 4984
rect 114143 5012 114155 5015
rect 114741 5015 114799 5021
rect 114741 5012 114753 5015
rect 114143 4984 114753 5012
rect 114143 4981 114155 4984
rect 114097 4975 114155 4981
rect 114741 4981 114753 4984
rect 114787 4981 114799 5015
rect 114741 4975 114799 4981
rect 115290 4972 115296 5024
rect 115348 5012 115354 5024
rect 117332 5012 117360 5052
rect 118050 5040 118056 5052
rect 118108 5040 118114 5092
rect 119893 5083 119951 5089
rect 119893 5080 119905 5083
rect 119172 5052 119905 5080
rect 115348 4984 117360 5012
rect 115348 4972 115354 4984
rect 117406 4972 117412 5024
rect 117464 5012 117470 5024
rect 119172 5012 119200 5052
rect 119893 5049 119905 5052
rect 119939 5049 119951 5083
rect 119893 5043 119951 5049
rect 120718 5040 120724 5092
rect 120776 5040 120782 5092
rect 117464 4984 119200 5012
rect 117464 4972 117470 4984
rect 119430 4972 119436 5024
rect 119488 5012 119494 5024
rect 120350 5012 120356 5024
rect 119488 4984 120356 5012
rect 119488 4972 119494 4984
rect 120350 4972 120356 4984
rect 120408 5012 120414 5024
rect 121656 5012 121684 5120
rect 122392 5089 122420 5120
rect 122377 5083 122435 5089
rect 122377 5049 122389 5083
rect 122423 5049 122435 5083
rect 122377 5043 122435 5049
rect 120408 4984 121684 5012
rect 120408 4972 120414 4984
rect 121914 4972 121920 5024
rect 121972 4972 121978 5024
rect 137986 5012 138014 5188
rect 149882 5176 149888 5228
rect 149940 5216 149946 5228
rect 150621 5219 150679 5225
rect 150621 5216 150633 5219
rect 149940 5188 150633 5216
rect 149940 5176 149946 5188
rect 150621 5185 150633 5188
rect 150667 5185 150679 5219
rect 157306 5216 157334 5324
rect 157794 5312 157800 5324
rect 157852 5352 157858 5364
rect 158165 5355 158223 5361
rect 158165 5352 158177 5355
rect 157852 5324 158177 5352
rect 157852 5312 157858 5324
rect 158165 5321 158177 5324
rect 158211 5352 158223 5355
rect 158211 5324 162716 5352
rect 158211 5321 158223 5324
rect 158165 5315 158223 5321
rect 159450 5244 159456 5296
rect 159508 5284 159514 5296
rect 162578 5284 162584 5296
rect 159508 5256 162584 5284
rect 159508 5244 159514 5256
rect 162578 5244 162584 5256
rect 162636 5244 162642 5296
rect 162688 5284 162716 5324
rect 163038 5312 163044 5364
rect 163096 5312 163102 5364
rect 163222 5312 163228 5364
rect 163280 5352 163286 5364
rect 175918 5352 175924 5364
rect 163280 5324 175924 5352
rect 163280 5312 163286 5324
rect 175918 5312 175924 5324
rect 175976 5312 175982 5364
rect 176626 5324 190454 5352
rect 176626 5284 176654 5324
rect 162688 5256 176654 5284
rect 188430 5244 188436 5296
rect 188488 5284 188494 5296
rect 188488 5256 188844 5284
rect 188488 5244 188494 5256
rect 150621 5179 150679 5185
rect 154500 5188 157334 5216
rect 150802 5108 150808 5160
rect 150860 5108 150866 5160
rect 150894 5108 150900 5160
rect 150952 5148 150958 5160
rect 150952 5120 151124 5148
rect 150952 5108 150958 5120
rect 151096 5080 151124 5120
rect 151354 5108 151360 5160
rect 151412 5148 151418 5160
rect 151722 5157 151728 5160
rect 151541 5151 151599 5157
rect 151541 5148 151553 5151
rect 151412 5120 151553 5148
rect 151412 5108 151418 5120
rect 151541 5117 151553 5120
rect 151587 5117 151599 5151
rect 151541 5111 151599 5117
rect 151679 5151 151728 5157
rect 151679 5117 151691 5151
rect 151725 5117 151728 5151
rect 151679 5111 151728 5117
rect 151722 5108 151728 5111
rect 151780 5108 151786 5160
rect 151814 5108 151820 5160
rect 151872 5108 151878 5160
rect 152366 5108 152372 5160
rect 152424 5148 152430 5160
rect 153105 5151 153163 5157
rect 153105 5148 153117 5151
rect 152424 5120 153117 5148
rect 152424 5108 152430 5120
rect 153105 5117 153117 5120
rect 153151 5117 153163 5151
rect 153565 5151 153623 5157
rect 153565 5148 153577 5151
rect 153105 5111 153163 5117
rect 153304 5120 153577 5148
rect 151265 5083 151323 5089
rect 151265 5080 151277 5083
rect 151096 5052 151277 5080
rect 151265 5049 151277 5052
rect 151311 5049 151323 5083
rect 151265 5043 151323 5049
rect 152737 5015 152795 5021
rect 152737 5012 152749 5015
rect 137986 4984 152749 5012
rect 152737 4981 152749 4984
rect 152783 5012 152795 5015
rect 153304 5012 153332 5120
rect 153565 5117 153577 5120
rect 153611 5148 153623 5151
rect 154500 5148 154528 5188
rect 161106 5176 161112 5228
rect 161164 5216 161170 5228
rect 161382 5216 161388 5228
rect 161164 5188 161388 5216
rect 161164 5176 161170 5188
rect 161382 5176 161388 5188
rect 161440 5176 161446 5228
rect 161566 5176 161572 5228
rect 161624 5176 161630 5228
rect 163133 5219 163191 5225
rect 163133 5216 163145 5219
rect 162136 5188 163145 5216
rect 153611 5120 154528 5148
rect 153611 5117 153623 5120
rect 153565 5111 153623 5117
rect 155862 5108 155868 5160
rect 155920 5148 155926 5160
rect 155920 5120 158208 5148
rect 155920 5108 155926 5120
rect 155405 5083 155463 5089
rect 155405 5080 155417 5083
rect 154546 5052 155417 5080
rect 152783 4984 153332 5012
rect 152783 4981 152795 4984
rect 152737 4975 152795 4981
rect 153746 4972 153752 5024
rect 153804 5012 153810 5024
rect 154546 5012 154574 5052
rect 155405 5049 155417 5052
rect 155451 5080 155463 5083
rect 158070 5080 158076 5092
rect 155451 5052 158076 5080
rect 155451 5049 155463 5052
rect 155405 5043 155463 5049
rect 158070 5040 158076 5052
rect 158128 5040 158134 5092
rect 158180 5080 158208 5120
rect 158254 5108 158260 5160
rect 158312 5108 158318 5160
rect 158441 5151 158499 5157
rect 158441 5117 158453 5151
rect 158487 5148 158499 5151
rect 158530 5148 158536 5160
rect 158487 5120 158536 5148
rect 158487 5117 158499 5120
rect 158441 5111 158499 5117
rect 158530 5108 158536 5120
rect 158588 5108 158594 5160
rect 160002 5108 160008 5160
rect 160060 5108 160066 5160
rect 162136 5092 162164 5188
rect 163133 5185 163145 5188
rect 163179 5216 163191 5219
rect 163179 5188 163452 5216
rect 163179 5185 163191 5188
rect 163133 5179 163191 5185
rect 162670 5148 162676 5160
rect 162596 5120 162676 5148
rect 161198 5080 161204 5092
rect 158180 5052 161204 5080
rect 161198 5040 161204 5052
rect 161256 5040 161262 5092
rect 162118 5040 162124 5092
rect 162176 5040 162182 5092
rect 162596 5089 162624 5120
rect 162670 5108 162676 5120
rect 162728 5108 162734 5160
rect 162581 5083 162639 5089
rect 162581 5049 162593 5083
rect 162627 5049 162639 5083
rect 162581 5043 162639 5049
rect 153804 4984 154574 5012
rect 153804 4972 153810 4984
rect 156046 4972 156052 5024
rect 156104 5012 156110 5024
rect 156782 5012 156788 5024
rect 156104 4984 156788 5012
rect 156104 4972 156110 4984
rect 156782 4972 156788 4984
rect 156840 5012 156846 5024
rect 158622 5012 158628 5024
rect 156840 4984 158628 5012
rect 156840 4972 156846 4984
rect 158622 4972 158628 4984
rect 158680 4972 158686 5024
rect 160002 4972 160008 5024
rect 160060 5012 160066 5024
rect 160465 5015 160523 5021
rect 160465 5012 160477 5015
rect 160060 4984 160477 5012
rect 160060 4972 160066 4984
rect 160465 4981 160477 4984
rect 160511 5012 160523 5015
rect 161566 5012 161572 5024
rect 160511 4984 161572 5012
rect 160511 4981 160523 4984
rect 160465 4975 160523 4981
rect 161566 4972 161572 4984
rect 161624 4972 161630 5024
rect 162946 4972 162952 5024
rect 163004 5012 163010 5024
rect 163317 5015 163375 5021
rect 163317 5012 163329 5015
rect 163004 4984 163329 5012
rect 163004 4972 163010 4984
rect 163317 4981 163329 4984
rect 163363 4981 163375 5015
rect 163424 5012 163452 5188
rect 163498 5176 163504 5228
rect 163556 5216 163562 5228
rect 180610 5216 180616 5228
rect 163556 5188 180616 5216
rect 163556 5176 163562 5188
rect 180610 5176 180616 5188
rect 180668 5176 180674 5228
rect 181993 5219 182051 5225
rect 181993 5185 182005 5219
rect 182039 5216 182051 5219
rect 182082 5216 182088 5228
rect 182039 5188 182088 5216
rect 182039 5185 182051 5188
rect 181993 5179 182051 5185
rect 182082 5176 182088 5188
rect 182140 5176 182146 5228
rect 182174 5176 182180 5228
rect 182232 5176 182238 5228
rect 182542 5176 182548 5228
rect 182600 5176 182606 5228
rect 188816 5225 188844 5256
rect 189166 5244 189172 5296
rect 189224 5244 189230 5296
rect 190426 5284 190454 5324
rect 212506 5324 215800 5352
rect 212506 5284 212534 5324
rect 190426 5256 212534 5284
rect 215772 5284 215800 5324
rect 215846 5312 215852 5364
rect 215904 5352 215910 5364
rect 218146 5352 218152 5364
rect 215904 5324 218152 5352
rect 215904 5312 215910 5324
rect 218146 5312 218152 5324
rect 218204 5312 218210 5364
rect 218900 5324 221136 5352
rect 218900 5293 218928 5324
rect 218241 5287 218299 5293
rect 218241 5284 218253 5287
rect 215772 5256 218253 5284
rect 218241 5253 218253 5256
rect 218287 5284 218299 5287
rect 218517 5287 218575 5293
rect 218517 5284 218529 5287
rect 218287 5256 218529 5284
rect 218287 5253 218299 5256
rect 218241 5247 218299 5253
rect 218517 5253 218529 5256
rect 218563 5284 218575 5287
rect 218885 5287 218943 5293
rect 218885 5284 218897 5287
rect 218563 5256 218897 5284
rect 218563 5253 218575 5256
rect 218517 5247 218575 5253
rect 218885 5253 218897 5256
rect 218931 5253 218943 5287
rect 218885 5247 218943 5253
rect 219437 5287 219495 5293
rect 219437 5253 219449 5287
rect 219483 5284 219495 5287
rect 220170 5284 220176 5296
rect 219483 5256 220176 5284
rect 219483 5253 219495 5256
rect 219437 5247 219495 5253
rect 220170 5244 220176 5256
rect 220228 5244 220234 5296
rect 221108 5293 221136 5324
rect 221752 5324 234614 5352
rect 221752 5293 221780 5324
rect 221093 5287 221151 5293
rect 221093 5253 221105 5287
rect 221139 5284 221151 5287
rect 221369 5287 221427 5293
rect 221369 5284 221381 5287
rect 221139 5256 221381 5284
rect 221139 5253 221151 5256
rect 221093 5247 221151 5253
rect 221369 5253 221381 5256
rect 221415 5284 221427 5287
rect 221737 5287 221795 5293
rect 221737 5284 221749 5287
rect 221415 5256 221749 5284
rect 221415 5253 221427 5256
rect 221369 5247 221427 5253
rect 221737 5253 221749 5256
rect 221783 5253 221795 5287
rect 224678 5284 224684 5296
rect 221737 5247 221795 5253
rect 222304 5256 224684 5284
rect 222304 5228 222332 5256
rect 224678 5244 224684 5256
rect 224736 5244 224742 5296
rect 227346 5284 227352 5296
rect 225708 5256 227352 5284
rect 188801 5219 188859 5225
rect 188801 5185 188813 5219
rect 188847 5216 188859 5219
rect 188847 5188 190454 5216
rect 188847 5185 188859 5188
rect 188801 5179 188859 5185
rect 177942 5148 177948 5160
rect 163608 5120 177948 5148
rect 163608 5012 163636 5120
rect 177942 5108 177948 5120
rect 178000 5108 178006 5160
rect 164234 5040 164240 5092
rect 164292 5080 164298 5092
rect 175826 5080 175832 5092
rect 164292 5052 175832 5080
rect 164292 5040 164298 5052
rect 175826 5040 175832 5052
rect 175884 5040 175890 5092
rect 182542 5040 182548 5092
rect 182600 5040 182606 5092
rect 190426 5080 190454 5188
rect 215772 5188 219204 5216
rect 214006 5108 214012 5160
rect 214064 5108 214070 5160
rect 214190 5108 214196 5160
rect 214248 5148 214254 5160
rect 215772 5148 215800 5188
rect 214248 5120 215800 5148
rect 215849 5151 215907 5157
rect 214248 5108 214254 5120
rect 215849 5117 215861 5151
rect 215895 5148 215907 5151
rect 216582 5148 216588 5160
rect 215895 5120 216588 5148
rect 215895 5117 215907 5120
rect 215849 5111 215907 5117
rect 216582 5108 216588 5120
rect 216640 5108 216646 5160
rect 219176 5148 219204 5188
rect 219250 5176 219256 5228
rect 219308 5176 219314 5228
rect 222286 5176 222292 5228
rect 222344 5176 222350 5228
rect 222378 5176 222384 5228
rect 222436 5216 222442 5228
rect 225708 5225 225736 5256
rect 227346 5244 227352 5256
rect 227404 5244 227410 5296
rect 227530 5244 227536 5296
rect 227588 5284 227594 5296
rect 228177 5287 228235 5293
rect 228177 5284 228189 5287
rect 227588 5256 228189 5284
rect 227588 5244 227594 5256
rect 228177 5253 228189 5256
rect 228223 5284 228235 5287
rect 228266 5284 228272 5296
rect 228223 5256 228272 5284
rect 228223 5253 228235 5256
rect 228177 5247 228235 5253
rect 228266 5244 228272 5256
rect 228324 5244 228330 5296
rect 228818 5284 228824 5296
rect 228468 5256 228824 5284
rect 228468 5225 228496 5256
rect 228818 5244 228824 5256
rect 228876 5284 228882 5296
rect 229925 5287 229983 5293
rect 229925 5284 229937 5287
rect 228876 5256 229937 5284
rect 228876 5244 228882 5256
rect 229925 5253 229937 5256
rect 229971 5253 229983 5287
rect 229925 5247 229983 5253
rect 230842 5244 230848 5296
rect 230900 5284 230906 5296
rect 231305 5287 231363 5293
rect 231305 5284 231317 5287
rect 230900 5256 231317 5284
rect 230900 5244 230906 5256
rect 231305 5253 231317 5256
rect 231351 5253 231363 5287
rect 234586 5284 234614 5324
rect 238662 5312 238668 5364
rect 238720 5352 238726 5364
rect 238720 5324 260328 5352
rect 238720 5312 238726 5324
rect 239214 5284 239220 5296
rect 234586 5256 239220 5284
rect 231305 5247 231363 5253
rect 239214 5244 239220 5256
rect 239272 5244 239278 5296
rect 239401 5287 239459 5293
rect 239401 5253 239413 5287
rect 239447 5284 239459 5287
rect 239447 5256 239536 5284
rect 239447 5253 239459 5256
rect 239401 5247 239459 5253
rect 222841 5219 222899 5225
rect 222841 5216 222853 5219
rect 222436 5188 222853 5216
rect 222436 5176 222442 5188
rect 222841 5185 222853 5188
rect 222887 5185 222899 5219
rect 222841 5179 222899 5185
rect 225693 5219 225751 5225
rect 225693 5185 225705 5219
rect 225739 5185 225751 5219
rect 225693 5179 225751 5185
rect 228453 5219 228511 5225
rect 228453 5185 228465 5219
rect 228499 5185 228511 5219
rect 228453 5179 228511 5185
rect 230014 5176 230020 5228
rect 230072 5176 230078 5228
rect 230474 5176 230480 5228
rect 230532 5216 230538 5228
rect 231854 5216 231860 5228
rect 230532 5188 231860 5216
rect 230532 5176 230538 5188
rect 231854 5176 231860 5188
rect 231912 5176 231918 5228
rect 238662 5176 238668 5228
rect 238720 5176 238726 5228
rect 238849 5219 238907 5225
rect 238849 5185 238861 5219
rect 238895 5216 238907 5219
rect 239306 5216 239312 5228
rect 238895 5188 239312 5216
rect 238895 5185 238907 5188
rect 238849 5179 238907 5185
rect 239306 5176 239312 5188
rect 239364 5176 239370 5228
rect 223025 5151 223083 5157
rect 223025 5148 223037 5151
rect 219176 5120 223037 5148
rect 223025 5117 223037 5120
rect 223071 5148 223083 5151
rect 223850 5148 223856 5160
rect 223071 5120 223856 5148
rect 223071 5117 223083 5120
rect 223025 5111 223083 5117
rect 223850 5108 223856 5120
rect 223908 5148 223914 5160
rect 225877 5151 225935 5157
rect 225877 5148 225889 5151
rect 223908 5120 225889 5148
rect 223908 5108 223914 5120
rect 225877 5117 225889 5120
rect 225923 5148 225935 5151
rect 225966 5148 225972 5160
rect 225923 5120 225972 5148
rect 225923 5117 225935 5120
rect 225877 5111 225935 5117
rect 225966 5108 225972 5120
rect 226024 5148 226030 5160
rect 226794 5148 226800 5160
rect 226024 5120 226800 5148
rect 226024 5108 226030 5120
rect 226794 5108 226800 5120
rect 226852 5148 226858 5160
rect 228729 5151 228787 5157
rect 228729 5148 228741 5151
rect 226852 5120 228741 5148
rect 226852 5108 226858 5120
rect 228729 5117 228741 5120
rect 228775 5117 228787 5151
rect 239214 5148 239220 5160
rect 228729 5111 228787 5117
rect 229296 5120 239220 5148
rect 215018 5080 215024 5092
rect 190426 5052 215024 5080
rect 215018 5040 215024 5052
rect 215076 5040 215082 5092
rect 215938 5040 215944 5092
rect 215996 5080 216002 5092
rect 215996 5052 218836 5080
rect 215996 5040 216002 5052
rect 163424 4984 163636 5012
rect 189169 5015 189227 5021
rect 163317 4975 163375 4981
rect 189169 4981 189181 5015
rect 189215 5012 189227 5015
rect 189258 5012 189264 5024
rect 189215 4984 189264 5012
rect 189215 4981 189227 4984
rect 189169 4975 189227 4981
rect 189258 4972 189264 4984
rect 189316 4972 189322 5024
rect 189353 5015 189411 5021
rect 189353 4981 189365 5015
rect 189399 5012 189411 5015
rect 189994 5012 190000 5024
rect 189399 4984 190000 5012
rect 189399 4981 189411 4984
rect 189353 4975 189411 4981
rect 189994 4972 190000 4984
rect 190052 4972 190058 5024
rect 210050 4972 210056 5024
rect 210108 5012 210114 5024
rect 218698 5012 218704 5024
rect 210108 4984 218704 5012
rect 210108 4972 210114 4984
rect 218698 4972 218704 4984
rect 218756 4972 218762 5024
rect 218808 5012 218836 5052
rect 226334 5040 226340 5092
rect 226392 5080 226398 5092
rect 229296 5080 229324 5120
rect 239214 5108 239220 5120
rect 239272 5108 239278 5160
rect 226392 5052 229324 5080
rect 226392 5040 226398 5052
rect 230658 5040 230664 5092
rect 230716 5080 230722 5092
rect 230937 5083 230995 5089
rect 230937 5080 230949 5083
rect 230716 5052 230949 5080
rect 230716 5040 230722 5052
rect 230937 5049 230949 5052
rect 230983 5049 230995 5083
rect 230937 5043 230995 5049
rect 231026 5040 231032 5092
rect 231084 5080 231090 5092
rect 239508 5080 239536 5256
rect 239674 5244 239680 5296
rect 239732 5284 239738 5296
rect 255774 5284 255780 5296
rect 239732 5256 255780 5284
rect 239732 5244 239738 5256
rect 255774 5244 255780 5256
rect 255832 5244 255838 5296
rect 239582 5176 239588 5228
rect 239640 5216 239646 5228
rect 240229 5219 240287 5225
rect 240229 5216 240241 5219
rect 239640 5188 240241 5216
rect 239640 5176 239646 5188
rect 240229 5185 240241 5188
rect 240275 5185 240287 5219
rect 251450 5216 251456 5228
rect 240229 5179 240287 5185
rect 240428 5188 251456 5216
rect 240428 5089 240456 5188
rect 251450 5176 251456 5188
rect 251508 5176 251514 5228
rect 253566 5148 253572 5160
rect 244246 5120 253572 5148
rect 240413 5083 240471 5089
rect 240413 5080 240425 5083
rect 231084 5052 240425 5080
rect 231084 5040 231090 5052
rect 240413 5049 240425 5052
rect 240459 5049 240471 5083
rect 244246 5080 244274 5120
rect 253566 5108 253572 5120
rect 253624 5108 253630 5160
rect 260300 5148 260328 5324
rect 262214 5312 262220 5364
rect 262272 5352 262278 5364
rect 264885 5355 264943 5361
rect 264885 5352 264897 5355
rect 262272 5324 264897 5352
rect 262272 5312 262278 5324
rect 264885 5321 264897 5324
rect 264931 5321 264943 5355
rect 264885 5315 264943 5321
rect 266722 5312 266728 5364
rect 266780 5352 266786 5364
rect 267093 5355 267151 5361
rect 267093 5352 267105 5355
rect 266780 5324 267105 5352
rect 266780 5312 266786 5324
rect 267093 5321 267105 5324
rect 267139 5321 267151 5355
rect 267093 5315 267151 5321
rect 267734 5312 267740 5364
rect 267792 5312 267798 5364
rect 267826 5312 267832 5364
rect 267884 5352 267890 5364
rect 268657 5355 268715 5361
rect 268657 5352 268669 5355
rect 267884 5324 268669 5352
rect 267884 5312 267890 5324
rect 268657 5321 268669 5324
rect 268703 5321 268715 5355
rect 268657 5315 268715 5321
rect 269022 5312 269028 5364
rect 269080 5352 269086 5364
rect 269669 5355 269727 5361
rect 269669 5352 269681 5355
rect 269080 5324 269681 5352
rect 269080 5312 269086 5324
rect 269669 5321 269681 5324
rect 269715 5321 269727 5355
rect 269669 5315 269727 5321
rect 271138 5312 271144 5364
rect 271196 5352 271202 5364
rect 271966 5352 271972 5364
rect 271196 5324 271972 5352
rect 271196 5312 271202 5324
rect 271966 5312 271972 5324
rect 272024 5312 272030 5364
rect 261849 5287 261907 5293
rect 261849 5284 261861 5287
rect 260392 5256 261861 5284
rect 260392 5225 260420 5256
rect 261849 5253 261861 5256
rect 261895 5253 261907 5287
rect 261849 5247 261907 5253
rect 261938 5244 261944 5296
rect 261996 5284 262002 5296
rect 266265 5287 266323 5293
rect 266265 5284 266277 5287
rect 261996 5256 266277 5284
rect 261996 5244 262002 5256
rect 266265 5253 266277 5256
rect 266311 5253 266323 5287
rect 266265 5247 266323 5253
rect 267274 5244 267280 5296
rect 267332 5284 267338 5296
rect 270497 5287 270555 5293
rect 270497 5284 270509 5287
rect 267332 5256 270509 5284
rect 267332 5244 267338 5256
rect 270497 5253 270509 5256
rect 270543 5253 270555 5287
rect 270497 5247 270555 5253
rect 260377 5219 260435 5225
rect 260377 5185 260389 5219
rect 260423 5185 260435 5219
rect 261665 5219 261723 5225
rect 261665 5216 261677 5219
rect 260377 5179 260435 5185
rect 260484 5188 261677 5216
rect 260484 5148 260512 5188
rect 261665 5185 261677 5188
rect 261711 5216 261723 5219
rect 262490 5216 262496 5228
rect 261711 5188 262496 5216
rect 261711 5185 261723 5188
rect 261665 5179 261723 5185
rect 262490 5176 262496 5188
rect 262548 5176 262554 5228
rect 262950 5176 262956 5228
rect 263008 5176 263014 5228
rect 264698 5176 264704 5228
rect 264756 5176 264762 5228
rect 265986 5176 265992 5228
rect 266044 5176 266050 5228
rect 266081 5219 266139 5225
rect 266081 5185 266093 5219
rect 266127 5216 266139 5219
rect 266170 5216 266176 5228
rect 266127 5188 266176 5216
rect 266127 5185 266139 5188
rect 266081 5179 266139 5185
rect 266170 5176 266176 5188
rect 266228 5216 266234 5228
rect 266909 5219 266967 5225
rect 266909 5216 266921 5219
rect 266228 5188 266921 5216
rect 266228 5176 266234 5188
rect 266909 5185 266921 5188
rect 266955 5185 266967 5219
rect 266909 5179 266967 5185
rect 267458 5176 267464 5228
rect 267516 5216 267522 5228
rect 267553 5219 267611 5225
rect 267553 5216 267565 5219
rect 267516 5188 267565 5216
rect 267516 5176 267522 5188
rect 267553 5185 267565 5188
rect 267599 5185 267611 5219
rect 267553 5179 267611 5185
rect 268473 5219 268531 5225
rect 268473 5185 268485 5219
rect 268519 5216 268531 5219
rect 268654 5216 268660 5228
rect 268519 5188 268660 5216
rect 268519 5185 268531 5188
rect 268473 5179 268531 5185
rect 268654 5176 268660 5188
rect 268712 5216 268718 5228
rect 269485 5219 269543 5225
rect 269485 5216 269497 5219
rect 268712 5188 269497 5216
rect 268712 5176 268718 5188
rect 269485 5185 269497 5188
rect 269531 5216 269543 5219
rect 269758 5216 269764 5228
rect 269531 5188 269764 5216
rect 269531 5185 269543 5188
rect 269485 5179 269543 5185
rect 269758 5176 269764 5188
rect 269816 5216 269822 5228
rect 270313 5219 270371 5225
rect 270313 5216 270325 5219
rect 269816 5188 270325 5216
rect 269816 5176 269822 5188
rect 270313 5185 270325 5188
rect 270359 5216 270371 5219
rect 270402 5216 270408 5228
rect 270359 5188 270408 5216
rect 270359 5185 270371 5188
rect 270313 5179 270371 5185
rect 270402 5176 270408 5188
rect 270460 5176 270466 5228
rect 260300 5120 260512 5148
rect 260650 5108 260656 5160
rect 260708 5108 260714 5160
rect 261481 5151 261539 5157
rect 261481 5117 261493 5151
rect 261527 5117 261539 5151
rect 261481 5111 261539 5117
rect 240413 5043 240471 5049
rect 241486 5052 244274 5080
rect 261496 5080 261524 5111
rect 263226 5108 263232 5160
rect 263284 5108 263290 5160
rect 264517 5151 264575 5157
rect 264517 5117 264529 5151
rect 264563 5117 264575 5151
rect 264517 5111 264575 5117
rect 264422 5080 264428 5092
rect 261496 5052 264428 5080
rect 224862 5012 224868 5024
rect 218808 4984 224868 5012
rect 224862 4972 224868 4984
rect 224920 4972 224926 5024
rect 225049 5015 225107 5021
rect 225049 4981 225061 5015
rect 225095 5012 225107 5015
rect 225230 5012 225236 5024
rect 225095 4984 225236 5012
rect 225095 4981 225107 4984
rect 225049 4975 225107 4981
rect 225230 4972 225236 4984
rect 225288 5012 225294 5024
rect 225417 5015 225475 5021
rect 225417 5012 225429 5015
rect 225288 4984 225429 5012
rect 225288 4972 225294 4984
rect 225417 4981 225429 4984
rect 225463 5012 225475 5015
rect 227530 5012 227536 5024
rect 225463 4984 227536 5012
rect 225463 4981 225475 4984
rect 225417 4975 225475 4981
rect 227530 4972 227536 4984
rect 227588 4972 227594 5024
rect 227714 4972 227720 5024
rect 227772 5012 227778 5024
rect 229002 5012 229008 5024
rect 227772 4984 229008 5012
rect 227772 4972 227778 4984
rect 229002 4972 229008 4984
rect 229060 4972 229066 5024
rect 231302 4972 231308 5024
rect 231360 4972 231366 5024
rect 231489 5015 231547 5021
rect 231489 4981 231501 5015
rect 231535 5012 231547 5015
rect 235626 5012 235632 5024
rect 231535 4984 235632 5012
rect 231535 4981 231547 4984
rect 231489 4975 231547 4981
rect 235626 4972 235632 4984
rect 235684 4972 235690 5024
rect 239214 4972 239220 5024
rect 239272 5012 239278 5024
rect 239493 5015 239551 5021
rect 239493 5012 239505 5015
rect 239272 4984 239505 5012
rect 239272 4972 239278 4984
rect 239493 4981 239505 4984
rect 239539 4981 239551 5015
rect 239493 4975 239551 4981
rect 239582 4972 239588 5024
rect 239640 5012 239646 5024
rect 241486 5012 241514 5052
rect 264422 5040 264428 5052
rect 264480 5040 264486 5092
rect 264532 5080 264560 5111
rect 265158 5108 265164 5160
rect 265216 5148 265222 5160
rect 266725 5151 266783 5157
rect 266725 5148 266737 5151
rect 265216 5120 266737 5148
rect 265216 5108 265222 5120
rect 266725 5117 266737 5120
rect 266771 5117 266783 5151
rect 266725 5111 266783 5117
rect 268286 5108 268292 5160
rect 268344 5108 268350 5160
rect 269298 5108 269304 5160
rect 269356 5108 269362 5160
rect 270129 5151 270187 5157
rect 270129 5117 270141 5151
rect 270175 5117 270187 5151
rect 270129 5111 270187 5117
rect 266630 5080 266636 5092
rect 264532 5052 266636 5080
rect 266630 5040 266636 5052
rect 266688 5040 266694 5092
rect 267458 5040 267464 5092
rect 267516 5080 267522 5092
rect 268838 5080 268844 5092
rect 267516 5052 268844 5080
rect 267516 5040 267522 5052
rect 268838 5040 268844 5052
rect 268896 5040 268902 5092
rect 269206 5040 269212 5092
rect 269264 5080 269270 5092
rect 270144 5080 270172 5111
rect 269264 5052 270172 5080
rect 269264 5040 269270 5052
rect 239640 4984 241514 5012
rect 241977 5015 242035 5021
rect 239640 4972 239646 4984
rect 241977 4981 241989 5015
rect 242023 5012 242035 5015
rect 242250 5012 242256 5024
rect 242023 4984 242256 5012
rect 242023 4981 242035 4984
rect 241977 4975 242035 4981
rect 242250 4972 242256 4984
rect 242308 4972 242314 5024
rect 242618 4972 242624 5024
rect 242676 4972 242682 5024
rect 242710 4972 242716 5024
rect 242768 5012 242774 5024
rect 245562 5012 245568 5024
rect 242768 4984 245568 5012
rect 242768 4972 242774 4984
rect 245562 4972 245568 4984
rect 245620 4972 245626 5024
rect 252462 4972 252468 5024
rect 252520 5012 252526 5024
rect 256878 5012 256884 5024
rect 252520 4984 256884 5012
rect 252520 4972 252526 4984
rect 256878 4972 256884 4984
rect 256936 4972 256942 5024
rect 258534 4972 258540 5024
rect 258592 5012 258598 5024
rect 259089 5015 259147 5021
rect 259089 5012 259101 5015
rect 258592 4984 259101 5012
rect 258592 4972 258598 4984
rect 259089 4981 259101 4984
rect 259135 4981 259147 5015
rect 259089 4975 259147 4981
rect 259454 4972 259460 5024
rect 259512 5012 259518 5024
rect 259825 5015 259883 5021
rect 259825 5012 259837 5015
rect 259512 4984 259837 5012
rect 259512 4972 259518 4984
rect 259825 4981 259837 4984
rect 259871 4981 259883 5015
rect 259825 4975 259883 4981
rect 266814 4972 266820 5024
rect 266872 5012 266878 5024
rect 271966 5012 271972 5024
rect 266872 4984 271972 5012
rect 266872 4972 266878 4984
rect 271966 4972 271972 4984
rect 272024 4972 272030 5024
rect 1104 4922 271492 4944
rect 1104 4870 34748 4922
rect 34800 4870 34812 4922
rect 34864 4870 34876 4922
rect 34928 4870 34940 4922
rect 34992 4870 35004 4922
rect 35056 4870 102345 4922
rect 102397 4870 102409 4922
rect 102461 4870 102473 4922
rect 102525 4870 102537 4922
rect 102589 4870 102601 4922
rect 102653 4870 169942 4922
rect 169994 4870 170006 4922
rect 170058 4870 170070 4922
rect 170122 4870 170134 4922
rect 170186 4870 170198 4922
rect 170250 4870 237539 4922
rect 237591 4870 237603 4922
rect 237655 4870 237667 4922
rect 237719 4870 237731 4922
rect 237783 4870 237795 4922
rect 237847 4870 271492 4922
rect 1104 4848 271492 4870
rect 12158 4768 12164 4820
rect 12216 4808 12222 4820
rect 35894 4808 35900 4820
rect 12216 4780 35900 4808
rect 12216 4768 12222 4780
rect 35894 4768 35900 4780
rect 35952 4768 35958 4820
rect 40954 4808 40960 4820
rect 39868 4780 40960 4808
rect 34606 4700 34612 4752
rect 34664 4740 34670 4752
rect 39758 4740 39764 4752
rect 34664 4712 39764 4740
rect 34664 4700 34670 4712
rect 39758 4700 39764 4712
rect 39816 4700 39822 4752
rect 33134 4632 33140 4684
rect 33192 4672 33198 4684
rect 39868 4672 39896 4780
rect 40954 4768 40960 4780
rect 41012 4768 41018 4820
rect 42518 4768 42524 4820
rect 42576 4808 42582 4820
rect 42613 4811 42671 4817
rect 42613 4808 42625 4811
rect 42576 4780 42625 4808
rect 42576 4768 42582 4780
rect 42613 4777 42625 4780
rect 42659 4777 42671 4811
rect 42613 4771 42671 4777
rect 48777 4811 48835 4817
rect 48777 4777 48789 4811
rect 48823 4808 48835 4811
rect 52086 4808 52092 4820
rect 48823 4780 52092 4808
rect 48823 4777 48835 4780
rect 48777 4771 48835 4777
rect 52086 4768 52092 4780
rect 52144 4768 52150 4820
rect 74534 4768 74540 4820
rect 74592 4808 74598 4820
rect 82906 4808 82912 4820
rect 74592 4780 82912 4808
rect 74592 4768 74598 4780
rect 82906 4768 82912 4780
rect 82964 4768 82970 4820
rect 84654 4768 84660 4820
rect 84712 4808 84718 4820
rect 84712 4780 89714 4808
rect 84712 4768 84718 4780
rect 51166 4700 51172 4752
rect 51224 4740 51230 4752
rect 51994 4740 52000 4752
rect 51224 4712 52000 4740
rect 51224 4700 51230 4712
rect 51994 4700 52000 4712
rect 52052 4700 52058 4752
rect 84746 4740 84752 4752
rect 64846 4712 84752 4740
rect 53104 4684 53156 4690
rect 33192 4644 39896 4672
rect 33192 4632 33198 4644
rect 41138 4632 41144 4684
rect 41196 4632 41202 4684
rect 44726 4672 44732 4684
rect 44022 4644 44732 4672
rect 44726 4632 44732 4644
rect 44784 4632 44790 4684
rect 48038 4632 48044 4684
rect 48096 4632 48102 4684
rect 53104 4626 53156 4632
rect 36538 4564 36544 4616
rect 36596 4604 36602 4616
rect 36596 4576 42748 4604
rect 36596 4564 36602 4576
rect 40052 4508 41184 4536
rect 8478 4428 8484 4480
rect 8536 4468 8542 4480
rect 40052 4477 40080 4508
rect 40037 4471 40095 4477
rect 40037 4468 40049 4471
rect 8536 4440 40049 4468
rect 8536 4428 8542 4440
rect 40037 4437 40049 4440
rect 40083 4437 40095 4471
rect 40037 4431 40095 4437
rect 40310 4428 40316 4480
rect 40368 4468 40374 4480
rect 40405 4471 40463 4477
rect 40405 4468 40417 4471
rect 40368 4440 40417 4468
rect 40368 4428 40374 4440
rect 40405 4437 40417 4440
rect 40451 4437 40463 4471
rect 40405 4431 40463 4437
rect 40954 4428 40960 4480
rect 41012 4428 41018 4480
rect 41156 4468 41184 4508
rect 41230 4496 41236 4548
rect 41288 4496 41294 4548
rect 41325 4539 41383 4545
rect 41325 4505 41337 4539
rect 41371 4536 41383 4539
rect 41598 4536 41604 4548
rect 41371 4508 41604 4536
rect 41371 4505 41383 4508
rect 41325 4499 41383 4505
rect 41598 4496 41604 4508
rect 41656 4496 41662 4548
rect 41693 4539 41751 4545
rect 41693 4505 41705 4539
rect 41739 4505 41751 4539
rect 41693 4499 41751 4505
rect 41708 4468 41736 4499
rect 42058 4496 42064 4548
rect 42116 4496 42122 4548
rect 42720 4536 42748 4576
rect 43254 4564 43260 4616
rect 43312 4564 43318 4616
rect 43349 4607 43407 4613
rect 43349 4573 43361 4607
rect 43395 4604 43407 4607
rect 43622 4604 43628 4616
rect 43395 4576 43628 4604
rect 43395 4573 43407 4576
rect 43349 4567 43407 4573
rect 43622 4564 43628 4576
rect 43680 4564 43686 4616
rect 47762 4564 47768 4616
rect 47820 4564 47826 4616
rect 48130 4564 48136 4616
rect 48188 4604 48194 4616
rect 48607 4607 48665 4613
rect 48607 4604 48619 4607
rect 48188 4576 48619 4604
rect 48188 4564 48194 4576
rect 48607 4573 48619 4576
rect 48653 4573 48665 4607
rect 48607 4567 48665 4573
rect 52365 4607 52423 4613
rect 52365 4573 52377 4607
rect 52411 4573 52423 4607
rect 52365 4567 52423 4573
rect 43717 4539 43775 4545
rect 42720 4508 43300 4536
rect 41156 4440 41736 4468
rect 42242 4428 42248 4480
rect 42300 4428 42306 4480
rect 42981 4471 43039 4477
rect 42981 4437 42993 4471
rect 43027 4468 43039 4471
rect 43070 4468 43076 4480
rect 43027 4440 43076 4468
rect 43027 4437 43039 4440
rect 42981 4431 43039 4437
rect 43070 4428 43076 4440
rect 43128 4428 43134 4480
rect 43272 4468 43300 4508
rect 43717 4505 43729 4539
rect 43763 4536 43775 4539
rect 43990 4536 43996 4548
rect 43763 4508 43996 4536
rect 43763 4505 43775 4508
rect 43717 4499 43775 4505
rect 43990 4496 43996 4508
rect 44048 4496 44054 4548
rect 45189 4539 45247 4545
rect 45189 4536 45201 4539
rect 44100 4508 45201 4536
rect 44100 4477 44128 4508
rect 45189 4505 45201 4508
rect 45235 4505 45247 4539
rect 45189 4499 45247 4505
rect 46842 4496 46848 4548
rect 46900 4536 46906 4548
rect 47210 4536 47216 4548
rect 46900 4508 47216 4536
rect 46900 4496 46906 4508
rect 47210 4496 47216 4508
rect 47268 4536 47274 4548
rect 47854 4536 47860 4548
rect 47268 4508 47860 4536
rect 47268 4496 47274 4508
rect 47854 4496 47860 4508
rect 47912 4496 47918 4548
rect 48222 4496 48228 4548
rect 48280 4496 48286 4548
rect 48866 4536 48872 4548
rect 48516 4508 48872 4536
rect 44085 4471 44143 4477
rect 44085 4468 44097 4471
rect 43272 4440 44097 4468
rect 44085 4437 44097 4440
rect 44131 4437 44143 4471
rect 44085 4431 44143 4437
rect 44266 4428 44272 4480
rect 44324 4428 44330 4480
rect 46934 4428 46940 4480
rect 46992 4428 46998 4480
rect 47489 4471 47547 4477
rect 47489 4437 47501 4471
rect 47535 4468 47547 4471
rect 48516 4468 48544 4508
rect 48866 4496 48872 4508
rect 48924 4496 48930 4548
rect 48976 4508 52224 4536
rect 47535 4440 48544 4468
rect 47535 4437 47547 4440
rect 47489 4431 47547 4437
rect 48590 4428 48596 4480
rect 48648 4468 48654 4480
rect 48976 4468 49004 4508
rect 48648 4440 49004 4468
rect 48648 4428 48654 4440
rect 50982 4428 50988 4480
rect 51040 4468 51046 4480
rect 51350 4468 51356 4480
rect 51040 4440 51356 4468
rect 51040 4428 51046 4440
rect 51350 4428 51356 4440
rect 51408 4428 51414 4480
rect 51994 4428 52000 4480
rect 52052 4468 52058 4480
rect 52089 4471 52147 4477
rect 52089 4468 52101 4471
rect 52052 4440 52101 4468
rect 52052 4428 52058 4440
rect 52089 4437 52101 4440
rect 52135 4437 52147 4471
rect 52196 4468 52224 4508
rect 52270 4496 52276 4548
rect 52328 4536 52334 4548
rect 52376 4536 52404 4567
rect 52328 4508 52404 4536
rect 52328 4496 52334 4508
rect 52454 4496 52460 4548
rect 52512 4496 52518 4548
rect 52822 4496 52828 4548
rect 52880 4496 52886 4548
rect 64846 4536 64874 4712
rect 84746 4700 84752 4712
rect 84804 4700 84810 4752
rect 85574 4700 85580 4752
rect 85632 4740 85638 4752
rect 86770 4740 86776 4752
rect 85632 4712 86776 4740
rect 85632 4700 85638 4712
rect 86770 4700 86776 4712
rect 86828 4700 86834 4752
rect 89686 4740 89714 4780
rect 91002 4768 91008 4820
rect 91060 4808 91066 4820
rect 91060 4780 113864 4808
rect 91060 4768 91066 4780
rect 99374 4740 99380 4752
rect 89686 4712 99380 4740
rect 99374 4700 99380 4712
rect 99432 4700 99438 4752
rect 99469 4743 99527 4749
rect 99469 4709 99481 4743
rect 99515 4740 99527 4743
rect 99834 4740 99840 4752
rect 99515 4712 99840 4740
rect 99515 4709 99527 4712
rect 99469 4703 99527 4709
rect 99834 4700 99840 4712
rect 99892 4700 99898 4752
rect 100938 4740 100944 4752
rect 99944 4712 100944 4740
rect 78122 4632 78128 4684
rect 78180 4672 78186 4684
rect 81713 4675 81771 4681
rect 81713 4672 81725 4675
rect 78180 4644 81725 4672
rect 78180 4632 78186 4644
rect 81713 4641 81725 4644
rect 81759 4641 81771 4675
rect 81713 4635 81771 4641
rect 81894 4632 81900 4684
rect 81952 4672 81958 4684
rect 92477 4675 92535 4681
rect 92477 4672 92489 4675
rect 81952 4644 92489 4672
rect 81952 4632 81958 4644
rect 92477 4641 92489 4644
rect 92523 4641 92535 4675
rect 92477 4635 92535 4641
rect 92658 4632 92664 4684
rect 92716 4632 92722 4684
rect 94317 4675 94375 4681
rect 94317 4641 94329 4675
rect 94363 4672 94375 4675
rect 95234 4672 95240 4684
rect 94363 4644 95240 4672
rect 94363 4641 94375 4644
rect 94317 4635 94375 4641
rect 95234 4632 95240 4644
rect 95292 4632 95298 4684
rect 99944 4681 99972 4712
rect 100938 4700 100944 4712
rect 100996 4700 101002 4752
rect 105538 4700 105544 4752
rect 105596 4740 105602 4752
rect 106642 4740 106648 4752
rect 105596 4712 106648 4740
rect 105596 4700 105602 4712
rect 106642 4700 106648 4712
rect 106700 4740 106706 4752
rect 107654 4740 107660 4752
rect 106700 4712 107660 4740
rect 106700 4700 106706 4712
rect 107654 4700 107660 4712
rect 107712 4700 107718 4752
rect 109402 4700 109408 4752
rect 109460 4740 109466 4752
rect 109460 4712 109816 4740
rect 109460 4700 109466 4712
rect 99929 4675 99987 4681
rect 99929 4641 99941 4675
rect 99975 4641 99987 4675
rect 99929 4635 99987 4641
rect 100021 4675 100079 4681
rect 100021 4641 100033 4675
rect 100067 4672 100079 4675
rect 100570 4672 100576 4684
rect 100067 4644 100576 4672
rect 100067 4641 100079 4644
rect 100021 4635 100079 4641
rect 100570 4632 100576 4644
rect 100628 4632 100634 4684
rect 106366 4632 106372 4684
rect 106424 4672 106430 4684
rect 107197 4675 107255 4681
rect 107197 4672 107209 4675
rect 106424 4644 107209 4672
rect 106424 4632 106430 4644
rect 107197 4641 107209 4644
rect 107243 4641 107255 4675
rect 107197 4635 107255 4641
rect 107933 4675 107991 4681
rect 107933 4641 107945 4675
rect 107979 4672 107991 4675
rect 108390 4672 108396 4684
rect 107979 4644 108396 4672
rect 107979 4641 107991 4644
rect 107933 4635 107991 4641
rect 108390 4632 108396 4644
rect 108448 4632 108454 4684
rect 109788 4681 109816 4712
rect 110230 4700 110236 4752
rect 110288 4740 110294 4752
rect 110417 4743 110475 4749
rect 110417 4740 110429 4743
rect 110288 4712 110429 4740
rect 110288 4700 110294 4712
rect 110417 4709 110429 4712
rect 110463 4709 110475 4743
rect 110417 4703 110475 4709
rect 111613 4743 111671 4749
rect 111613 4709 111625 4743
rect 111659 4740 111671 4743
rect 111794 4740 111800 4752
rect 111659 4712 111800 4740
rect 111659 4709 111671 4712
rect 111613 4703 111671 4709
rect 111794 4700 111800 4712
rect 111852 4700 111858 4752
rect 112990 4700 112996 4752
rect 113048 4740 113054 4752
rect 113726 4740 113732 4752
rect 113048 4712 113732 4740
rect 113048 4700 113054 4712
rect 113726 4700 113732 4712
rect 113784 4700 113790 4752
rect 113836 4740 113864 4780
rect 113910 4768 113916 4820
rect 113968 4808 113974 4820
rect 118878 4808 118884 4820
rect 113968 4780 118884 4808
rect 113968 4768 113974 4780
rect 118878 4768 118884 4780
rect 118936 4768 118942 4820
rect 121825 4811 121883 4817
rect 121825 4808 121837 4811
rect 118988 4780 121837 4808
rect 118988 4740 119016 4780
rect 121825 4777 121837 4780
rect 121871 4777 121883 4811
rect 121825 4771 121883 4777
rect 113836 4712 119016 4740
rect 120718 4700 120724 4752
rect 120776 4740 120782 4752
rect 121840 4740 121868 4771
rect 139302 4768 139308 4820
rect 139360 4808 139366 4820
rect 153746 4808 153752 4820
rect 139360 4780 153752 4808
rect 139360 4768 139366 4780
rect 153746 4768 153752 4780
rect 153804 4768 153810 4820
rect 155405 4811 155463 4817
rect 153856 4780 155356 4808
rect 142798 4740 142804 4752
rect 120776 4712 120948 4740
rect 121840 4712 122972 4740
rect 120776 4700 120782 4712
rect 109773 4675 109831 4681
rect 109773 4641 109785 4675
rect 109819 4641 109831 4675
rect 109773 4635 109831 4641
rect 110690 4632 110696 4684
rect 110748 4632 110754 4684
rect 110831 4675 110889 4681
rect 110831 4641 110843 4675
rect 110877 4672 110889 4675
rect 110877 4644 112484 4672
rect 110877 4641 110889 4644
rect 110831 4635 110889 4641
rect 84010 4564 84016 4616
rect 84068 4564 84074 4616
rect 85853 4607 85911 4613
rect 85853 4573 85865 4607
rect 85899 4604 85911 4607
rect 85899 4576 86540 4604
rect 85899 4573 85911 4576
rect 85853 4567 85911 4573
rect 53116 4508 64874 4536
rect 53116 4468 53144 4508
rect 81618 4496 81624 4548
rect 81676 4536 81682 4548
rect 81897 4539 81955 4545
rect 81897 4536 81909 4539
rect 81676 4508 81909 4536
rect 81676 4496 81682 4508
rect 81897 4505 81909 4508
rect 81943 4505 81955 4539
rect 81897 4499 81955 4505
rect 83553 4539 83611 4545
rect 83553 4505 83565 4539
rect 83599 4505 83611 4539
rect 83553 4499 83611 4505
rect 84197 4539 84255 4545
rect 84197 4505 84209 4539
rect 84243 4536 84255 4539
rect 85574 4536 85580 4548
rect 84243 4508 85580 4536
rect 84243 4505 84255 4508
rect 84197 4499 84255 4505
rect 52196 4440 53144 4468
rect 52089 4431 52147 4437
rect 53190 4428 53196 4480
rect 53248 4428 53254 4480
rect 53374 4428 53380 4480
rect 53432 4428 53438 4480
rect 80333 4471 80391 4477
rect 80333 4437 80345 4471
rect 80379 4468 80391 4471
rect 80701 4471 80759 4477
rect 80701 4468 80713 4471
rect 80379 4440 80713 4468
rect 80379 4437 80391 4440
rect 80333 4431 80391 4437
rect 80701 4437 80713 4440
rect 80747 4468 80759 4471
rect 81437 4471 81495 4477
rect 81437 4468 81449 4471
rect 80747 4440 81449 4468
rect 80747 4437 80759 4440
rect 80701 4431 80759 4437
rect 81437 4437 81449 4440
rect 81483 4468 81495 4471
rect 83568 4468 83596 4499
rect 85574 4496 85580 4508
rect 85632 4496 85638 4548
rect 86402 4496 86408 4548
rect 86460 4496 86466 4548
rect 86420 4468 86448 4496
rect 86512 4477 86540 4576
rect 87874 4564 87880 4616
rect 87932 4564 87938 4616
rect 89272 4576 92520 4604
rect 86678 4496 86684 4548
rect 86736 4536 86742 4548
rect 86736 4508 87644 4536
rect 86736 4496 86742 4508
rect 81483 4440 86448 4468
rect 86497 4471 86555 4477
rect 81483 4437 81495 4440
rect 81437 4431 81495 4437
rect 86497 4437 86509 4471
rect 86543 4468 86555 4471
rect 86865 4471 86923 4477
rect 86865 4468 86877 4471
rect 86543 4440 86877 4468
rect 86543 4437 86555 4440
rect 86497 4431 86555 4437
rect 86865 4437 86877 4440
rect 86911 4468 86923 4471
rect 87233 4471 87291 4477
rect 87233 4468 87245 4471
rect 86911 4440 87245 4468
rect 86911 4437 86923 4440
rect 86865 4431 86923 4437
rect 87233 4437 87245 4440
rect 87279 4468 87291 4471
rect 87506 4468 87512 4480
rect 87279 4440 87512 4468
rect 87279 4437 87291 4440
rect 87233 4431 87291 4437
rect 87506 4428 87512 4440
rect 87564 4428 87570 4480
rect 87616 4468 87644 4508
rect 88058 4496 88064 4548
rect 88116 4496 88122 4548
rect 89272 4468 89300 4576
rect 89717 4539 89775 4545
rect 89717 4505 89729 4539
rect 89763 4536 89775 4539
rect 92492 4536 92520 4576
rect 94406 4564 94412 4616
rect 94464 4564 94470 4616
rect 94501 4607 94559 4613
rect 94501 4573 94513 4607
rect 94547 4604 94559 4607
rect 94869 4607 94927 4613
rect 94869 4604 94881 4607
rect 94547 4576 94881 4604
rect 94547 4573 94559 4576
rect 94501 4567 94559 4573
rect 94869 4573 94881 4576
rect 94915 4573 94927 4607
rect 94869 4567 94927 4573
rect 94958 4564 94964 4616
rect 95016 4604 95022 4616
rect 105814 4604 105820 4616
rect 95016 4576 105820 4604
rect 95016 4564 95022 4576
rect 105814 4564 105820 4576
rect 105872 4564 105878 4616
rect 106274 4564 106280 4616
rect 106332 4604 106338 4616
rect 108114 4613 108120 4616
rect 107013 4607 107071 4613
rect 107013 4604 107025 4607
rect 106332 4576 107025 4604
rect 106332 4564 106338 4576
rect 107013 4573 107025 4576
rect 107059 4573 107071 4607
rect 107013 4567 107071 4573
rect 108071 4607 108120 4613
rect 108071 4573 108083 4607
rect 108117 4573 108120 4607
rect 108071 4567 108120 4573
rect 108114 4564 108120 4567
rect 108172 4564 108178 4616
rect 108206 4564 108212 4616
rect 108264 4564 108270 4616
rect 109954 4564 109960 4616
rect 110012 4564 110018 4616
rect 110966 4564 110972 4616
rect 111024 4564 111030 4616
rect 89763 4508 90128 4536
rect 92492 4508 92612 4536
rect 89763 4505 89775 4508
rect 89717 4499 89775 4505
rect 90100 4477 90128 4508
rect 87616 4440 89300 4468
rect 90085 4471 90143 4477
rect 90085 4437 90097 4471
rect 90131 4468 90143 4471
rect 90453 4471 90511 4477
rect 90453 4468 90465 4471
rect 90131 4440 90465 4468
rect 90131 4437 90143 4440
rect 90085 4431 90143 4437
rect 90453 4437 90465 4440
rect 90499 4468 90511 4471
rect 90821 4471 90879 4477
rect 90821 4468 90833 4471
rect 90499 4440 90833 4468
rect 90499 4437 90511 4440
rect 90453 4431 90511 4437
rect 90821 4437 90833 4440
rect 90867 4468 90879 4471
rect 92474 4468 92480 4480
rect 90867 4440 92480 4468
rect 90867 4437 90879 4440
rect 90821 4431 90879 4437
rect 92474 4428 92480 4440
rect 92532 4428 92538 4480
rect 92584 4468 92612 4508
rect 95050 4496 95056 4548
rect 95108 4536 95114 4548
rect 95237 4539 95295 4545
rect 95237 4536 95249 4539
rect 95108 4508 95249 4536
rect 95108 4496 95114 4508
rect 95237 4505 95249 4508
rect 95283 4505 95295 4539
rect 95237 4499 95295 4505
rect 99466 4496 99472 4548
rect 99524 4496 99530 4548
rect 105446 4536 105452 4548
rect 99852 4508 105452 4536
rect 99852 4468 99880 4508
rect 105446 4496 105452 4508
rect 105504 4496 105510 4548
rect 108758 4496 108764 4548
rect 108816 4536 108822 4548
rect 109862 4536 109868 4548
rect 108816 4508 109868 4536
rect 108816 4496 108822 4508
rect 109862 4496 109868 4508
rect 109920 4496 109926 4548
rect 112456 4536 112484 4644
rect 113634 4632 113640 4684
rect 113692 4672 113698 4684
rect 114097 4675 114155 4681
rect 114097 4672 114109 4675
rect 113692 4644 114109 4672
rect 113692 4632 113698 4644
rect 114097 4641 114109 4644
rect 114143 4641 114155 4675
rect 114097 4635 114155 4641
rect 114281 4675 114339 4681
rect 114281 4641 114293 4675
rect 114327 4672 114339 4675
rect 114370 4672 114376 4684
rect 114327 4644 114376 4672
rect 114327 4641 114339 4644
rect 114281 4635 114339 4641
rect 114370 4632 114376 4644
rect 114428 4632 114434 4684
rect 114462 4632 114468 4684
rect 114520 4672 114526 4684
rect 114557 4675 114615 4681
rect 114557 4672 114569 4675
rect 114520 4644 114569 4672
rect 114520 4632 114526 4644
rect 114557 4641 114569 4644
rect 114603 4672 114615 4675
rect 116210 4672 116216 4684
rect 114603 4644 116216 4672
rect 114603 4641 114615 4644
rect 114557 4635 114615 4641
rect 116210 4632 116216 4644
rect 116268 4632 116274 4684
rect 118234 4632 118240 4684
rect 118292 4632 118298 4684
rect 118881 4675 118939 4681
rect 118881 4672 118893 4675
rect 118344 4644 118893 4672
rect 112530 4564 112536 4616
rect 112588 4604 112594 4616
rect 113910 4604 113916 4616
rect 112588 4576 113916 4604
rect 112588 4564 112594 4576
rect 113910 4564 113916 4576
rect 113968 4564 113974 4616
rect 118050 4564 118056 4616
rect 118108 4604 118114 4616
rect 118344 4604 118372 4644
rect 118881 4641 118893 4644
rect 118927 4672 118939 4675
rect 119798 4672 119804 4684
rect 118927 4644 119804 4672
rect 118927 4641 118939 4644
rect 118881 4635 118939 4641
rect 119798 4632 119804 4644
rect 119856 4672 119862 4684
rect 120920 4681 120948 4712
rect 120905 4675 120963 4681
rect 120905 4672 120917 4675
rect 119856 4644 120917 4672
rect 119856 4632 119862 4644
rect 120905 4641 120917 4644
rect 120951 4641 120963 4675
rect 120905 4635 120963 4641
rect 121914 4632 121920 4684
rect 121972 4672 121978 4684
rect 122944 4681 122972 4712
rect 128326 4712 142804 4740
rect 122469 4675 122527 4681
rect 122469 4672 122481 4675
rect 121972 4644 122481 4672
rect 121972 4632 121978 4644
rect 122469 4641 122481 4644
rect 122515 4641 122527 4675
rect 122469 4635 122527 4641
rect 122929 4675 122987 4681
rect 122929 4641 122941 4675
rect 122975 4672 122987 4675
rect 124585 4675 124643 4681
rect 124585 4672 124597 4675
rect 122975 4644 124597 4672
rect 122975 4641 122987 4644
rect 122929 4635 122987 4641
rect 124585 4641 124597 4644
rect 124631 4672 124643 4675
rect 128326 4672 128354 4712
rect 142798 4700 142804 4712
rect 142856 4700 142862 4752
rect 151078 4700 151084 4752
rect 151136 4740 151142 4752
rect 151136 4712 151308 4740
rect 151136 4700 151142 4712
rect 124631 4644 128354 4672
rect 143077 4675 143135 4681
rect 124631 4641 124643 4644
rect 124585 4635 124643 4641
rect 143077 4641 143089 4675
rect 143123 4672 143135 4675
rect 144822 4672 144828 4684
rect 143123 4644 144828 4672
rect 143123 4641 143135 4644
rect 143077 4635 143135 4641
rect 144822 4632 144828 4644
rect 144880 4632 144886 4684
rect 150434 4632 150440 4684
rect 150492 4672 150498 4684
rect 150529 4675 150587 4681
rect 150529 4672 150541 4675
rect 150492 4644 150541 4672
rect 150492 4632 150498 4644
rect 150529 4641 150541 4644
rect 150575 4641 150587 4675
rect 150529 4635 150587 4641
rect 150894 4632 150900 4684
rect 150952 4672 150958 4684
rect 151170 4672 151176 4684
rect 150952 4644 151176 4672
rect 150952 4632 150958 4644
rect 151170 4632 151176 4644
rect 151228 4632 151234 4684
rect 151280 4672 151308 4712
rect 152458 4700 152464 4752
rect 152516 4740 152522 4752
rect 153856 4749 153884 4780
rect 153841 4743 153899 4749
rect 153841 4740 153853 4743
rect 152516 4712 153853 4740
rect 152516 4700 152522 4712
rect 153841 4709 153853 4712
rect 153887 4709 153899 4743
rect 155328 4740 155356 4780
rect 155405 4777 155417 4811
rect 155451 4808 155463 4811
rect 156598 4808 156604 4820
rect 155451 4780 156604 4808
rect 155451 4777 155463 4780
rect 155405 4771 155463 4777
rect 156598 4768 156604 4780
rect 156656 4808 156662 4820
rect 157242 4808 157248 4820
rect 156656 4780 157248 4808
rect 156656 4768 156662 4780
rect 157242 4768 157248 4780
rect 157300 4768 157306 4820
rect 158530 4808 158536 4820
rect 157536 4780 158536 4808
rect 156046 4740 156052 4752
rect 155328 4712 156052 4740
rect 153841 4703 153899 4709
rect 156046 4700 156052 4712
rect 156104 4700 156110 4752
rect 151725 4675 151783 4681
rect 151725 4672 151737 4675
rect 151280 4644 151737 4672
rect 151725 4641 151737 4644
rect 151771 4641 151783 4675
rect 151725 4635 151783 4641
rect 151906 4632 151912 4684
rect 151964 4672 151970 4684
rect 153197 4675 153255 4681
rect 153197 4672 153209 4675
rect 151964 4644 153209 4672
rect 151964 4632 151970 4644
rect 153197 4641 153209 4644
rect 153243 4641 153255 4675
rect 157536 4672 157564 4780
rect 158530 4768 158536 4780
rect 158588 4768 158594 4820
rect 160002 4768 160008 4820
rect 160060 4808 160066 4820
rect 163222 4808 163228 4820
rect 160060 4780 163228 4808
rect 160060 4768 160066 4780
rect 163222 4768 163228 4780
rect 163280 4768 163286 4820
rect 179874 4808 179880 4820
rect 166966 4780 179880 4808
rect 166966 4672 166994 4780
rect 179874 4768 179880 4780
rect 179932 4768 179938 4820
rect 213914 4808 213920 4820
rect 212552 4780 213920 4808
rect 153197 4635 153255 4641
rect 153304 4644 157564 4672
rect 157720 4644 166994 4672
rect 118108 4576 118372 4604
rect 118108 4564 118114 4576
rect 118418 4564 118424 4616
rect 118476 4564 118482 4616
rect 119154 4564 119160 4616
rect 119212 4564 119218 4616
rect 119246 4564 119252 4616
rect 119304 4613 119310 4616
rect 119304 4607 119332 4613
rect 119320 4573 119332 4607
rect 119304 4567 119332 4573
rect 119304 4564 119310 4567
rect 119430 4564 119436 4616
rect 119488 4564 119494 4616
rect 120445 4607 120503 4613
rect 120445 4573 120457 4607
rect 120491 4604 120503 4607
rect 120721 4607 120779 4613
rect 120721 4604 120733 4607
rect 120491 4576 120733 4604
rect 120491 4573 120503 4576
rect 120445 4567 120503 4573
rect 120721 4573 120733 4576
rect 120767 4604 120779 4607
rect 120767 4576 122052 4604
rect 120767 4573 120779 4576
rect 120721 4567 120779 4573
rect 115014 4536 115020 4548
rect 112456 4508 115020 4536
rect 115014 4496 115020 4508
rect 115072 4496 115078 4548
rect 120460 4536 120488 4567
rect 119908 4508 120488 4536
rect 92584 4440 99880 4468
rect 100202 4428 100208 4480
rect 100260 4428 100266 4480
rect 101306 4428 101312 4480
rect 101364 4468 101370 4480
rect 106274 4468 106280 4480
rect 101364 4440 106280 4468
rect 101364 4428 101370 4440
rect 106274 4428 106280 4440
rect 106332 4428 106338 4480
rect 108850 4428 108856 4480
rect 108908 4428 108914 4480
rect 110966 4428 110972 4480
rect 111024 4468 111030 4480
rect 113174 4468 113180 4480
rect 111024 4440 113180 4468
rect 111024 4428 111030 4440
rect 113174 4428 113180 4440
rect 113232 4428 113238 4480
rect 113358 4428 113364 4480
rect 113416 4468 113422 4480
rect 113729 4471 113787 4477
rect 113729 4468 113741 4471
rect 113416 4440 113741 4468
rect 113416 4428 113422 4440
rect 113729 4437 113741 4440
rect 113775 4468 113787 4471
rect 114462 4468 114468 4480
rect 113775 4440 114468 4468
rect 113775 4437 113787 4440
rect 113729 4431 113787 4437
rect 114462 4428 114468 4440
rect 114520 4428 114526 4480
rect 114646 4428 114652 4480
rect 114704 4468 114710 4480
rect 116394 4468 116400 4480
rect 114704 4440 116400 4468
rect 114704 4428 114710 4440
rect 116394 4428 116400 4440
rect 116452 4428 116458 4480
rect 118878 4428 118884 4480
rect 118936 4468 118942 4480
rect 119908 4468 119936 4508
rect 118936 4440 119936 4468
rect 120077 4471 120135 4477
rect 118936 4428 118942 4440
rect 120077 4437 120089 4471
rect 120123 4468 120135 4471
rect 120258 4468 120264 4480
rect 120123 4440 120264 4468
rect 120123 4437 120135 4440
rect 120077 4431 120135 4437
rect 120258 4428 120264 4440
rect 120316 4428 120322 4480
rect 122024 4468 122052 4576
rect 150710 4564 150716 4616
rect 150768 4564 150774 4616
rect 151446 4564 151452 4616
rect 151504 4564 151510 4616
rect 151630 4613 151636 4616
rect 151587 4607 151636 4613
rect 151587 4573 151599 4607
rect 151633 4573 151636 4607
rect 151587 4567 151636 4573
rect 151630 4564 151636 4567
rect 151688 4564 151694 4616
rect 152366 4564 152372 4616
rect 152424 4564 152430 4616
rect 122650 4496 122656 4548
rect 122708 4496 122714 4548
rect 142154 4496 142160 4548
rect 142212 4536 142218 4548
rect 143261 4539 143319 4545
rect 143261 4536 143273 4539
rect 142212 4508 143273 4536
rect 142212 4496 142218 4508
rect 143261 4505 143273 4508
rect 143307 4536 143319 4539
rect 143350 4536 143356 4548
rect 143307 4508 143356 4536
rect 143307 4505 143319 4508
rect 143261 4499 143319 4505
rect 143350 4496 143356 4508
rect 143408 4496 143414 4548
rect 144917 4539 144975 4545
rect 144917 4505 144929 4539
rect 144963 4536 144975 4539
rect 145190 4536 145196 4548
rect 144963 4508 145196 4536
rect 144963 4505 144975 4508
rect 144917 4499 144975 4505
rect 129918 4468 129924 4480
rect 122024 4440 129924 4468
rect 129918 4428 129924 4440
rect 129976 4428 129982 4480
rect 142430 4428 142436 4480
rect 142488 4468 142494 4480
rect 144932 4468 144960 4499
rect 145190 4496 145196 4508
rect 145248 4496 145254 4548
rect 152274 4496 152280 4548
rect 152332 4536 152338 4548
rect 153304 4536 153332 4644
rect 153378 4564 153384 4616
rect 153436 4564 153442 4616
rect 154114 4564 154120 4616
rect 154172 4564 154178 4616
rect 154298 4613 154304 4616
rect 154255 4607 154304 4613
rect 154255 4573 154267 4607
rect 154301 4573 154304 4607
rect 154255 4567 154304 4573
rect 154298 4564 154304 4567
rect 154356 4564 154362 4616
rect 154390 4564 154396 4616
rect 154448 4564 154454 4616
rect 155037 4607 155095 4613
rect 155037 4573 155049 4607
rect 155083 4604 155095 4607
rect 155957 4607 156015 4613
rect 155957 4604 155969 4607
rect 155083 4576 155969 4604
rect 155083 4573 155095 4576
rect 155037 4567 155095 4573
rect 155957 4573 155969 4576
rect 156003 4573 156015 4607
rect 155957 4567 156015 4573
rect 152332 4508 153332 4536
rect 152332 4496 152338 4508
rect 155862 4496 155868 4548
rect 155920 4536 155926 4548
rect 156141 4539 156199 4545
rect 156141 4536 156153 4539
rect 155920 4508 156153 4536
rect 155920 4496 155926 4508
rect 156141 4505 156153 4508
rect 156187 4505 156199 4539
rect 156141 4499 156199 4505
rect 156414 4496 156420 4548
rect 156472 4536 156478 4548
rect 157720 4536 157748 4644
rect 210694 4632 210700 4684
rect 210752 4672 210758 4684
rect 212552 4681 212580 4780
rect 213914 4768 213920 4780
rect 213972 4768 213978 4820
rect 214006 4768 214012 4820
rect 214064 4808 214070 4820
rect 217045 4811 217103 4817
rect 217045 4808 217057 4811
rect 214064 4780 217057 4808
rect 214064 4768 214070 4780
rect 217045 4777 217057 4780
rect 217091 4777 217103 4811
rect 217045 4771 217103 4777
rect 219710 4768 219716 4820
rect 219768 4808 219774 4820
rect 222470 4808 222476 4820
rect 219768 4780 222476 4808
rect 219768 4768 219774 4780
rect 222470 4768 222476 4780
rect 222528 4808 222534 4820
rect 222749 4811 222807 4817
rect 222749 4808 222761 4811
rect 222528 4780 222761 4808
rect 222528 4768 222534 4780
rect 222749 4777 222761 4780
rect 222795 4808 222807 4811
rect 223117 4811 223175 4817
rect 223117 4808 223129 4811
rect 222795 4780 223129 4808
rect 222795 4777 222807 4780
rect 222749 4771 222807 4777
rect 223117 4777 223129 4780
rect 223163 4808 223175 4811
rect 223206 4808 223212 4820
rect 223163 4780 223212 4808
rect 223163 4777 223175 4780
rect 223117 4771 223175 4777
rect 223206 4768 223212 4780
rect 223264 4768 223270 4820
rect 224678 4768 224684 4820
rect 224736 4808 224742 4820
rect 225049 4811 225107 4817
rect 225049 4808 225061 4811
rect 224736 4780 225061 4808
rect 224736 4768 224742 4780
rect 225049 4777 225061 4780
rect 225095 4777 225107 4811
rect 225049 4771 225107 4777
rect 226334 4768 226340 4820
rect 226392 4808 226398 4820
rect 226392 4780 228404 4808
rect 226392 4768 226398 4780
rect 213454 4700 213460 4752
rect 213512 4740 213518 4752
rect 215478 4740 215484 4752
rect 213512 4712 215484 4740
rect 213512 4700 213518 4712
rect 215478 4700 215484 4712
rect 215536 4740 215542 4752
rect 215846 4740 215852 4752
rect 215536 4712 215852 4740
rect 215536 4700 215542 4712
rect 215846 4700 215852 4712
rect 215904 4700 215910 4752
rect 217410 4700 217416 4752
rect 217468 4740 217474 4752
rect 217468 4712 220768 4740
rect 217468 4700 217474 4712
rect 212537 4675 212595 4681
rect 212537 4672 212549 4675
rect 210752 4644 212549 4672
rect 210752 4632 210758 4644
rect 212537 4641 212549 4644
rect 212583 4641 212595 4675
rect 212537 4635 212595 4641
rect 213270 4632 213276 4684
rect 213328 4672 213334 4684
rect 215205 4675 215263 4681
rect 215205 4672 215217 4675
rect 213328 4644 215217 4672
rect 213328 4632 213334 4644
rect 215205 4641 215217 4644
rect 215251 4641 215263 4675
rect 215205 4635 215263 4641
rect 216398 4632 216404 4684
rect 216456 4632 216462 4684
rect 220630 4632 220636 4684
rect 220688 4632 220694 4684
rect 220740 4672 220768 4712
rect 222010 4700 222016 4752
rect 222068 4740 222074 4752
rect 228266 4740 228272 4752
rect 222068 4712 228272 4740
rect 222068 4700 222074 4712
rect 228266 4700 228272 4712
rect 228324 4700 228330 4752
rect 228376 4740 228404 4780
rect 229738 4768 229744 4820
rect 229796 4808 229802 4820
rect 237190 4808 237196 4820
rect 229796 4780 237196 4808
rect 229796 4768 229802 4780
rect 237190 4768 237196 4780
rect 237248 4768 237254 4820
rect 237282 4768 237288 4820
rect 237340 4808 237346 4820
rect 238297 4811 238355 4817
rect 238297 4808 238309 4811
rect 237340 4780 238309 4808
rect 237340 4768 237346 4780
rect 238297 4777 238309 4780
rect 238343 4808 238355 4811
rect 238665 4811 238723 4817
rect 238665 4808 238677 4811
rect 238343 4780 238677 4808
rect 238343 4777 238355 4780
rect 238297 4771 238355 4777
rect 238665 4777 238677 4780
rect 238711 4808 238723 4811
rect 239953 4811 240011 4817
rect 239953 4808 239965 4811
rect 238711 4780 239965 4808
rect 238711 4777 238723 4780
rect 238665 4771 238723 4777
rect 230750 4740 230756 4752
rect 228376 4712 230756 4740
rect 230750 4700 230756 4712
rect 230808 4700 230814 4752
rect 238772 4672 238800 4780
rect 239953 4777 239965 4780
rect 239999 4777 240011 4811
rect 239953 4771 240011 4777
rect 240318 4768 240324 4820
rect 240376 4808 240382 4820
rect 240962 4808 240968 4820
rect 240376 4780 240968 4808
rect 240376 4768 240382 4780
rect 240962 4768 240968 4780
rect 241020 4808 241026 4820
rect 241885 4811 241943 4817
rect 241885 4808 241897 4811
rect 241020 4780 241897 4808
rect 241020 4768 241026 4780
rect 241885 4777 241897 4780
rect 241931 4808 241943 4811
rect 242618 4808 242624 4820
rect 241931 4780 242624 4808
rect 241931 4777 241943 4780
rect 241885 4771 241943 4777
rect 242618 4768 242624 4780
rect 242676 4768 242682 4820
rect 244274 4768 244280 4820
rect 244332 4808 244338 4820
rect 252462 4808 252468 4820
rect 244332 4780 252468 4808
rect 244332 4768 244338 4780
rect 252462 4768 252468 4780
rect 252520 4768 252526 4820
rect 253566 4768 253572 4820
rect 253624 4808 253630 4820
rect 253624 4780 253934 4808
rect 253624 4768 253630 4780
rect 246482 4740 246488 4752
rect 239140 4712 246488 4740
rect 239033 4675 239091 4681
rect 239033 4672 239045 4675
rect 220740 4644 234614 4672
rect 238772 4644 239045 4672
rect 157886 4564 157892 4616
rect 157944 4604 157950 4616
rect 158349 4607 158407 4613
rect 158349 4604 158361 4607
rect 157944 4576 158361 4604
rect 157944 4564 157950 4576
rect 158349 4573 158361 4576
rect 158395 4573 158407 4607
rect 158349 4567 158407 4573
rect 159744 4576 160968 4604
rect 156472 4508 157748 4536
rect 157797 4539 157855 4545
rect 156472 4496 156478 4508
rect 157797 4505 157809 4539
rect 157843 4536 157855 4539
rect 158070 4536 158076 4548
rect 157843 4508 158076 4536
rect 157843 4505 157855 4508
rect 157797 4499 157855 4505
rect 158070 4496 158076 4508
rect 158128 4496 158134 4548
rect 158530 4496 158536 4548
rect 158588 4536 158594 4548
rect 159744 4536 159772 4576
rect 158588 4508 159772 4536
rect 160189 4539 160247 4545
rect 158588 4496 158594 4508
rect 160189 4505 160201 4539
rect 160235 4536 160247 4539
rect 160557 4539 160615 4545
rect 160557 4536 160569 4539
rect 160235 4508 160569 4536
rect 160235 4505 160247 4508
rect 160189 4499 160247 4505
rect 160557 4505 160569 4508
rect 160603 4536 160615 4539
rect 160830 4536 160836 4548
rect 160603 4508 160836 4536
rect 160603 4505 160615 4508
rect 160557 4499 160615 4505
rect 142488 4440 144960 4468
rect 142488 4428 142494 4440
rect 148962 4428 148968 4480
rect 149020 4468 149026 4480
rect 151814 4468 151820 4480
rect 149020 4440 151820 4468
rect 149020 4428 149026 4440
rect 151814 4428 151820 4440
rect 151872 4468 151878 4480
rect 155218 4468 155224 4480
rect 151872 4440 155224 4468
rect 151872 4428 151878 4440
rect 155218 4428 155224 4440
rect 155276 4468 155282 4480
rect 156322 4468 156328 4480
rect 155276 4440 156328 4468
rect 155276 4428 155282 4440
rect 156322 4428 156328 4440
rect 156380 4428 156386 4480
rect 158162 4428 158168 4480
rect 158220 4468 158226 4480
rect 160204 4468 160232 4499
rect 160830 4496 160836 4508
rect 160888 4496 160894 4548
rect 158220 4440 160232 4468
rect 160940 4468 160968 4576
rect 161014 4564 161020 4616
rect 161072 4564 161078 4616
rect 212353 4607 212411 4613
rect 212353 4573 212365 4607
rect 212399 4573 212411 4607
rect 212353 4567 212411 4573
rect 161198 4496 161204 4548
rect 161256 4496 161262 4548
rect 161382 4496 161388 4548
rect 161440 4536 161446 4548
rect 162857 4539 162915 4545
rect 162857 4536 162869 4539
rect 161440 4508 162869 4536
rect 161440 4496 161446 4508
rect 162857 4505 162869 4508
rect 162903 4536 162915 4539
rect 163130 4536 163136 4548
rect 162903 4508 163136 4536
rect 162903 4505 162915 4508
rect 162857 4499 162915 4505
rect 163130 4496 163136 4508
rect 163188 4496 163194 4548
rect 162026 4468 162032 4480
rect 160940 4440 162032 4468
rect 158220 4428 158226 4440
rect 162026 4428 162032 4440
rect 162084 4428 162090 4480
rect 212368 4468 212396 4567
rect 213914 4564 213920 4616
rect 213972 4604 213978 4616
rect 213972 4576 214328 4604
rect 213972 4564 213978 4576
rect 214098 4496 214104 4548
rect 214156 4536 214162 4548
rect 214193 4539 214251 4545
rect 214193 4536 214205 4539
rect 214156 4508 214205 4536
rect 214156 4496 214162 4508
rect 214193 4505 214205 4508
rect 214239 4505 214251 4539
rect 214300 4536 214328 4576
rect 214558 4564 214564 4616
rect 214616 4604 214622 4616
rect 215389 4607 215447 4613
rect 215389 4604 215401 4607
rect 214616 4576 215401 4604
rect 214616 4564 214622 4576
rect 215389 4573 215401 4576
rect 215435 4573 215447 4607
rect 215389 4567 215447 4573
rect 216122 4564 216128 4616
rect 216180 4564 216186 4616
rect 216306 4613 216312 4616
rect 216263 4607 216312 4613
rect 216263 4573 216275 4607
rect 216309 4573 216312 4607
rect 216263 4567 216312 4573
rect 216306 4564 216312 4567
rect 216364 4564 216370 4616
rect 222470 4564 222476 4616
rect 222528 4564 222534 4616
rect 226150 4564 226156 4616
rect 226208 4604 226214 4616
rect 226521 4607 226579 4613
rect 226521 4604 226533 4607
rect 226208 4576 226533 4604
rect 226208 4564 226214 4576
rect 226521 4573 226533 4576
rect 226567 4573 226579 4607
rect 226521 4567 226579 4573
rect 228818 4564 228824 4616
rect 228876 4564 228882 4616
rect 231210 4564 231216 4616
rect 231268 4564 231274 4616
rect 231305 4607 231363 4613
rect 231305 4573 231317 4607
rect 231351 4604 231363 4607
rect 231486 4604 231492 4616
rect 231351 4576 231492 4604
rect 231351 4573 231363 4576
rect 231305 4567 231363 4573
rect 231486 4564 231492 4576
rect 231544 4564 231550 4616
rect 234586 4604 234614 4644
rect 239033 4641 239045 4644
rect 239079 4641 239091 4675
rect 239033 4635 239091 4641
rect 239140 4604 239168 4712
rect 246482 4700 246488 4712
rect 246540 4700 246546 4752
rect 241149 4675 241207 4681
rect 241149 4672 241161 4675
rect 240888 4644 241161 4672
rect 234586 4576 239168 4604
rect 239214 4564 239220 4616
rect 239272 4604 239278 4616
rect 240888 4604 240916 4644
rect 241149 4641 241161 4644
rect 241195 4672 241207 4675
rect 242805 4675 242863 4681
rect 242805 4672 242817 4675
rect 241195 4644 242817 4672
rect 241195 4641 241207 4644
rect 241149 4635 241207 4641
rect 242805 4641 242817 4644
rect 242851 4672 242863 4675
rect 244093 4675 244151 4681
rect 244093 4672 244105 4675
rect 242851 4644 244105 4672
rect 242851 4641 242863 4644
rect 242805 4635 242863 4641
rect 244093 4641 244105 4644
rect 244139 4672 244151 4675
rect 244139 4644 244274 4672
rect 244139 4641 244151 4644
rect 244093 4635 244151 4641
rect 239272 4576 240916 4604
rect 239272 4564 239278 4576
rect 240962 4564 240968 4616
rect 241020 4564 241026 4616
rect 242250 4564 242256 4616
rect 242308 4604 242314 4616
rect 242621 4607 242679 4613
rect 242621 4604 242633 4607
rect 242308 4576 242633 4604
rect 242308 4564 242314 4576
rect 242621 4573 242633 4576
rect 242667 4573 242679 4607
rect 242621 4567 242679 4573
rect 243909 4607 243967 4613
rect 243909 4573 243921 4607
rect 243955 4573 243967 4607
rect 244246 4604 244274 4644
rect 250622 4632 250628 4684
rect 250680 4672 250686 4684
rect 251269 4675 251327 4681
rect 251269 4672 251281 4675
rect 250680 4644 251281 4672
rect 250680 4632 250686 4644
rect 251269 4641 251281 4644
rect 251315 4672 251327 4675
rect 252189 4675 252247 4681
rect 252189 4672 252201 4675
rect 251315 4644 252201 4672
rect 251315 4641 251327 4644
rect 251269 4635 251327 4641
rect 252189 4641 252201 4644
rect 252235 4641 252247 4675
rect 253906 4672 253934 4780
rect 255774 4768 255780 4820
rect 255832 4808 255838 4820
rect 256694 4808 256700 4820
rect 255832 4780 256700 4808
rect 255832 4768 255838 4780
rect 256694 4768 256700 4780
rect 256752 4808 256758 4820
rect 257985 4811 258043 4817
rect 257985 4808 257997 4811
rect 256752 4780 257997 4808
rect 256752 4768 256758 4780
rect 257985 4777 257997 4780
rect 258031 4808 258043 4811
rect 259454 4808 259460 4820
rect 258031 4780 259460 4808
rect 258031 4777 258043 4780
rect 257985 4771 258043 4777
rect 259454 4768 259460 4780
rect 259512 4768 259518 4820
rect 263042 4768 263048 4820
rect 263100 4768 263106 4820
rect 265158 4768 265164 4820
rect 265216 4768 265222 4820
rect 266906 4768 266912 4820
rect 266964 4768 266970 4820
rect 268562 4768 268568 4820
rect 268620 4808 268626 4820
rect 270313 4811 270371 4817
rect 270313 4808 270325 4811
rect 268620 4780 270325 4808
rect 268620 4768 268626 4780
rect 270313 4777 270325 4780
rect 270359 4777 270371 4811
rect 270313 4771 270371 4777
rect 270497 4811 270555 4817
rect 270497 4777 270509 4811
rect 270543 4808 270555 4811
rect 270954 4808 270960 4820
rect 270543 4780 270960 4808
rect 270543 4777 270555 4780
rect 270497 4771 270555 4777
rect 270954 4768 270960 4780
rect 271012 4768 271018 4820
rect 255314 4740 255320 4752
rect 254412 4712 255320 4740
rect 254412 4681 254440 4712
rect 255314 4700 255320 4712
rect 255372 4700 255378 4752
rect 259270 4700 259276 4752
rect 259328 4740 259334 4752
rect 260745 4743 260803 4749
rect 259328 4712 259684 4740
rect 259328 4700 259334 4712
rect 259656 4681 259684 4712
rect 260745 4709 260757 4743
rect 260791 4740 260803 4743
rect 264054 4740 264060 4752
rect 260791 4712 264060 4740
rect 260791 4709 260803 4712
rect 260745 4703 260803 4709
rect 264054 4700 264060 4712
rect 264112 4700 264118 4752
rect 264238 4700 264244 4752
rect 264296 4740 264302 4752
rect 269669 4743 269727 4749
rect 269669 4740 269681 4743
rect 264296 4712 269681 4740
rect 264296 4700 264302 4712
rect 269669 4709 269681 4712
rect 269715 4709 269727 4743
rect 269669 4703 269727 4709
rect 254029 4675 254087 4681
rect 254029 4672 254041 4675
rect 253906 4644 254041 4672
rect 252189 4635 252247 4641
rect 254029 4641 254041 4644
rect 254075 4672 254087 4675
rect 254397 4675 254455 4681
rect 254397 4672 254409 4675
rect 254075 4644 254409 4672
rect 254075 4641 254087 4644
rect 254029 4635 254087 4641
rect 254397 4641 254409 4644
rect 254443 4641 254455 4675
rect 259641 4675 259699 4681
rect 254397 4635 254455 4641
rect 255516 4644 257844 4672
rect 251358 4604 251364 4616
rect 244246 4576 251364 4604
rect 243909 4567 243967 4573
rect 214300 4508 215294 4536
rect 214193 4499 214251 4505
rect 215110 4468 215116 4480
rect 212368 4440 215116 4468
rect 215110 4428 215116 4440
rect 215168 4428 215174 4480
rect 215266 4468 215294 4508
rect 220170 4496 220176 4548
rect 220228 4536 220234 4548
rect 220817 4539 220875 4545
rect 220817 4536 220829 4539
rect 220228 4508 220829 4536
rect 220228 4496 220234 4508
rect 220817 4505 220829 4508
rect 220863 4536 220875 4539
rect 222010 4536 222016 4548
rect 220863 4508 222016 4536
rect 220863 4505 220875 4508
rect 220817 4499 220875 4505
rect 222010 4496 222016 4508
rect 222068 4496 222074 4548
rect 223666 4496 223672 4548
rect 223724 4536 223730 4548
rect 225877 4539 225935 4545
rect 223724 4508 224954 4536
rect 223724 4496 223730 4508
rect 218882 4468 218888 4480
rect 215266 4440 218888 4468
rect 218882 4428 218888 4440
rect 218940 4428 218946 4480
rect 224926 4468 224954 4508
rect 225877 4505 225889 4539
rect 225923 4536 225935 4539
rect 226242 4536 226248 4548
rect 225923 4508 226248 4536
rect 225923 4505 225935 4508
rect 225877 4499 225935 4505
rect 226242 4496 226248 4508
rect 226300 4496 226306 4548
rect 226705 4539 226763 4545
rect 226705 4505 226717 4539
rect 226751 4536 226763 4539
rect 226794 4536 226800 4548
rect 226751 4508 226800 4536
rect 226751 4505 226763 4508
rect 226705 4499 226763 4505
rect 226794 4496 226800 4508
rect 226852 4496 226858 4548
rect 228361 4539 228419 4545
rect 228361 4505 228373 4539
rect 228407 4536 228419 4539
rect 228726 4536 228732 4548
rect 228407 4508 228732 4536
rect 228407 4505 228419 4508
rect 228361 4499 228419 4505
rect 228726 4496 228732 4508
rect 228784 4496 228790 4548
rect 229557 4539 229615 4545
rect 229557 4505 229569 4539
rect 229603 4505 229615 4539
rect 229557 4499 229615 4505
rect 226610 4468 226616 4480
rect 224926 4440 226616 4468
rect 226610 4428 226616 4440
rect 226668 4428 226674 4480
rect 228266 4428 228272 4480
rect 228324 4468 228330 4480
rect 229572 4468 229600 4499
rect 230750 4496 230756 4548
rect 230808 4496 230814 4548
rect 243541 4539 243599 4545
rect 243541 4536 243553 4539
rect 230860 4508 243553 4536
rect 228324 4440 229600 4468
rect 228324 4428 228330 4440
rect 230290 4428 230296 4480
rect 230348 4468 230354 4480
rect 230860 4468 230888 4508
rect 243541 4505 243553 4508
rect 243587 4536 243599 4539
rect 243924 4536 243952 4567
rect 251358 4564 251364 4576
rect 251416 4564 251422 4616
rect 251450 4564 251456 4616
rect 251508 4564 251514 4616
rect 255038 4564 255044 4616
rect 255096 4564 255102 4616
rect 255516 4604 255544 4644
rect 255240 4576 255544 4604
rect 244553 4539 244611 4545
rect 243587 4508 244274 4536
rect 243587 4505 243599 4508
rect 243541 4499 243599 4505
rect 230348 4440 230888 4468
rect 230348 4428 230354 4440
rect 231486 4428 231492 4480
rect 231544 4428 231550 4480
rect 239674 4428 239680 4480
rect 239732 4428 239738 4480
rect 241606 4428 241612 4480
rect 241664 4428 241670 4480
rect 243262 4428 243268 4480
rect 243320 4428 243326 4480
rect 244246 4468 244274 4508
rect 244553 4505 244565 4539
rect 244599 4536 244611 4539
rect 245105 4539 245163 4545
rect 245105 4536 245117 4539
rect 244599 4508 245117 4536
rect 244599 4505 244611 4508
rect 244553 4499 244611 4505
rect 245105 4505 245117 4508
rect 245151 4505 245163 4539
rect 251468 4536 251496 4564
rect 251468 4508 253934 4536
rect 245105 4499 245163 4505
rect 244829 4471 244887 4477
rect 244829 4468 244841 4471
rect 244246 4440 244841 4468
rect 244829 4437 244841 4440
rect 244875 4437 244887 4471
rect 244829 4431 244887 4437
rect 245378 4428 245384 4480
rect 245436 4428 245442 4480
rect 251910 4428 251916 4480
rect 251968 4428 251974 4480
rect 253906 4468 253934 4508
rect 254026 4496 254032 4548
rect 254084 4536 254090 4548
rect 254489 4539 254547 4545
rect 254489 4536 254501 4539
rect 254084 4508 254501 4536
rect 254084 4496 254090 4508
rect 254489 4505 254501 4508
rect 254535 4536 254547 4539
rect 255240 4536 255268 4576
rect 256694 4564 256700 4616
rect 256752 4604 256758 4616
rect 257065 4607 257123 4613
rect 257065 4604 257077 4607
rect 256752 4576 257077 4604
rect 256752 4564 256758 4576
rect 257065 4573 257077 4576
rect 257111 4573 257123 4607
rect 257065 4567 257123 4573
rect 257249 4607 257307 4613
rect 257249 4573 257261 4607
rect 257295 4573 257307 4607
rect 257249 4567 257307 4573
rect 254535 4508 255268 4536
rect 254535 4505 254547 4508
rect 254489 4499 254547 4505
rect 255314 4496 255320 4548
rect 255372 4496 255378 4548
rect 257264 4536 257292 4567
rect 257816 4548 257844 4644
rect 259641 4641 259653 4675
rect 259687 4641 259699 4675
rect 266173 4675 266231 4681
rect 266173 4672 266185 4675
rect 259641 4635 259699 4641
rect 263796 4644 266185 4672
rect 258166 4564 258172 4616
rect 258224 4564 258230 4616
rect 258353 4607 258411 4613
rect 258353 4573 258365 4607
rect 258399 4604 258411 4607
rect 259825 4607 259883 4613
rect 259825 4604 259837 4607
rect 258399 4576 259837 4604
rect 258399 4573 258411 4576
rect 258353 4567 258411 4573
rect 259825 4573 259837 4576
rect 259871 4573 259883 4607
rect 259825 4567 259883 4573
rect 263229 4607 263287 4613
rect 263229 4573 263241 4607
rect 263275 4604 263287 4607
rect 263318 4604 263324 4616
rect 263275 4576 263324 4604
rect 263275 4573 263287 4576
rect 263229 4567 263287 4573
rect 256712 4508 257292 4536
rect 256712 4480 256740 4508
rect 257798 4496 257804 4548
rect 257856 4536 257862 4548
rect 258368 4536 258396 4567
rect 263318 4564 263324 4576
rect 263376 4564 263382 4616
rect 263796 4613 263824 4644
rect 266173 4641 266185 4644
rect 266219 4641 266231 4675
rect 266173 4635 266231 4641
rect 266262 4632 266268 4684
rect 266320 4672 266326 4684
rect 267734 4672 267740 4684
rect 266320 4644 267740 4672
rect 266320 4632 266326 4644
rect 267734 4632 267740 4644
rect 267792 4632 267798 4684
rect 263781 4607 263839 4613
rect 263781 4573 263793 4607
rect 263827 4573 263839 4607
rect 263781 4567 263839 4573
rect 265345 4607 265403 4613
rect 265345 4573 265357 4607
rect 265391 4573 265403 4607
rect 265345 4567 265403 4573
rect 257856 4508 258396 4536
rect 258813 4539 258871 4545
rect 257856 4496 257862 4508
rect 258813 4505 258825 4539
rect 258859 4536 258871 4539
rect 259730 4536 259736 4548
rect 258859 4508 259736 4536
rect 258859 4505 258871 4508
rect 258813 4499 258871 4505
rect 259730 4496 259736 4508
rect 259788 4496 259794 4548
rect 260098 4496 260104 4548
rect 260156 4536 260162 4548
rect 260469 4539 260527 4545
rect 260469 4536 260481 4539
rect 260156 4508 260481 4536
rect 260156 4496 260162 4508
rect 260469 4505 260481 4508
rect 260515 4505 260527 4539
rect 260469 4499 260527 4505
rect 264146 4496 264152 4548
rect 264204 4496 264210 4548
rect 265360 4536 265388 4567
rect 265802 4564 265808 4616
rect 265860 4564 265866 4616
rect 265894 4564 265900 4616
rect 265952 4604 265958 4616
rect 265989 4607 266047 4613
rect 265989 4604 266001 4607
rect 265952 4576 266001 4604
rect 265952 4564 265958 4576
rect 265989 4573 266001 4576
rect 266035 4573 266047 4607
rect 265989 4567 266047 4573
rect 266078 4564 266084 4616
rect 266136 4604 266142 4616
rect 266725 4607 266783 4613
rect 266725 4604 266737 4607
rect 266136 4576 266737 4604
rect 266136 4564 266142 4576
rect 266725 4573 266737 4576
rect 266771 4573 266783 4607
rect 266725 4567 266783 4573
rect 267366 4564 267372 4616
rect 267424 4604 267430 4616
rect 267461 4607 267519 4613
rect 267461 4604 267473 4607
rect 267424 4576 267473 4604
rect 267424 4564 267430 4576
rect 267461 4573 267473 4576
rect 267507 4573 267519 4607
rect 267461 4567 267519 4573
rect 267550 4564 267556 4616
rect 267608 4604 267614 4616
rect 267645 4607 267703 4613
rect 267645 4604 267657 4607
rect 267608 4576 267657 4604
rect 267608 4564 267614 4576
rect 267645 4573 267657 4576
rect 267691 4573 267703 4607
rect 267645 4567 267703 4573
rect 268194 4564 268200 4616
rect 268252 4564 268258 4616
rect 269114 4564 269120 4616
rect 269172 4604 269178 4616
rect 269301 4607 269359 4613
rect 269301 4604 269313 4607
rect 269172 4576 269313 4604
rect 269172 4564 269178 4576
rect 269301 4573 269313 4576
rect 269347 4573 269359 4607
rect 269301 4567 269359 4573
rect 269485 4607 269543 4613
rect 269485 4573 269497 4607
rect 269531 4604 269543 4607
rect 269758 4604 269764 4616
rect 269531 4576 269764 4604
rect 269531 4573 269543 4576
rect 269485 4567 269543 4573
rect 269758 4564 269764 4576
rect 269816 4564 269822 4616
rect 271138 4564 271144 4616
rect 271196 4604 271202 4616
rect 272150 4604 272156 4616
rect 271196 4576 272156 4604
rect 271196 4564 271202 4576
rect 272150 4564 272156 4576
rect 272208 4564 272214 4616
rect 268470 4536 268476 4548
rect 265360 4508 268476 4536
rect 268470 4496 268476 4508
rect 268528 4496 268534 4548
rect 268562 4496 268568 4548
rect 268620 4496 268626 4548
rect 270129 4539 270187 4545
rect 270129 4536 270141 4539
rect 268856 4508 270141 4536
rect 256694 4468 256700 4480
rect 253906 4440 256700 4468
rect 256694 4428 256700 4440
rect 256752 4428 256758 4480
rect 257706 4428 257712 4480
rect 257764 4428 257770 4480
rect 260282 4428 260288 4480
rect 260340 4428 260346 4480
rect 267553 4471 267611 4477
rect 267553 4437 267565 4471
rect 267599 4468 267611 4471
rect 268856 4468 268884 4508
rect 270129 4505 270141 4508
rect 270175 4505 270187 4539
rect 270129 4499 270187 4505
rect 270218 4496 270224 4548
rect 270276 4536 270282 4548
rect 270329 4539 270387 4545
rect 270329 4536 270341 4539
rect 270276 4508 270341 4536
rect 270276 4496 270282 4508
rect 270329 4505 270341 4508
rect 270375 4505 270387 4539
rect 270329 4499 270387 4505
rect 267599 4440 268884 4468
rect 267599 4437 267611 4440
rect 267553 4431 267611 4437
rect 1104 4378 271651 4400
rect 1104 4326 68546 4378
rect 68598 4326 68610 4378
rect 68662 4326 68674 4378
rect 68726 4326 68738 4378
rect 68790 4326 68802 4378
rect 68854 4326 136143 4378
rect 136195 4326 136207 4378
rect 136259 4326 136271 4378
rect 136323 4326 136335 4378
rect 136387 4326 136399 4378
rect 136451 4326 203740 4378
rect 203792 4326 203804 4378
rect 203856 4326 203868 4378
rect 203920 4326 203932 4378
rect 203984 4326 203996 4378
rect 204048 4326 271337 4378
rect 271389 4326 271401 4378
rect 271453 4326 271465 4378
rect 271517 4326 271529 4378
rect 271581 4326 271593 4378
rect 271645 4326 271651 4378
rect 1104 4304 271651 4326
rect 23290 4224 23296 4276
rect 23348 4264 23354 4276
rect 23348 4236 31754 4264
rect 23348 4224 23354 4236
rect 31726 4196 31754 4236
rect 40052 4236 41368 4264
rect 40052 4205 40080 4236
rect 40037 4199 40095 4205
rect 40037 4196 40049 4199
rect 25700 4168 25912 4196
rect 31726 4168 40049 4196
rect 23566 4088 23572 4140
rect 23624 4128 23630 4140
rect 25700 4128 25728 4168
rect 23624 4100 25728 4128
rect 23624 4088 23630 4100
rect 25774 4088 25780 4140
rect 25832 4088 25838 4140
rect 25884 4128 25912 4168
rect 40037 4165 40049 4168
rect 40083 4165 40095 4199
rect 40037 4159 40095 4165
rect 40218 4156 40224 4208
rect 40276 4196 40282 4208
rect 40276 4168 40540 4196
rect 40276 4156 40282 4168
rect 38930 4128 38936 4140
rect 25884 4100 38936 4128
rect 38930 4088 38936 4100
rect 38988 4088 38994 4140
rect 40512 4128 40540 4168
rect 40586 4156 40592 4208
rect 40644 4156 40650 4208
rect 40957 4199 41015 4205
rect 40957 4196 40969 4199
rect 40788 4168 40969 4196
rect 40788 4128 40816 4168
rect 40957 4165 40969 4168
rect 41003 4196 41015 4199
rect 41230 4196 41236 4208
rect 41003 4168 41236 4196
rect 41003 4165 41015 4168
rect 40957 4159 41015 4165
rect 41230 4156 41236 4168
rect 41288 4156 41294 4208
rect 41340 4205 41368 4236
rect 42886 4224 42892 4276
rect 42944 4264 42950 4276
rect 48590 4264 48596 4276
rect 42944 4236 48596 4264
rect 42944 4224 42950 4236
rect 48590 4224 48596 4236
rect 48648 4224 48654 4276
rect 49050 4224 49056 4276
rect 49108 4264 49114 4276
rect 50065 4267 50123 4273
rect 50065 4264 50077 4267
rect 49108 4236 50077 4264
rect 49108 4224 49114 4236
rect 50065 4233 50077 4236
rect 50111 4233 50123 4267
rect 50065 4227 50123 4233
rect 50249 4267 50307 4273
rect 50249 4233 50261 4267
rect 50295 4264 50307 4267
rect 51166 4264 51172 4276
rect 50295 4236 51172 4264
rect 50295 4233 50307 4236
rect 50249 4227 50307 4233
rect 51166 4224 51172 4236
rect 51224 4224 51230 4276
rect 53374 4224 53380 4276
rect 53432 4264 53438 4276
rect 53432 4236 84194 4264
rect 53432 4224 53438 4236
rect 41325 4199 41383 4205
rect 41325 4165 41337 4199
rect 41371 4165 41383 4199
rect 41693 4199 41751 4205
rect 41693 4196 41705 4199
rect 41325 4159 41383 4165
rect 41432 4168 41705 4196
rect 40512 4100 40816 4128
rect 40862 4088 40868 4140
rect 40920 4088 40926 4140
rect 41046 4088 41052 4140
rect 41104 4128 41110 4140
rect 41432 4128 41460 4168
rect 41693 4165 41705 4168
rect 41739 4165 41751 4199
rect 41693 4159 41751 4165
rect 42610 4156 42616 4208
rect 42668 4196 42674 4208
rect 42668 4168 45508 4196
rect 42668 4156 42674 4168
rect 41104 4100 41460 4128
rect 45480 4128 45508 4168
rect 48038 4156 48044 4208
rect 48096 4196 48102 4208
rect 48133 4199 48191 4205
rect 48133 4196 48145 4199
rect 48096 4168 48145 4196
rect 48096 4156 48102 4168
rect 48133 4165 48145 4168
rect 48179 4165 48191 4199
rect 48133 4159 48191 4165
rect 48961 4199 49019 4205
rect 48961 4165 48973 4199
rect 49007 4196 49019 4199
rect 49142 4196 49148 4208
rect 49007 4168 49148 4196
rect 49007 4165 49019 4168
rect 48961 4159 49019 4165
rect 49142 4156 49148 4168
rect 49200 4156 49206 4208
rect 49234 4156 49240 4208
rect 49292 4156 49298 4208
rect 49326 4156 49332 4208
rect 49384 4156 49390 4208
rect 49697 4199 49755 4205
rect 49697 4165 49709 4199
rect 49743 4196 49755 4199
rect 49878 4196 49884 4208
rect 49743 4168 49884 4196
rect 49743 4165 49755 4168
rect 49697 4159 49755 4165
rect 49878 4156 49884 4168
rect 49936 4156 49942 4208
rect 50985 4199 51043 4205
rect 50985 4165 50997 4199
rect 51031 4196 51043 4199
rect 51534 4196 51540 4208
rect 51031 4168 51540 4196
rect 51031 4165 51043 4168
rect 50985 4159 51043 4165
rect 51534 4156 51540 4168
rect 51592 4156 51598 4208
rect 51718 4156 51724 4208
rect 51776 4156 51782 4208
rect 51810 4156 51816 4208
rect 51868 4196 51874 4208
rect 52089 4199 52147 4205
rect 52089 4196 52101 4199
rect 51868 4168 52101 4196
rect 51868 4156 51874 4168
rect 52089 4165 52101 4168
rect 52135 4165 52147 4199
rect 52089 4159 52147 4165
rect 53009 4199 53067 4205
rect 53009 4165 53021 4199
rect 53055 4196 53067 4199
rect 80882 4196 80888 4208
rect 53055 4168 80888 4196
rect 53055 4165 53067 4168
rect 53009 4159 53067 4165
rect 80882 4156 80888 4168
rect 80940 4156 80946 4208
rect 81618 4156 81624 4208
rect 81676 4196 81682 4208
rect 83642 4196 83648 4208
rect 81676 4168 83648 4196
rect 81676 4156 81682 4168
rect 83642 4156 83648 4168
rect 83700 4156 83706 4208
rect 47857 4131 47915 4137
rect 47857 4128 47869 4131
rect 45480 4100 47869 4128
rect 41104 4088 41110 4100
rect 47857 4097 47869 4100
rect 47903 4128 47915 4131
rect 47903 4100 49832 4128
rect 47903 4097 47915 4100
rect 47857 4091 47915 4097
rect 49804 4072 49832 4100
rect 51258 4088 51264 4140
rect 51316 4088 51322 4140
rect 51350 4088 51356 4140
rect 51408 4128 51414 4140
rect 52454 4128 52460 4140
rect 51408 4100 52460 4128
rect 51408 4088 51414 4100
rect 52454 4088 52460 4100
rect 52512 4128 52518 4140
rect 53193 4131 53251 4137
rect 53193 4128 53205 4131
rect 52512 4100 53205 4128
rect 52512 4088 52518 4100
rect 53193 4097 53205 4100
rect 53239 4097 53251 4131
rect 84166 4128 84194 4236
rect 87506 4224 87512 4276
rect 87564 4264 87570 4276
rect 112990 4264 112996 4276
rect 87564 4236 112996 4264
rect 87564 4224 87570 4236
rect 112990 4224 112996 4236
rect 113048 4224 113054 4276
rect 113174 4224 113180 4276
rect 113232 4264 113238 4276
rect 123386 4264 123392 4276
rect 113232 4236 123392 4264
rect 113232 4224 113238 4236
rect 123386 4224 123392 4236
rect 123444 4224 123450 4276
rect 142430 4264 142436 4276
rect 123588 4236 142436 4264
rect 84930 4156 84936 4208
rect 84988 4156 84994 4208
rect 96062 4156 96068 4208
rect 96120 4196 96126 4208
rect 102042 4196 102048 4208
rect 96120 4168 102048 4196
rect 96120 4156 96126 4168
rect 102042 4156 102048 4168
rect 102100 4156 102106 4208
rect 109862 4156 109868 4208
rect 109920 4196 109926 4208
rect 112530 4196 112536 4208
rect 109920 4168 112536 4196
rect 109920 4156 109926 4168
rect 112530 4156 112536 4168
rect 112588 4156 112594 4208
rect 116394 4156 116400 4208
rect 116452 4196 116458 4208
rect 116452 4168 123340 4196
rect 116452 4156 116458 4168
rect 84749 4131 84807 4137
rect 84749 4128 84761 4131
rect 84166 4100 84761 4128
rect 53193 4091 53251 4097
rect 84749 4097 84761 4100
rect 84795 4097 84807 4131
rect 84749 4091 84807 4097
rect 86589 4131 86647 4137
rect 86589 4097 86601 4131
rect 86635 4128 86647 4131
rect 86957 4131 87015 4137
rect 86957 4128 86969 4131
rect 86635 4100 86969 4128
rect 86635 4097 86647 4100
rect 86589 4091 86647 4097
rect 86957 4097 86969 4100
rect 87003 4128 87015 4131
rect 91002 4128 91008 4140
rect 87003 4100 91008 4128
rect 87003 4097 87015 4100
rect 86957 4091 87015 4097
rect 14366 4020 14372 4072
rect 14424 4060 14430 4072
rect 14424 4032 36676 4060
rect 14424 4020 14430 4032
rect 9214 3952 9220 4004
rect 9272 3992 9278 4004
rect 36538 3992 36544 4004
rect 9272 3964 36544 3992
rect 9272 3952 9278 3964
rect 36538 3952 36544 3964
rect 36596 3952 36602 4004
rect 24486 3884 24492 3936
rect 24544 3924 24550 3936
rect 25961 3927 26019 3933
rect 25961 3924 25973 3927
rect 24544 3896 25973 3924
rect 24544 3884 24550 3896
rect 25961 3893 25973 3896
rect 26007 3893 26019 3927
rect 36648 3924 36676 4032
rect 40770 4020 40776 4072
rect 40828 4020 40834 4072
rect 49786 4020 49792 4072
rect 49844 4020 49850 4072
rect 51626 4020 51632 4072
rect 51684 4020 51690 4072
rect 81434 4020 81440 4072
rect 81492 4020 81498 4072
rect 83277 4063 83335 4069
rect 83277 4029 83289 4063
rect 83323 4060 83335 4063
rect 83323 4032 83964 4060
rect 83323 4029 83335 4032
rect 83277 4023 83335 4029
rect 80793 3995 80851 4001
rect 80793 3961 80805 3995
rect 80839 3992 80851 3995
rect 81161 3995 81219 4001
rect 81161 3992 81173 3995
rect 80839 3964 81173 3992
rect 80839 3961 80851 3964
rect 80793 3955 80851 3961
rect 81161 3961 81173 3964
rect 81207 3992 81219 3995
rect 83292 3992 83320 4023
rect 81207 3964 83320 3992
rect 81207 3961 81219 3964
rect 81161 3955 81219 3961
rect 83936 3936 83964 4032
rect 84473 3995 84531 4001
rect 84473 3961 84485 3995
rect 84519 3992 84531 3995
rect 86604 3992 86632 4091
rect 91002 4088 91008 4100
rect 91060 4088 91066 4140
rect 94314 4088 94320 4140
rect 94372 4088 94378 4140
rect 104897 4131 104955 4137
rect 104897 4097 104909 4131
rect 104943 4128 104955 4131
rect 104986 4128 104992 4140
rect 104943 4100 104992 4128
rect 104943 4097 104955 4100
rect 104897 4091 104955 4097
rect 104986 4088 104992 4100
rect 105044 4088 105050 4140
rect 105814 4088 105820 4140
rect 105872 4088 105878 4140
rect 106734 4088 106740 4140
rect 106792 4128 106798 4140
rect 107197 4131 107255 4137
rect 107197 4128 107209 4131
rect 106792 4100 107209 4128
rect 106792 4088 106798 4100
rect 107197 4097 107209 4100
rect 107243 4097 107255 4131
rect 107197 4091 107255 4097
rect 108390 4088 108396 4140
rect 108448 4088 108454 4140
rect 112346 4088 112352 4140
rect 112404 4088 112410 4140
rect 113542 4088 113548 4140
rect 113600 4088 113606 4140
rect 114186 4088 114192 4140
rect 114244 4088 114250 4140
rect 114649 4131 114707 4137
rect 114649 4097 114661 4131
rect 114695 4128 114707 4131
rect 114738 4128 114744 4140
rect 114695 4100 114744 4128
rect 114695 4097 114707 4100
rect 114649 4091 114707 4097
rect 114738 4088 114744 4100
rect 114796 4088 114802 4140
rect 115566 4088 115572 4140
rect 115624 4088 115630 4140
rect 123312 4128 123340 4168
rect 123588 4128 123616 4236
rect 142430 4224 142436 4236
rect 142488 4224 142494 4276
rect 151078 4224 151084 4276
rect 151136 4264 151142 4276
rect 154390 4264 154396 4276
rect 151136 4236 154396 4264
rect 151136 4224 151142 4236
rect 154390 4224 154396 4236
rect 154448 4224 154454 4276
rect 213914 4264 213920 4276
rect 157306 4236 213920 4264
rect 123662 4156 123668 4208
rect 123720 4196 123726 4208
rect 147490 4196 147496 4208
rect 123720 4168 147496 4196
rect 123720 4156 123726 4168
rect 145024 4137 145052 4168
rect 147490 4156 147496 4168
rect 147548 4156 147554 4208
rect 148410 4196 148416 4208
rect 147646 4168 148416 4196
rect 123312 4100 123616 4128
rect 145009 4131 145067 4137
rect 145009 4097 145021 4131
rect 145055 4097 145067 4131
rect 147646 4128 147674 4168
rect 148410 4156 148416 4168
rect 148468 4196 148474 4208
rect 148870 4196 148876 4208
rect 148468 4168 148876 4196
rect 148468 4156 148474 4168
rect 148870 4156 148876 4168
rect 148928 4196 148934 4208
rect 151814 4196 151820 4208
rect 148928 4168 151820 4196
rect 148928 4156 148934 4168
rect 151814 4156 151820 4168
rect 151872 4156 151878 4208
rect 154666 4156 154672 4208
rect 154724 4196 154730 4208
rect 157306 4196 157334 4236
rect 213914 4224 213920 4236
rect 213972 4224 213978 4276
rect 215110 4224 215116 4276
rect 215168 4264 215174 4276
rect 216769 4267 216827 4273
rect 216769 4264 216781 4267
rect 215168 4236 216781 4264
rect 215168 4224 215174 4236
rect 216769 4233 216781 4236
rect 216815 4233 216827 4267
rect 216769 4227 216827 4233
rect 219066 4224 219072 4276
rect 219124 4264 219130 4276
rect 222010 4264 222016 4276
rect 219124 4236 222016 4264
rect 219124 4224 219130 4236
rect 222010 4224 222016 4236
rect 222068 4224 222074 4276
rect 240042 4264 240048 4276
rect 222212 4236 240048 4264
rect 154724 4168 157334 4196
rect 154724 4156 154730 4168
rect 157794 4156 157800 4208
rect 157852 4196 157858 4208
rect 158073 4199 158131 4205
rect 158073 4196 158085 4199
rect 157852 4168 158085 4196
rect 157852 4156 157858 4168
rect 158073 4165 158085 4168
rect 158119 4165 158131 4199
rect 158073 4159 158131 4165
rect 161290 4156 161296 4208
rect 161348 4156 161354 4208
rect 189994 4156 190000 4208
rect 190052 4156 190058 4208
rect 209682 4156 209688 4208
rect 209740 4196 209746 4208
rect 209740 4168 209820 4196
rect 209740 4156 209746 4168
rect 145009 4091 145067 4097
rect 147416 4100 147674 4128
rect 93762 4020 93768 4072
rect 93820 4060 93826 4072
rect 94501 4063 94559 4069
rect 94501 4060 94513 4063
rect 93820 4032 94513 4060
rect 93820 4020 93826 4032
rect 94501 4029 94513 4032
rect 94547 4029 94559 4063
rect 94501 4023 94559 4029
rect 96154 4020 96160 4072
rect 96212 4020 96218 4072
rect 98546 4020 98552 4072
rect 98604 4060 98610 4072
rect 99377 4063 99435 4069
rect 99377 4060 99389 4063
rect 98604 4032 99389 4060
rect 98604 4020 98610 4032
rect 99377 4029 99389 4032
rect 99423 4029 99435 4063
rect 99377 4023 99435 4029
rect 99561 4063 99619 4069
rect 99561 4029 99573 4063
rect 99607 4060 99619 4063
rect 99742 4060 99748 4072
rect 99607 4032 99748 4060
rect 99607 4029 99619 4032
rect 99561 4023 99619 4029
rect 99742 4020 99748 4032
rect 99800 4020 99806 4072
rect 101217 4063 101275 4069
rect 101217 4029 101229 4063
rect 101263 4029 101275 4063
rect 101217 4023 101275 4029
rect 84519 3964 86632 3992
rect 84519 3961 84531 3964
rect 84473 3955 84531 3961
rect 92290 3952 92296 4004
rect 92348 3992 92354 4004
rect 98914 3992 98920 4004
rect 92348 3964 98920 3992
rect 92348 3952 92354 3964
rect 98914 3952 98920 3964
rect 98972 3952 98978 4004
rect 40402 3924 40408 3936
rect 36648 3896 40408 3924
rect 25961 3887 26019 3893
rect 40402 3884 40408 3896
rect 40460 3884 40466 3936
rect 41874 3884 41880 3936
rect 41932 3884 41938 3936
rect 42794 3884 42800 3936
rect 42852 3924 42858 3936
rect 47394 3924 47400 3936
rect 42852 3896 47400 3924
rect 42852 3884 42858 3896
rect 47394 3884 47400 3896
rect 47452 3884 47458 3936
rect 52270 3884 52276 3936
rect 52328 3884 52334 3936
rect 83918 3884 83924 3936
rect 83976 3884 83982 3936
rect 87690 3884 87696 3936
rect 87748 3924 87754 3936
rect 96890 3924 96896 3936
rect 87748 3896 96896 3924
rect 87748 3884 87754 3896
rect 96890 3884 96896 3896
rect 96948 3884 96954 3936
rect 98178 3884 98184 3936
rect 98236 3924 98242 3936
rect 98641 3927 98699 3933
rect 98641 3924 98653 3927
rect 98236 3896 98653 3924
rect 98236 3884 98242 3896
rect 98641 3893 98653 3896
rect 98687 3924 98699 3927
rect 101232 3924 101260 4023
rect 102226 4020 102232 4072
rect 102284 4060 102290 4072
rect 102284 4032 104756 4060
rect 102284 4020 102290 4032
rect 102870 3952 102876 4004
rect 102928 3992 102934 4004
rect 104728 3992 104756 4032
rect 105078 4020 105084 4072
rect 105136 4020 105142 4072
rect 105538 4020 105544 4072
rect 105596 4020 105602 4072
rect 105998 4069 106004 4072
rect 105955 4063 106004 4069
rect 105955 4029 105967 4063
rect 106001 4029 106004 4063
rect 105955 4023 106004 4029
rect 105998 4020 106004 4023
rect 106056 4020 106062 4072
rect 106093 4063 106151 4069
rect 106093 4029 106105 4063
rect 106139 4060 106151 4063
rect 107286 4060 107292 4072
rect 106139 4032 107292 4060
rect 106139 4029 106151 4032
rect 106093 4023 106151 4029
rect 105556 3992 105584 4020
rect 102928 3964 104664 3992
rect 104728 3964 105584 3992
rect 102928 3952 102934 3964
rect 101582 3924 101588 3936
rect 98687 3896 101588 3924
rect 98687 3893 98699 3896
rect 98641 3887 98699 3893
rect 101582 3884 101588 3896
rect 101640 3884 101646 3936
rect 104069 3927 104127 3933
rect 104069 3893 104081 3927
rect 104115 3924 104127 3927
rect 104526 3924 104532 3936
rect 104115 3896 104532 3924
rect 104115 3893 104127 3896
rect 104069 3887 104127 3893
rect 104526 3884 104532 3896
rect 104584 3884 104590 3936
rect 104636 3924 104664 3964
rect 106476 3924 106504 4032
rect 107286 4020 107292 4032
rect 107344 4020 107350 4072
rect 107378 4020 107384 4072
rect 107436 4020 107442 4072
rect 108117 4063 108175 4069
rect 108117 4060 108129 4063
rect 107948 4032 108129 4060
rect 106918 3952 106924 4004
rect 106976 3992 106982 4004
rect 107746 3992 107752 4004
rect 106976 3964 107752 3992
rect 106976 3952 106982 3964
rect 107746 3952 107752 3964
rect 107804 3992 107810 4004
rect 107841 3995 107899 4001
rect 107841 3992 107853 3995
rect 107804 3964 107853 3992
rect 107804 3952 107810 3964
rect 107841 3961 107853 3964
rect 107887 3961 107899 3995
rect 107841 3955 107899 3961
rect 104636 3896 106504 3924
rect 106737 3927 106795 3933
rect 106737 3893 106749 3927
rect 106783 3924 106795 3927
rect 107102 3924 107108 3936
rect 106783 3896 107108 3924
rect 106783 3893 106795 3896
rect 106737 3887 106795 3893
rect 107102 3884 107108 3896
rect 107160 3884 107166 3936
rect 107948 3924 107976 4032
rect 108117 4029 108129 4032
rect 108163 4029 108175 4063
rect 108117 4023 108175 4029
rect 108255 4063 108313 4069
rect 108255 4029 108267 4063
rect 108301 4060 108313 4063
rect 111334 4060 111340 4072
rect 108301 4032 111340 4060
rect 108301 4029 108313 4032
rect 108255 4023 108313 4029
rect 111334 4020 111340 4032
rect 111392 4020 111398 4072
rect 112530 4020 112536 4072
rect 112588 4020 112594 4072
rect 113450 4069 113456 4072
rect 113269 4063 113327 4069
rect 113269 4060 113281 4063
rect 113100 4032 113281 4060
rect 112438 3952 112444 4004
rect 112496 3992 112502 4004
rect 112990 3992 112996 4004
rect 112496 3964 112996 3992
rect 112496 3952 112502 3964
rect 112990 3952 112996 3964
rect 113048 3952 113054 4004
rect 108942 3924 108948 3936
rect 107948 3896 108948 3924
rect 108942 3884 108948 3896
rect 109000 3884 109006 3936
rect 109037 3927 109095 3933
rect 109037 3893 109049 3927
rect 109083 3924 109095 3927
rect 110230 3924 110236 3936
rect 109083 3896 110236 3924
rect 109083 3893 109095 3896
rect 109037 3887 109095 3893
rect 110230 3884 110236 3896
rect 110288 3884 110294 3936
rect 113100 3924 113128 4032
rect 113269 4029 113281 4032
rect 113315 4029 113327 4063
rect 113269 4023 113327 4029
rect 113407 4063 113456 4069
rect 113407 4029 113419 4063
rect 113453 4029 113456 4063
rect 113407 4023 113456 4029
rect 113450 4020 113456 4023
rect 113508 4020 113514 4072
rect 114830 4020 114836 4072
rect 114888 4020 114894 4072
rect 115686 4063 115744 4069
rect 115686 4060 115698 4063
rect 115400 4032 115698 4060
rect 115290 3952 115296 4004
rect 115348 3952 115354 4004
rect 114554 3924 114560 3936
rect 113100 3896 114560 3924
rect 114554 3884 114560 3896
rect 114612 3884 114618 3936
rect 115400 3924 115428 4032
rect 115686 4029 115698 4032
rect 115732 4029 115744 4063
rect 115686 4023 115744 4029
rect 115845 4063 115903 4069
rect 115845 4029 115857 4063
rect 115891 4060 115903 4063
rect 116026 4060 116032 4072
rect 115891 4032 116032 4060
rect 115891 4029 115903 4032
rect 115845 4023 115903 4029
rect 116026 4020 116032 4032
rect 116084 4020 116090 4072
rect 116762 4020 116768 4072
rect 116820 4060 116826 4072
rect 117501 4063 117559 4069
rect 117501 4060 117513 4063
rect 116820 4032 117513 4060
rect 116820 4020 116826 4032
rect 117501 4029 117513 4032
rect 117547 4029 117559 4063
rect 117501 4023 117559 4029
rect 117682 4020 117688 4072
rect 117740 4020 117746 4072
rect 117961 4063 118019 4069
rect 117961 4029 117973 4063
rect 118007 4029 118019 4063
rect 117961 4023 118019 4029
rect 117976 3992 118004 4023
rect 120994 4020 121000 4072
rect 121052 4060 121058 4072
rect 121733 4063 121791 4069
rect 121733 4060 121745 4063
rect 121052 4032 121745 4060
rect 121052 4020 121058 4032
rect 121733 4029 121745 4032
rect 121779 4029 121791 4063
rect 121733 4023 121791 4029
rect 121914 4020 121920 4072
rect 121972 4060 121978 4072
rect 122650 4060 122656 4072
rect 121972 4032 122656 4060
rect 121972 4020 121978 4032
rect 122650 4020 122656 4032
rect 122708 4020 122714 4072
rect 123573 4063 123631 4069
rect 123573 4029 123585 4063
rect 123619 4060 123631 4063
rect 123619 4032 123984 4060
rect 123619 4029 123631 4032
rect 123573 4023 123631 4029
rect 117148 3964 118694 3992
rect 116394 3924 116400 3936
rect 115400 3896 116400 3924
rect 116394 3884 116400 3896
rect 116452 3884 116458 3936
rect 116486 3884 116492 3936
rect 116544 3884 116550 3936
rect 116670 3884 116676 3936
rect 116728 3924 116734 3936
rect 117148 3933 117176 3964
rect 116765 3927 116823 3933
rect 116765 3924 116777 3927
rect 116728 3896 116777 3924
rect 116728 3884 116734 3896
rect 116765 3893 116777 3896
rect 116811 3924 116823 3927
rect 117133 3927 117191 3933
rect 117133 3924 117145 3927
rect 116811 3896 117145 3924
rect 116811 3893 116823 3896
rect 116765 3887 116823 3893
rect 117133 3893 117145 3896
rect 117179 3893 117191 3927
rect 118666 3924 118694 3964
rect 120902 3952 120908 4004
rect 120960 3992 120966 4004
rect 121089 3995 121147 4001
rect 121089 3992 121101 3995
rect 120960 3964 121101 3992
rect 120960 3952 120966 3964
rect 121089 3961 121101 3964
rect 121135 3992 121147 3995
rect 121457 3995 121515 4001
rect 121457 3992 121469 3995
rect 121135 3964 121469 3992
rect 121135 3961 121147 3964
rect 121089 3955 121147 3961
rect 121457 3961 121469 3964
rect 121503 3992 121515 3995
rect 123588 3992 123616 4023
rect 121503 3964 123616 3992
rect 121503 3961 121515 3964
rect 121457 3955 121515 3961
rect 119982 3924 119988 3936
rect 118666 3896 119988 3924
rect 117133 3887 117191 3893
rect 119982 3884 119988 3896
rect 120040 3884 120046 3936
rect 123956 3933 123984 4032
rect 124306 4020 124312 4072
rect 124364 4060 124370 4072
rect 139302 4060 139308 4072
rect 124364 4032 139308 4060
rect 124364 4020 124370 4032
rect 139302 4020 139308 4032
rect 139360 4020 139366 4072
rect 141786 4020 141792 4072
rect 141844 4020 141850 4072
rect 141973 4063 142031 4069
rect 141973 4029 141985 4063
rect 142019 4060 142031 4063
rect 142154 4060 142160 4072
rect 142019 4032 142160 4060
rect 142019 4029 142031 4032
rect 141973 4023 142031 4029
rect 142154 4020 142160 4032
rect 142212 4020 142218 4072
rect 142249 4063 142307 4069
rect 142249 4029 142261 4063
rect 142295 4029 142307 4063
rect 142249 4023 142307 4029
rect 142264 3992 142292 4023
rect 145650 4020 145656 4072
rect 145708 4020 145714 4072
rect 145837 4063 145895 4069
rect 145837 4029 145849 4063
rect 145883 4060 145895 4063
rect 147416 4060 147444 4100
rect 150894 4088 150900 4140
rect 150952 4128 150958 4140
rect 151909 4131 151967 4137
rect 151909 4128 151921 4131
rect 150952 4100 151921 4128
rect 150952 4088 150958 4100
rect 151909 4097 151921 4100
rect 151955 4097 151967 4131
rect 151909 4091 151967 4097
rect 152642 4088 152648 4140
rect 152700 4088 152706 4140
rect 154482 4088 154488 4140
rect 154540 4128 154546 4140
rect 154577 4131 154635 4137
rect 154577 4128 154589 4131
rect 154540 4100 154589 4128
rect 154540 4088 154546 4100
rect 154577 4097 154589 4100
rect 154623 4097 154635 4131
rect 155678 4128 155684 4140
rect 154577 4091 154635 4097
rect 154684 4100 155684 4128
rect 145883 4032 147444 4060
rect 145883 4029 145895 4032
rect 145837 4023 145895 4029
rect 147950 4020 147956 4072
rect 148008 4020 148014 4072
rect 148134 4020 148140 4072
rect 148192 4020 148198 4072
rect 149054 4020 149060 4072
rect 149112 4060 149118 4072
rect 149790 4060 149796 4072
rect 149112 4032 149796 4060
rect 149112 4020 149118 4032
rect 149790 4020 149796 4032
rect 149848 4020 149854 4072
rect 151262 4020 151268 4072
rect 151320 4060 151326 4072
rect 151725 4063 151783 4069
rect 151725 4060 151737 4063
rect 151320 4032 151737 4060
rect 151320 4020 151326 4032
rect 151725 4029 151737 4032
rect 151771 4029 151783 4063
rect 151725 4023 151783 4029
rect 152369 4063 152427 4069
rect 152369 4029 152381 4063
rect 152415 4060 152427 4063
rect 152458 4060 152464 4072
rect 152415 4032 152464 4060
rect 152415 4029 152427 4032
rect 152369 4023 152427 4029
rect 152458 4020 152464 4032
rect 152516 4020 152522 4072
rect 152826 4069 152832 4072
rect 152783 4063 152832 4069
rect 152783 4029 152795 4063
rect 152829 4029 152832 4063
rect 152783 4023 152832 4029
rect 152826 4020 152832 4023
rect 152884 4020 152890 4072
rect 152918 4020 152924 4072
rect 152976 4020 152982 4072
rect 153565 4063 153623 4069
rect 153565 4029 153577 4063
rect 153611 4060 153623 4063
rect 154684 4060 154712 4100
rect 155678 4088 155684 4100
rect 155736 4088 155742 4140
rect 156322 4128 156328 4140
rect 155788 4100 156328 4128
rect 153611 4032 154712 4060
rect 153611 4029 153623 4032
rect 153565 4023 153623 4029
rect 154850 4020 154856 4072
rect 154908 4060 154914 4072
rect 155788 4060 155816 4100
rect 156322 4088 156328 4100
rect 156380 4088 156386 4140
rect 158441 4131 158499 4137
rect 158441 4128 158453 4131
rect 157306 4100 158453 4128
rect 154908 4032 155816 4060
rect 154908 4020 154914 4032
rect 156230 4020 156236 4072
rect 156288 4060 156294 4072
rect 157306 4060 157334 4100
rect 158441 4097 158453 4100
rect 158487 4097 158499 4131
rect 158441 4091 158499 4097
rect 159174 4088 159180 4140
rect 159232 4088 159238 4140
rect 159450 4088 159456 4140
rect 159508 4088 159514 4140
rect 160738 4128 160744 4140
rect 160020 4100 160744 4128
rect 156288 4032 157334 4060
rect 156288 4020 156294 4032
rect 157702 4020 157708 4072
rect 157760 4060 157766 4072
rect 158257 4063 158315 4069
rect 158257 4060 158269 4063
rect 157760 4032 158269 4060
rect 157760 4020 157766 4032
rect 158257 4029 158269 4032
rect 158303 4029 158315 4063
rect 158257 4023 158315 4029
rect 158622 4020 158628 4072
rect 158680 4060 158686 4072
rect 158901 4063 158959 4069
rect 158901 4060 158913 4063
rect 158680 4032 158913 4060
rect 158680 4020 158686 4032
rect 158901 4029 158913 4032
rect 158947 4029 158959 4063
rect 158901 4023 158959 4029
rect 159315 4063 159373 4069
rect 159315 4029 159327 4063
rect 159361 4060 159373 4063
rect 160020 4060 160048 4100
rect 160738 4088 160744 4100
rect 160796 4088 160802 4140
rect 162486 4088 162492 4140
rect 162544 4128 162550 4140
rect 190365 4131 190423 4137
rect 162544 4100 166994 4128
rect 162544 4088 162550 4100
rect 159361 4032 160048 4060
rect 160097 4063 160155 4069
rect 159361 4029 159373 4032
rect 159315 4023 159373 4029
rect 160097 4029 160109 4063
rect 160143 4060 160155 4063
rect 161109 4063 161167 4069
rect 161109 4060 161121 4063
rect 160143 4032 161121 4060
rect 160143 4029 160155 4032
rect 160097 4023 160155 4029
rect 161109 4029 161121 4032
rect 161155 4029 161167 4063
rect 161109 4023 161167 4029
rect 161382 4020 161388 4072
rect 161440 4060 161446 4072
rect 162949 4063 163007 4069
rect 162949 4060 162961 4063
rect 161440 4032 162961 4060
rect 161440 4020 161446 4032
rect 162949 4029 162961 4032
rect 162995 4060 163007 4063
rect 163317 4063 163375 4069
rect 163317 4060 163329 4063
rect 162995 4032 163329 4060
rect 162995 4029 163007 4032
rect 162949 4023 163007 4029
rect 163317 4029 163329 4032
rect 163363 4060 163375 4063
rect 163682 4060 163688 4072
rect 163363 4032 163688 4060
rect 163363 4029 163375 4032
rect 163317 4023 163375 4029
rect 163682 4020 163688 4032
rect 163740 4020 163746 4072
rect 166966 4060 166994 4100
rect 190365 4097 190377 4131
rect 190411 4128 190423 4131
rect 190914 4128 190920 4140
rect 190411 4100 190920 4128
rect 190411 4097 190423 4100
rect 190365 4091 190423 4097
rect 190914 4088 190920 4100
rect 190972 4088 190978 4140
rect 209314 4088 209320 4140
rect 209372 4088 209378 4140
rect 209792 4137 209820 4168
rect 216858 4156 216864 4208
rect 216916 4196 216922 4208
rect 216916 4168 219480 4196
rect 216916 4156 216922 4168
rect 209777 4131 209835 4137
rect 209777 4097 209789 4131
rect 209823 4097 209835 4131
rect 209777 4091 209835 4097
rect 212626 4088 212632 4140
rect 212684 4128 212690 4140
rect 212813 4131 212871 4137
rect 212813 4128 212825 4131
rect 212684 4100 212825 4128
rect 212684 4088 212690 4100
rect 212813 4097 212825 4100
rect 212859 4097 212871 4131
rect 212813 4091 212871 4097
rect 214006 4088 214012 4140
rect 214064 4088 214070 4140
rect 214926 4088 214932 4140
rect 214984 4088 214990 4140
rect 215846 4088 215852 4140
rect 215904 4088 215910 4140
rect 216122 4088 216128 4140
rect 216180 4088 216186 4140
rect 219452 4128 219480 4168
rect 222212 4128 222240 4236
rect 240042 4224 240048 4236
rect 240100 4224 240106 4276
rect 242986 4264 242992 4276
rect 240520 4236 242992 4264
rect 226610 4156 226616 4208
rect 226668 4196 226674 4208
rect 226705 4199 226763 4205
rect 226705 4196 226717 4199
rect 226668 4168 226717 4196
rect 226668 4156 226674 4168
rect 226705 4165 226717 4168
rect 226751 4196 226763 4199
rect 231026 4196 231032 4208
rect 226751 4168 231032 4196
rect 226751 4165 226763 4168
rect 226705 4159 226763 4165
rect 231026 4156 231032 4168
rect 231084 4156 231090 4208
rect 235626 4156 235632 4208
rect 235684 4156 235690 4208
rect 239674 4156 239680 4208
rect 239732 4196 239738 4208
rect 240413 4199 240471 4205
rect 240413 4196 240425 4199
rect 239732 4168 240425 4196
rect 239732 4156 239738 4168
rect 240413 4165 240425 4168
rect 240459 4165 240471 4199
rect 240413 4159 240471 4165
rect 219452 4100 222240 4128
rect 224037 4131 224095 4137
rect 224037 4097 224049 4131
rect 224083 4128 224095 4131
rect 224083 4100 224632 4128
rect 224083 4097 224095 4100
rect 224037 4091 224095 4097
rect 166966 4032 171134 4060
rect 143905 3995 143963 4001
rect 143905 3992 143917 3995
rect 141436 3964 143917 3992
rect 141436 3936 141464 3964
rect 143905 3961 143917 3964
rect 143951 3961 143963 3995
rect 171106 3992 171134 4032
rect 207474 4020 207480 4072
rect 207532 4020 207538 4072
rect 207661 4063 207719 4069
rect 207661 4029 207673 4063
rect 207707 4060 207719 4063
rect 207750 4060 207756 4072
rect 207707 4032 207756 4060
rect 207707 4029 207719 4032
rect 207661 4023 207719 4029
rect 207750 4020 207756 4032
rect 207808 4060 207814 4072
rect 209958 4060 209964 4072
rect 207808 4032 209964 4060
rect 207808 4020 207814 4032
rect 209958 4020 209964 4032
rect 210016 4020 210022 4072
rect 211617 4063 211675 4069
rect 211617 4029 211629 4063
rect 211663 4029 211675 4063
rect 211617 4023 211675 4029
rect 206465 3995 206523 4001
rect 206465 3992 206477 3995
rect 143905 3955 143963 3961
rect 147416 3964 152504 3992
rect 123941 3927 123999 3933
rect 123941 3893 123953 3927
rect 123987 3924 123999 3927
rect 124030 3924 124036 3936
rect 123987 3896 124036 3924
rect 123987 3893 123999 3896
rect 123941 3887 123999 3893
rect 124030 3884 124036 3896
rect 124088 3884 124094 3936
rect 141418 3884 141424 3936
rect 141476 3884 141482 3936
rect 143920 3924 143948 3955
rect 147416 3924 147444 3964
rect 143920 3896 147444 3924
rect 147490 3884 147496 3936
rect 147548 3924 147554 3936
rect 147861 3927 147919 3933
rect 147861 3924 147873 3927
rect 147548 3896 147873 3924
rect 147548 3884 147554 3896
rect 147861 3893 147873 3896
rect 147907 3924 147919 3927
rect 150986 3924 150992 3936
rect 147907 3896 150992 3924
rect 147907 3893 147919 3896
rect 147861 3887 147919 3893
rect 150986 3884 150992 3896
rect 151044 3884 151050 3936
rect 152476 3924 152504 3964
rect 153304 3964 158852 3992
rect 153304 3924 153332 3964
rect 152476 3896 153332 3924
rect 155405 3927 155463 3933
rect 155405 3893 155417 3927
rect 155451 3924 155463 3927
rect 156966 3924 156972 3936
rect 155451 3896 156972 3924
rect 155451 3893 155463 3896
rect 155405 3887 155463 3893
rect 156966 3884 156972 3896
rect 157024 3884 157030 3936
rect 158824 3924 158852 3964
rect 160020 3964 166994 3992
rect 171106 3964 206477 3992
rect 160020 3924 160048 3964
rect 158824 3896 160048 3924
rect 160462 3884 160468 3936
rect 160520 3924 160526 3936
rect 160557 3927 160615 3933
rect 160557 3924 160569 3927
rect 160520 3896 160569 3924
rect 160520 3884 160526 3896
rect 160557 3893 160569 3896
rect 160603 3924 160615 3927
rect 161382 3924 161388 3936
rect 160603 3896 161388 3924
rect 160603 3893 160615 3896
rect 160557 3887 160615 3893
rect 161382 3884 161388 3896
rect 161440 3884 161446 3936
rect 166966 3924 166994 3964
rect 206465 3961 206477 3964
rect 206511 3992 206523 3995
rect 206833 3995 206891 4001
rect 206833 3992 206845 3995
rect 206511 3964 206845 3992
rect 206511 3961 206523 3964
rect 206465 3955 206523 3961
rect 206833 3961 206845 3964
rect 206879 3992 206891 3995
rect 206879 3964 207888 3992
rect 206879 3961 206891 3964
rect 206833 3955 206891 3961
rect 207658 3924 207664 3936
rect 166966 3896 207664 3924
rect 207658 3884 207664 3896
rect 207716 3884 207722 3936
rect 207860 3924 207888 3964
rect 208026 3952 208032 4004
rect 208084 3992 208090 4004
rect 211632 3992 211660 4023
rect 211798 4020 211804 4072
rect 211856 4060 211862 4072
rect 212997 4063 213055 4069
rect 212997 4060 213009 4063
rect 211856 4032 213009 4060
rect 211856 4020 211862 4032
rect 212997 4029 213009 4032
rect 213043 4029 213055 4063
rect 212997 4023 213055 4029
rect 213086 4020 213092 4072
rect 213144 4060 213150 4072
rect 213454 4060 213460 4072
rect 213144 4032 213460 4060
rect 213144 4020 213150 4032
rect 213454 4020 213460 4032
rect 213512 4020 213518 4072
rect 213733 4063 213791 4069
rect 213733 4060 213745 4063
rect 213564 4032 213745 4060
rect 208084 3964 211660 3992
rect 208084 3952 208090 3964
rect 209314 3924 209320 3936
rect 207860 3896 209320 3924
rect 209314 3884 209320 3896
rect 209372 3924 209378 3936
rect 210878 3924 210884 3936
rect 209372 3896 210884 3924
rect 209372 3884 209378 3896
rect 210878 3884 210884 3896
rect 210936 3884 210942 3936
rect 211632 3924 211660 3964
rect 211985 3927 212043 3933
rect 211985 3924 211997 3927
rect 211632 3896 211997 3924
rect 211985 3893 211997 3896
rect 212031 3924 212043 3927
rect 212721 3927 212779 3933
rect 212721 3924 212733 3927
rect 212031 3896 212733 3924
rect 212031 3893 212043 3896
rect 211985 3887 212043 3893
rect 212721 3893 212733 3896
rect 212767 3924 212779 3927
rect 213270 3924 213276 3936
rect 212767 3896 213276 3924
rect 212767 3893 212779 3896
rect 212721 3887 212779 3893
rect 213270 3884 213276 3896
rect 213328 3884 213334 3936
rect 213564 3924 213592 4032
rect 213733 4029 213745 4032
rect 213779 4029 213791 4063
rect 213733 4023 213791 4029
rect 213822 4020 213828 4072
rect 213880 4069 213886 4072
rect 213880 4063 213908 4069
rect 213896 4029 213908 4063
rect 213880 4023 213908 4029
rect 213880 4020 213886 4023
rect 214190 4020 214196 4072
rect 214248 4060 214254 4072
rect 215113 4063 215171 4069
rect 215113 4060 215125 4063
rect 214248 4032 215125 4060
rect 214248 4020 214254 4032
rect 215113 4029 215125 4032
rect 215159 4029 215171 4063
rect 215113 4023 215171 4029
rect 215478 4020 215484 4072
rect 215536 4060 215542 4072
rect 215573 4063 215631 4069
rect 215573 4060 215585 4063
rect 215536 4032 215585 4060
rect 215536 4020 215542 4032
rect 215573 4029 215585 4032
rect 215619 4029 215631 4063
rect 215573 4023 215631 4029
rect 215987 4063 216045 4069
rect 215987 4029 215999 4063
rect 216033 4060 216045 4063
rect 221642 4060 221648 4072
rect 216033 4032 221648 4060
rect 216033 4029 216045 4032
rect 215987 4023 216045 4029
rect 221642 4020 221648 4032
rect 221700 4020 221706 4072
rect 222930 4020 222936 4072
rect 222988 4060 222994 4072
rect 224313 4063 224371 4069
rect 224313 4060 224325 4063
rect 222988 4032 224325 4060
rect 222988 4020 222994 4032
rect 224313 4029 224325 4032
rect 224359 4029 224371 4063
rect 224313 4023 224371 4029
rect 224494 4020 224500 4072
rect 224552 4020 224558 4072
rect 224604 4060 224632 4100
rect 226150 4088 226156 4140
rect 226208 4088 226214 4140
rect 229830 4088 229836 4140
rect 229888 4128 229894 4140
rect 230385 4131 230443 4137
rect 230385 4128 230397 4131
rect 229888 4100 230397 4128
rect 229888 4088 229894 4100
rect 230385 4097 230397 4100
rect 230431 4128 230443 4131
rect 231302 4128 231308 4140
rect 230431 4100 231308 4128
rect 230431 4097 230443 4100
rect 230385 4091 230443 4097
rect 231302 4088 231308 4100
rect 231360 4088 231366 4140
rect 236914 4088 236920 4140
rect 236972 4128 236978 4140
rect 240520 4128 240548 4236
rect 242986 4224 242992 4236
rect 243044 4224 243050 4276
rect 245378 4224 245384 4276
rect 245436 4264 245442 4276
rect 264882 4264 264888 4276
rect 245436 4236 264888 4264
rect 245436 4224 245442 4236
rect 264882 4224 264888 4236
rect 264940 4224 264946 4276
rect 265069 4267 265127 4273
rect 265069 4233 265081 4267
rect 265115 4264 265127 4267
rect 265802 4264 265808 4276
rect 265115 4236 265808 4264
rect 265115 4233 265127 4236
rect 265069 4227 265127 4233
rect 265802 4224 265808 4236
rect 265860 4224 265866 4276
rect 266170 4224 266176 4276
rect 266228 4264 266234 4276
rect 268102 4264 268108 4276
rect 266228 4236 268108 4264
rect 266228 4224 266234 4236
rect 268102 4224 268108 4236
rect 268160 4224 268166 4276
rect 268194 4224 268200 4276
rect 268252 4264 268258 4276
rect 268749 4267 268807 4273
rect 268749 4264 268761 4267
rect 268252 4236 268761 4264
rect 268252 4224 268258 4236
rect 268749 4233 268761 4236
rect 268795 4233 268807 4267
rect 268749 4227 268807 4233
rect 241606 4156 241612 4208
rect 241664 4196 241670 4208
rect 242253 4199 242311 4205
rect 242253 4196 242265 4199
rect 241664 4168 242265 4196
rect 241664 4156 241670 4168
rect 242253 4165 242265 4168
rect 242299 4165 242311 4199
rect 242253 4159 242311 4165
rect 243262 4156 243268 4208
rect 243320 4196 243326 4208
rect 243909 4199 243967 4205
rect 243909 4196 243921 4199
rect 243320 4168 243921 4196
rect 243320 4156 243326 4168
rect 243909 4165 243921 4168
rect 243955 4165 243967 4199
rect 243909 4159 243967 4165
rect 251358 4156 251364 4208
rect 251416 4196 251422 4208
rect 252097 4199 252155 4205
rect 252097 4196 252109 4199
rect 251416 4168 252109 4196
rect 251416 4156 251422 4168
rect 252097 4165 252109 4168
rect 252143 4196 252155 4199
rect 254026 4196 254032 4208
rect 252143 4168 254032 4196
rect 252143 4165 252155 4168
rect 252097 4159 252155 4165
rect 254026 4156 254032 4168
rect 254084 4156 254090 4208
rect 255314 4156 255320 4208
rect 255372 4196 255378 4208
rect 255685 4199 255743 4205
rect 255685 4196 255697 4199
rect 255372 4168 255697 4196
rect 255372 4156 255378 4168
rect 255685 4165 255697 4168
rect 255731 4165 255743 4199
rect 255685 4159 255743 4165
rect 257706 4156 257712 4208
rect 257764 4196 257770 4208
rect 259641 4199 259699 4205
rect 259641 4196 259653 4199
rect 257764 4168 259653 4196
rect 257764 4156 257770 4168
rect 259641 4165 259653 4168
rect 259687 4165 259699 4199
rect 259641 4159 259699 4165
rect 260190 4156 260196 4208
rect 260248 4156 260254 4208
rect 260282 4156 260288 4208
rect 260340 4196 260346 4208
rect 260929 4199 260987 4205
rect 260929 4196 260941 4199
rect 260340 4168 260941 4196
rect 260340 4156 260346 4168
rect 260929 4165 260941 4168
rect 260975 4165 260987 4199
rect 264974 4196 264980 4208
rect 260929 4159 260987 4165
rect 264624 4168 264980 4196
rect 236972 4100 240548 4128
rect 236972 4088 236978 4100
rect 240778 4088 240784 4140
rect 240836 4088 240842 4140
rect 254581 4131 254639 4137
rect 254581 4097 254593 4131
rect 254627 4128 254639 4131
rect 260006 4128 260012 4140
rect 254627 4100 260012 4128
rect 254627 4097 254639 4100
rect 254581 4091 254639 4097
rect 260006 4088 260012 4100
rect 260064 4088 260070 4140
rect 264624 4137 264652 4168
rect 264974 4156 264980 4168
rect 265032 4156 265038 4208
rect 268838 4196 268844 4208
rect 265268 4168 268844 4196
rect 265268 4137 265296 4168
rect 268838 4156 268844 4168
rect 268896 4156 268902 4208
rect 271690 4196 271696 4208
rect 269224 4168 271696 4196
rect 264609 4131 264667 4137
rect 264609 4097 264621 4131
rect 264655 4097 264667 4131
rect 264609 4091 264667 4097
rect 265253 4131 265311 4137
rect 265253 4097 265265 4131
rect 265299 4097 265311 4131
rect 265253 4091 265311 4097
rect 265894 4088 265900 4140
rect 265952 4088 265958 4140
rect 266541 4131 266599 4137
rect 266541 4097 266553 4131
rect 266587 4128 266599 4131
rect 267090 4128 267096 4140
rect 266587 4100 267096 4128
rect 266587 4097 266599 4100
rect 266541 4091 266599 4097
rect 267090 4088 267096 4100
rect 267148 4088 267154 4140
rect 267182 4088 267188 4140
rect 267240 4088 267246 4140
rect 267642 4088 267648 4140
rect 267700 4088 267706 4140
rect 268565 4131 268623 4137
rect 268565 4097 268577 4131
rect 268611 4128 268623 4131
rect 268654 4128 268660 4140
rect 268611 4100 268660 4128
rect 268611 4097 268623 4100
rect 268565 4091 268623 4097
rect 268654 4088 268660 4100
rect 268712 4088 268718 4140
rect 269224 4128 269252 4168
rect 271690 4156 271696 4168
rect 271748 4156 271754 4208
rect 268856 4100 269252 4128
rect 269301 4131 269359 4137
rect 268856 4072 268884 4100
rect 269301 4097 269313 4131
rect 269347 4128 269359 4131
rect 269666 4128 269672 4140
rect 269347 4100 269672 4128
rect 269347 4097 269359 4100
rect 269301 4091 269359 4097
rect 269666 4088 269672 4100
rect 269724 4088 269730 4140
rect 270037 4131 270095 4137
rect 270037 4097 270049 4131
rect 270083 4128 270095 4131
rect 270678 4128 270684 4140
rect 270083 4100 270684 4128
rect 270083 4097 270095 4100
rect 270037 4091 270095 4097
rect 270678 4088 270684 4100
rect 270736 4088 270742 4140
rect 270773 4131 270831 4137
rect 270773 4097 270785 4131
rect 270819 4097 270831 4131
rect 270773 4091 270831 4097
rect 225230 4060 225236 4072
rect 224604 4032 225236 4060
rect 225230 4020 225236 4032
rect 225288 4020 225294 4072
rect 225322 4020 225328 4072
rect 225380 4069 225386 4072
rect 225380 4063 225408 4069
rect 225396 4029 225408 4063
rect 225380 4023 225408 4029
rect 225509 4063 225567 4069
rect 225509 4029 225521 4063
rect 225555 4060 225567 4063
rect 225555 4032 226012 4060
rect 225555 4029 225567 4032
rect 225509 4023 225567 4029
rect 225380 4020 225386 4023
rect 214576 3964 215294 3992
rect 214576 3924 214604 3964
rect 213564 3896 214604 3924
rect 214650 3884 214656 3936
rect 214708 3884 214714 3936
rect 215266 3924 215294 3964
rect 216508 3964 222194 3992
rect 216508 3924 216536 3964
rect 215266 3896 216536 3924
rect 216582 3884 216588 3936
rect 216640 3924 216646 3936
rect 218146 3924 218152 3936
rect 216640 3896 218152 3924
rect 216640 3884 216646 3896
rect 218146 3884 218152 3896
rect 218204 3884 218210 3936
rect 222166 3924 222194 3964
rect 224954 3952 224960 4004
rect 225012 3952 225018 4004
rect 225984 3992 226012 4032
rect 226058 4020 226064 4072
rect 226116 4060 226122 4072
rect 226978 4060 226984 4072
rect 226116 4032 226984 4060
rect 226116 4020 226122 4032
rect 226978 4020 226984 4032
rect 227036 4020 227042 4072
rect 227346 4020 227352 4072
rect 227404 4060 227410 4072
rect 228085 4063 228143 4069
rect 228085 4060 228097 4063
rect 227404 4032 228097 4060
rect 227404 4020 227410 4032
rect 228085 4029 228097 4032
rect 228131 4029 228143 4063
rect 228085 4023 228143 4029
rect 228266 4020 228272 4072
rect 228324 4020 228330 4072
rect 229094 4020 229100 4072
rect 229152 4060 229158 4072
rect 230201 4063 230259 4069
rect 230201 4060 230213 4063
rect 229152 4032 230213 4060
rect 229152 4020 229158 4032
rect 230201 4029 230213 4032
rect 230247 4060 230259 4063
rect 230290 4060 230296 4072
rect 230247 4032 230296 4060
rect 230247 4029 230259 4032
rect 230201 4023 230259 4029
rect 230290 4020 230296 4032
rect 230348 4020 230354 4072
rect 230750 4060 230756 4072
rect 230584 4032 230756 4060
rect 226610 3992 226616 4004
rect 225984 3964 226616 3992
rect 226610 3952 226616 3964
rect 226668 3952 226674 4004
rect 230474 3992 230480 4004
rect 226720 3964 230480 3992
rect 226720 3924 226748 3964
rect 230474 3952 230480 3964
rect 230532 3952 230538 4004
rect 230584 4001 230612 4032
rect 230750 4020 230756 4032
rect 230808 4020 230814 4072
rect 237374 4020 237380 4072
rect 237432 4060 237438 4072
rect 251450 4060 251456 4072
rect 237432 4032 251456 4060
rect 237432 4020 237438 4032
rect 251450 4020 251456 4032
rect 251508 4020 251514 4072
rect 252005 4063 252063 4069
rect 252005 4060 252017 4063
rect 251560 4032 252017 4060
rect 230569 3995 230627 4001
rect 230569 3961 230581 3995
rect 230615 3961 230627 3995
rect 230569 3955 230627 3961
rect 230658 3952 230664 4004
rect 230716 3992 230722 4004
rect 235905 3995 235963 4001
rect 230716 3964 235856 3992
rect 230716 3952 230722 3964
rect 222166 3896 226748 3924
rect 226794 3884 226800 3936
rect 226852 3884 226858 3936
rect 226886 3884 226892 3936
rect 226944 3924 226950 3936
rect 227438 3924 227444 3936
rect 226944 3896 227444 3924
rect 226944 3884 226950 3896
rect 227438 3884 227444 3896
rect 227496 3884 227502 3936
rect 231026 3884 231032 3936
rect 231084 3924 231090 3936
rect 235534 3924 235540 3936
rect 231084 3896 235540 3924
rect 231084 3884 231090 3896
rect 235534 3884 235540 3896
rect 235592 3884 235598 3936
rect 235828 3924 235856 3964
rect 235905 3961 235917 3995
rect 235951 3992 235963 3995
rect 243170 3992 243176 4004
rect 235951 3964 243176 3992
rect 235951 3961 235963 3964
rect 235905 3955 235963 3961
rect 243170 3952 243176 3964
rect 243228 3952 243234 4004
rect 244182 3952 244188 4004
rect 244240 3952 244246 4004
rect 242434 3924 242440 3936
rect 235828 3896 242440 3924
rect 242434 3884 242440 3896
rect 242492 3884 242498 3936
rect 242526 3884 242532 3936
rect 242584 3884 242590 3936
rect 242802 3884 242808 3936
rect 242860 3924 242866 3936
rect 251560 3933 251588 4032
rect 252005 4029 252017 4032
rect 252051 4060 252063 4063
rect 252925 4063 252983 4069
rect 252925 4060 252937 4063
rect 252051 4032 252937 4060
rect 252051 4029 252063 4032
rect 252005 4023 252063 4029
rect 252925 4029 252937 4032
rect 252971 4029 252983 4063
rect 252925 4023 252983 4029
rect 253934 4020 253940 4072
rect 253992 4060 253998 4072
rect 253992 4032 254992 4060
rect 253992 4020 253998 4032
rect 254964 4001 254992 4032
rect 256510 4020 256516 4072
rect 256568 4020 256574 4072
rect 256694 4020 256700 4072
rect 256752 4020 256758 4072
rect 257614 4020 257620 4072
rect 257672 4020 257678 4072
rect 257798 4020 257804 4072
rect 257856 4020 257862 4072
rect 258166 4020 258172 4072
rect 258224 4060 258230 4072
rect 259089 4063 259147 4069
rect 259089 4060 259101 4063
rect 258224 4032 259101 4060
rect 258224 4020 258230 4032
rect 259089 4029 259101 4032
rect 259135 4029 259147 4063
rect 259089 4023 259147 4029
rect 261205 4063 261263 4069
rect 261205 4029 261217 4063
rect 261251 4060 261263 4063
rect 265618 4060 265624 4072
rect 261251 4032 265624 4060
rect 261251 4029 261263 4032
rect 261205 4023 261263 4029
rect 265618 4020 265624 4032
rect 265676 4020 265682 4072
rect 265728 4032 268332 4060
rect 252557 3995 252615 4001
rect 252557 3961 252569 3995
rect 252603 3992 252615 3995
rect 254949 3995 255007 4001
rect 252603 3964 253934 3992
rect 252603 3961 252615 3964
rect 252557 3955 252615 3961
rect 250809 3927 250867 3933
rect 250809 3924 250821 3927
rect 242860 3896 250821 3924
rect 242860 3884 242866 3896
rect 250809 3893 250821 3896
rect 250855 3924 250867 3927
rect 251177 3927 251235 3933
rect 251177 3924 251189 3927
rect 250855 3896 251189 3924
rect 250855 3893 250867 3896
rect 250809 3887 250867 3893
rect 251177 3893 251189 3896
rect 251223 3924 251235 3927
rect 251545 3927 251603 3933
rect 251545 3924 251557 3927
rect 251223 3896 251557 3924
rect 251223 3893 251235 3896
rect 251177 3887 251235 3893
rect 251545 3893 251557 3896
rect 251591 3893 251603 3927
rect 253906 3924 253934 3964
rect 254949 3961 254961 3995
rect 254995 3992 255007 3995
rect 255317 3995 255375 4001
rect 255317 3992 255329 3995
rect 254995 3964 255329 3992
rect 254995 3961 255007 3964
rect 254949 3955 255007 3961
rect 255317 3961 255329 3964
rect 255363 3992 255375 3995
rect 256053 3995 256111 4001
rect 256053 3992 256065 3995
rect 255363 3964 256065 3992
rect 255363 3961 255375 3964
rect 255317 3955 255375 3961
rect 256053 3961 256065 3964
rect 256099 3961 256111 3995
rect 260098 3992 260104 4004
rect 256053 3955 256111 3961
rect 256160 3964 260104 3992
rect 256160 3924 256188 3964
rect 260098 3952 260104 3964
rect 260156 3952 260162 4004
rect 265728 4001 265756 4032
rect 260469 3995 260527 4001
rect 260469 3961 260481 3995
rect 260515 3992 260527 3995
rect 265713 3995 265771 4001
rect 260515 3964 265664 3992
rect 260515 3961 260527 3964
rect 260469 3955 260527 3961
rect 253906 3896 256188 3924
rect 257157 3927 257215 3933
rect 251545 3887 251603 3893
rect 257157 3893 257169 3927
rect 257203 3924 257215 3927
rect 258074 3924 258080 3936
rect 257203 3896 258080 3924
rect 257203 3893 257215 3896
rect 257157 3887 257215 3893
rect 258074 3884 258080 3896
rect 258132 3884 258138 3936
rect 258258 3884 258264 3936
rect 258316 3884 258322 3936
rect 258534 3884 258540 3936
rect 258592 3884 258598 3936
rect 259914 3884 259920 3936
rect 259972 3884 259978 3936
rect 264425 3927 264483 3933
rect 264425 3893 264437 3927
rect 264471 3924 264483 3927
rect 264790 3924 264796 3936
rect 264471 3896 264796 3924
rect 264471 3893 264483 3896
rect 264425 3887 264483 3893
rect 264790 3884 264796 3896
rect 264848 3884 264854 3936
rect 265636 3924 265664 3964
rect 265713 3961 265725 3995
rect 265759 3961 265771 3995
rect 265713 3955 265771 3961
rect 266280 3964 266952 3992
rect 266280 3924 266308 3964
rect 265636 3896 266308 3924
rect 266354 3884 266360 3936
rect 266412 3884 266418 3936
rect 266924 3924 266952 3964
rect 266998 3952 267004 4004
rect 267056 3952 267062 4004
rect 267829 3995 267887 4001
rect 267829 3961 267841 3995
rect 267875 3992 267887 3995
rect 267918 3992 267924 4004
rect 267875 3964 267924 3992
rect 267875 3961 267887 3964
rect 267829 3955 267887 3961
rect 267918 3952 267924 3964
rect 267976 3952 267982 4004
rect 268304 3992 268332 4032
rect 268378 4020 268384 4072
rect 268436 4020 268442 4072
rect 268838 4020 268844 4072
rect 268896 4020 268902 4072
rect 270788 3992 270816 4091
rect 270862 4088 270868 4140
rect 270920 4088 270926 4140
rect 268304 3964 270816 3992
rect 269022 3924 269028 3936
rect 266924 3896 269028 3924
rect 269022 3884 269028 3896
rect 269080 3884 269086 3936
rect 269390 3884 269396 3936
rect 269448 3924 269454 3936
rect 269485 3927 269543 3933
rect 269485 3924 269497 3927
rect 269448 3896 269497 3924
rect 269448 3884 269454 3896
rect 269485 3893 269497 3896
rect 269531 3893 269543 3927
rect 269485 3887 269543 3893
rect 270221 3927 270279 3933
rect 270221 3893 270233 3927
rect 270267 3924 270279 3927
rect 270494 3924 270500 3936
rect 270267 3896 270500 3924
rect 270267 3893 270279 3896
rect 270221 3887 270279 3893
rect 270494 3884 270500 3896
rect 270552 3884 270558 3936
rect 1104 3834 271492 3856
rect 1104 3782 34748 3834
rect 34800 3782 34812 3834
rect 34864 3782 34876 3834
rect 34928 3782 34940 3834
rect 34992 3782 35004 3834
rect 35056 3782 102345 3834
rect 102397 3782 102409 3834
rect 102461 3782 102473 3834
rect 102525 3782 102537 3834
rect 102589 3782 102601 3834
rect 102653 3782 169942 3834
rect 169994 3782 170006 3834
rect 170058 3782 170070 3834
rect 170122 3782 170134 3834
rect 170186 3782 170198 3834
rect 170250 3782 237539 3834
rect 237591 3782 237603 3834
rect 237655 3782 237667 3834
rect 237719 3782 237731 3834
rect 237783 3782 237795 3834
rect 237847 3782 271492 3834
rect 1104 3760 271492 3782
rect 3326 3680 3332 3732
rect 3384 3720 3390 3732
rect 36446 3720 36452 3732
rect 3384 3692 36452 3720
rect 3384 3680 3390 3692
rect 36446 3680 36452 3692
rect 36504 3680 36510 3732
rect 39942 3680 39948 3732
rect 40000 3720 40006 3732
rect 40000 3692 40816 3720
rect 40000 3680 40006 3692
rect 40788 3664 40816 3692
rect 66714 3680 66720 3732
rect 66772 3720 66778 3732
rect 67177 3723 67235 3729
rect 67177 3720 67189 3723
rect 66772 3692 67189 3720
rect 66772 3680 66778 3692
rect 67177 3689 67189 3692
rect 67223 3689 67235 3723
rect 67177 3683 67235 3689
rect 79226 3680 79232 3732
rect 79284 3720 79290 3732
rect 84010 3720 84016 3732
rect 79284 3692 84016 3720
rect 79284 3680 79290 3692
rect 84010 3680 84016 3692
rect 84068 3680 84074 3732
rect 87506 3680 87512 3732
rect 87564 3720 87570 3732
rect 88153 3723 88211 3729
rect 88153 3720 88165 3723
rect 87564 3692 88165 3720
rect 87564 3680 87570 3692
rect 88153 3689 88165 3692
rect 88199 3689 88211 3723
rect 98822 3720 98828 3732
rect 88153 3683 88211 3689
rect 96540 3692 98828 3720
rect 37737 3655 37795 3661
rect 37737 3621 37749 3655
rect 37783 3652 37795 3655
rect 40034 3652 40040 3664
rect 37783 3624 40040 3652
rect 37783 3621 37795 3624
rect 37737 3615 37795 3621
rect 40034 3612 40040 3624
rect 40092 3612 40098 3664
rect 40770 3612 40776 3664
rect 40828 3652 40834 3664
rect 42521 3655 42579 3661
rect 40828 3624 41092 3652
rect 40828 3612 40834 3624
rect 15102 3544 15108 3596
rect 15160 3584 15166 3596
rect 19334 3584 19340 3596
rect 15160 3556 19340 3584
rect 15160 3544 15166 3556
rect 19334 3544 19340 3556
rect 19392 3544 19398 3596
rect 24946 3544 24952 3596
rect 25004 3544 25010 3596
rect 25038 3476 25044 3528
rect 25096 3516 25102 3528
rect 25133 3519 25191 3525
rect 25133 3516 25145 3519
rect 25096 3488 25145 3516
rect 25096 3476 25102 3488
rect 25133 3485 25145 3488
rect 25179 3516 25191 3519
rect 25406 3516 25412 3528
rect 25179 3488 25412 3516
rect 25179 3485 25191 3488
rect 25133 3479 25191 3485
rect 25406 3476 25412 3488
rect 25464 3476 25470 3528
rect 25777 3519 25835 3525
rect 25777 3485 25789 3519
rect 25823 3516 25835 3519
rect 26234 3516 26240 3528
rect 25823 3488 26240 3516
rect 25823 3485 25835 3488
rect 25777 3479 25835 3485
rect 26234 3476 26240 3488
rect 26292 3476 26298 3528
rect 26510 3476 26516 3528
rect 26568 3476 26574 3528
rect 27249 3519 27307 3525
rect 27249 3485 27261 3519
rect 27295 3516 27307 3519
rect 27522 3516 27528 3528
rect 27295 3488 27528 3516
rect 27295 3485 27307 3488
rect 27249 3479 27307 3485
rect 27522 3476 27528 3488
rect 27580 3476 27586 3528
rect 36630 3476 36636 3528
rect 36688 3516 36694 3528
rect 36725 3519 36783 3525
rect 36725 3516 36737 3519
rect 36688 3488 36737 3516
rect 36688 3476 36694 3488
rect 36725 3485 36737 3488
rect 36771 3485 36783 3519
rect 36725 3479 36783 3485
rect 36817 3519 36875 3525
rect 36817 3485 36829 3519
rect 36863 3516 36875 3519
rect 37274 3516 37280 3528
rect 36863 3488 37280 3516
rect 36863 3485 36875 3488
rect 36817 3479 36875 3485
rect 37274 3476 37280 3488
rect 37332 3476 37338 3528
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 20714 3448 20720 3460
rect 11204 3420 20720 3448
rect 11204 3408 11210 3420
rect 20714 3408 20720 3420
rect 20772 3408 20778 3460
rect 22738 3408 22744 3460
rect 22796 3448 22802 3460
rect 27614 3448 27620 3460
rect 22796 3420 27620 3448
rect 22796 3408 22802 3420
rect 27614 3408 27620 3420
rect 27672 3408 27678 3460
rect 37185 3451 37243 3457
rect 37185 3448 37197 3451
rect 35912 3420 37197 3448
rect 35912 3392 35940 3420
rect 37185 3417 37197 3420
rect 37231 3417 37243 3451
rect 37476 3448 37504 3570
rect 37550 3544 37556 3596
rect 37608 3584 37614 3596
rect 37608 3556 41000 3584
rect 41064 3570 41092 3624
rect 42521 3621 42533 3655
rect 42567 3621 42579 3655
rect 42521 3615 42579 3621
rect 47949 3655 48007 3661
rect 47949 3621 47961 3655
rect 47995 3652 48007 3655
rect 47995 3624 51074 3652
rect 47995 3621 48007 3624
rect 47949 3615 48007 3621
rect 37608 3544 37614 3556
rect 40972 3516 41000 3556
rect 42536 3516 42564 3615
rect 48038 3584 48044 3596
rect 47702 3556 48044 3584
rect 48038 3544 48044 3556
rect 48096 3544 48102 3596
rect 40972 3488 42380 3516
rect 42536 3488 47900 3516
rect 38470 3448 38476 3460
rect 37476 3420 38476 3448
rect 37185 3411 37243 3417
rect 38470 3408 38476 3420
rect 38528 3408 38534 3460
rect 40221 3451 40279 3457
rect 40221 3417 40233 3451
rect 40267 3448 40279 3451
rect 40865 3451 40923 3457
rect 40865 3448 40877 3451
rect 40267 3420 40877 3448
rect 40267 3417 40279 3420
rect 40221 3411 40279 3417
rect 40865 3417 40877 3420
rect 40911 3448 40923 3451
rect 40954 3448 40960 3460
rect 40911 3420 40960 3448
rect 40911 3417 40923 3420
rect 40865 3411 40923 3417
rect 40954 3408 40960 3420
rect 41012 3408 41018 3460
rect 41064 3420 41414 3448
rect 23750 3340 23756 3392
rect 23808 3380 23814 3392
rect 25317 3383 25375 3389
rect 25317 3380 25329 3383
rect 23808 3352 25329 3380
rect 23808 3340 23814 3352
rect 25317 3349 25329 3352
rect 25363 3349 25375 3383
rect 25317 3343 25375 3349
rect 25958 3340 25964 3392
rect 26016 3340 26022 3392
rect 26694 3340 26700 3392
rect 26752 3340 26758 3392
rect 27430 3340 27436 3392
rect 27488 3340 27494 3392
rect 35894 3340 35900 3392
rect 35952 3340 35958 3392
rect 36078 3340 36084 3392
rect 36136 3380 36142 3392
rect 36449 3383 36507 3389
rect 36449 3380 36461 3383
rect 36136 3352 36461 3380
rect 36136 3340 36142 3352
rect 36449 3349 36461 3352
rect 36495 3349 36507 3383
rect 36449 3343 36507 3349
rect 37550 3340 37556 3392
rect 37608 3340 37614 3392
rect 38654 3340 38660 3392
rect 38712 3380 38718 3392
rect 40313 3383 40371 3389
rect 40313 3380 40325 3383
rect 38712 3352 40325 3380
rect 38712 3340 38718 3352
rect 40313 3349 40325 3352
rect 40359 3349 40371 3383
rect 40313 3343 40371 3349
rect 40402 3340 40408 3392
rect 40460 3380 40466 3392
rect 41064 3380 41092 3420
rect 40460 3352 41092 3380
rect 40460 3340 40466 3352
rect 41230 3340 41236 3392
rect 41288 3340 41294 3392
rect 41386 3380 41414 3420
rect 41506 3408 41512 3460
rect 41564 3408 41570 3460
rect 41598 3408 41604 3460
rect 41656 3408 41662 3460
rect 41966 3408 41972 3460
rect 42024 3408 42030 3460
rect 42352 3457 42380 3488
rect 42337 3451 42395 3457
rect 42337 3417 42349 3451
rect 42383 3417 42395 3451
rect 42337 3411 42395 3417
rect 46658 3408 46664 3460
rect 46716 3408 46722 3460
rect 46934 3408 46940 3460
rect 46992 3408 46998 3460
rect 47029 3451 47087 3457
rect 47029 3417 47041 3451
rect 47075 3448 47087 3451
rect 47210 3448 47216 3460
rect 47075 3420 47216 3448
rect 47075 3417 47087 3420
rect 47029 3411 47087 3417
rect 47210 3408 47216 3420
rect 47268 3408 47274 3460
rect 47394 3408 47400 3460
rect 47452 3408 47458 3460
rect 46109 3383 46167 3389
rect 46109 3380 46121 3383
rect 41386 3352 46121 3380
rect 46109 3349 46121 3352
rect 46155 3380 46167 3383
rect 47765 3383 47823 3389
rect 47765 3380 47777 3383
rect 46155 3352 47777 3380
rect 46155 3349 46167 3352
rect 46109 3343 46167 3349
rect 47765 3349 47777 3352
rect 47811 3349 47823 3383
rect 47872 3380 47900 3488
rect 51046 3448 51074 3624
rect 60734 3612 60740 3664
rect 60792 3652 60798 3664
rect 94222 3652 94228 3664
rect 60792 3624 94228 3652
rect 60792 3612 60798 3624
rect 94222 3612 94228 3624
rect 94280 3612 94286 3664
rect 77294 3584 77300 3596
rect 67100 3556 77300 3584
rect 51902 3476 51908 3528
rect 51960 3516 51966 3528
rect 66990 3516 66996 3528
rect 51960 3488 66996 3516
rect 51960 3476 51966 3488
rect 66990 3476 66996 3488
rect 67048 3476 67054 3528
rect 67100 3525 67128 3556
rect 77294 3544 77300 3556
rect 77352 3544 77358 3596
rect 82817 3587 82875 3593
rect 82817 3553 82829 3587
rect 82863 3584 82875 3587
rect 83185 3587 83243 3593
rect 83185 3584 83197 3587
rect 82863 3556 83197 3584
rect 82863 3553 82875 3556
rect 82817 3547 82875 3553
rect 83185 3553 83197 3556
rect 83231 3584 83243 3587
rect 94041 3587 94099 3593
rect 94041 3584 94053 3587
rect 83231 3556 85344 3584
rect 83231 3553 83243 3556
rect 83185 3547 83243 3553
rect 67085 3519 67143 3525
rect 67085 3485 67097 3519
rect 67131 3485 67143 3519
rect 67085 3479 67143 3485
rect 67174 3476 67180 3528
rect 67232 3516 67238 3528
rect 83461 3519 83519 3525
rect 83461 3516 83473 3519
rect 67232 3488 83473 3516
rect 67232 3476 67238 3488
rect 83461 3485 83473 3488
rect 83507 3485 83519 3519
rect 83461 3479 83519 3485
rect 79226 3448 79232 3460
rect 51046 3420 79232 3448
rect 79226 3408 79232 3420
rect 79284 3408 79290 3460
rect 79336 3420 83228 3448
rect 79336 3380 79364 3420
rect 47872 3352 79364 3380
rect 83200 3380 83228 3420
rect 83642 3408 83648 3460
rect 83700 3448 83706 3460
rect 84470 3448 84476 3460
rect 83700 3420 84476 3448
rect 83700 3408 83706 3420
rect 84470 3408 84476 3420
rect 84528 3448 84534 3460
rect 84930 3448 84936 3460
rect 84528 3420 84936 3448
rect 84528 3408 84534 3420
rect 84930 3408 84936 3420
rect 84988 3408 84994 3460
rect 85316 3457 85344 3556
rect 85500 3556 94053 3584
rect 85301 3451 85359 3457
rect 85301 3417 85313 3451
rect 85347 3448 85359 3451
rect 85390 3448 85396 3460
rect 85347 3420 85396 3448
rect 85347 3417 85359 3420
rect 85301 3411 85359 3417
rect 85390 3408 85396 3420
rect 85448 3408 85454 3460
rect 85500 3380 85528 3556
rect 94041 3553 94053 3556
rect 94087 3553 94099 3587
rect 94041 3547 94099 3553
rect 87969 3519 88027 3525
rect 87969 3485 87981 3519
rect 88015 3516 88027 3519
rect 88242 3516 88248 3528
rect 88015 3488 88248 3516
rect 88015 3485 88027 3488
rect 87969 3479 88027 3485
rect 88242 3476 88248 3488
rect 88300 3476 88306 3528
rect 91741 3519 91799 3525
rect 91741 3516 91753 3519
rect 88352 3488 91753 3516
rect 83200 3352 85528 3380
rect 47765 3343 47823 3349
rect 85666 3340 85672 3392
rect 85724 3340 85730 3392
rect 86034 3340 86040 3392
rect 86092 3380 86098 3392
rect 88352 3380 88380 3488
rect 91741 3485 91753 3488
rect 91787 3485 91799 3519
rect 91741 3479 91799 3485
rect 95878 3476 95884 3528
rect 95936 3476 95942 3528
rect 91646 3408 91652 3460
rect 91704 3448 91710 3460
rect 91922 3448 91928 3460
rect 91704 3420 91928 3448
rect 91704 3408 91710 3420
rect 91922 3408 91928 3420
rect 91980 3408 91986 3460
rect 93581 3451 93639 3457
rect 93581 3417 93593 3451
rect 93627 3417 93639 3451
rect 93581 3411 93639 3417
rect 94225 3451 94283 3457
rect 94225 3417 94237 3451
rect 94271 3448 94283 3451
rect 95050 3448 95056 3460
rect 94271 3420 95056 3448
rect 94271 3417 94283 3420
rect 94225 3411 94283 3417
rect 86092 3352 88380 3380
rect 89073 3383 89131 3389
rect 86092 3340 86098 3352
rect 89073 3349 89085 3383
rect 89119 3380 89131 3383
rect 89806 3380 89812 3392
rect 89119 3352 89812 3380
rect 89119 3349 89131 3352
rect 89073 3343 89131 3349
rect 89806 3340 89812 3352
rect 89864 3340 89870 3392
rect 93596 3380 93624 3411
rect 95050 3408 95056 3420
rect 95108 3408 95114 3460
rect 96540 3380 96568 3692
rect 98822 3680 98828 3692
rect 98880 3680 98886 3732
rect 98914 3680 98920 3732
rect 98972 3720 98978 3732
rect 104253 3723 104311 3729
rect 104253 3720 104265 3723
rect 98972 3692 104265 3720
rect 98972 3680 98978 3692
rect 104253 3689 104265 3692
rect 104299 3689 104311 3723
rect 104253 3683 104311 3689
rect 98638 3612 98644 3664
rect 98696 3652 98702 3664
rect 99098 3652 99104 3664
rect 98696 3624 99104 3652
rect 98696 3612 98702 3624
rect 99098 3612 99104 3624
rect 99156 3612 99162 3664
rect 99466 3612 99472 3664
rect 99524 3652 99530 3664
rect 104158 3652 104164 3664
rect 99524 3624 104164 3652
rect 99524 3612 99530 3624
rect 104158 3612 104164 3624
rect 104216 3612 104222 3664
rect 104268 3652 104296 3683
rect 104526 3680 104532 3732
rect 104584 3720 104590 3732
rect 104584 3692 112944 3720
rect 104584 3680 104590 3692
rect 104268 3624 105400 3652
rect 96614 3544 96620 3596
rect 96672 3544 96678 3596
rect 97258 3544 97264 3596
rect 97316 3544 97322 3596
rect 97534 3544 97540 3596
rect 97592 3544 97598 3596
rect 97675 3587 97733 3593
rect 97675 3553 97687 3587
rect 97721 3584 97733 3587
rect 100570 3584 100576 3596
rect 97721 3556 100576 3584
rect 97721 3553 97733 3556
rect 97675 3547 97733 3553
rect 100570 3544 100576 3556
rect 100628 3544 100634 3596
rect 101306 3544 101312 3596
rect 101364 3544 101370 3596
rect 101398 3544 101404 3596
rect 101456 3584 101462 3596
rect 102870 3584 102876 3596
rect 101456 3556 102876 3584
rect 101456 3544 101462 3556
rect 102870 3544 102876 3556
rect 102928 3544 102934 3596
rect 103790 3544 103796 3596
rect 103848 3584 103854 3596
rect 104526 3584 104532 3596
rect 103848 3556 104532 3584
rect 103848 3544 103854 3556
rect 104526 3544 104532 3556
rect 104584 3544 104590 3596
rect 104621 3587 104679 3593
rect 104621 3553 104633 3587
rect 104667 3584 104679 3587
rect 105262 3584 105268 3596
rect 104667 3556 105268 3584
rect 104667 3553 104679 3556
rect 104621 3547 104679 3553
rect 105262 3544 105268 3556
rect 105320 3544 105326 3596
rect 105372 3593 105400 3624
rect 105446 3612 105452 3664
rect 105504 3652 105510 3664
rect 112714 3652 112720 3664
rect 105504 3624 112720 3652
rect 105504 3612 105510 3624
rect 112714 3612 112720 3624
rect 112772 3612 112778 3664
rect 105357 3587 105415 3593
rect 105357 3553 105369 3587
rect 105403 3584 105415 3587
rect 107013 3587 107071 3593
rect 107013 3584 107025 3587
rect 105403 3556 107025 3584
rect 105403 3553 105415 3556
rect 105357 3547 105415 3553
rect 107013 3553 107025 3556
rect 107059 3553 107071 3587
rect 107013 3547 107071 3553
rect 96706 3476 96712 3528
rect 96764 3516 96770 3528
rect 96801 3519 96859 3525
rect 96801 3516 96813 3519
rect 96764 3488 96813 3516
rect 96764 3476 96770 3488
rect 96801 3485 96813 3488
rect 96847 3485 96859 3519
rect 96801 3479 96859 3485
rect 97810 3476 97816 3528
rect 97868 3476 97874 3528
rect 98730 3476 98736 3528
rect 98788 3516 98794 3528
rect 99469 3519 99527 3525
rect 99469 3516 99481 3519
rect 98788 3488 99481 3516
rect 98788 3476 98794 3488
rect 99469 3485 99481 3488
rect 99515 3485 99527 3519
rect 99469 3479 99527 3485
rect 101490 3476 101496 3528
rect 101548 3516 101554 3528
rect 101953 3519 102011 3525
rect 101953 3516 101965 3519
rect 101548 3488 101965 3516
rect 101548 3476 101554 3488
rect 101953 3485 101965 3488
rect 101999 3485 102011 3519
rect 101953 3479 102011 3485
rect 104158 3476 104164 3528
rect 104216 3516 104222 3528
rect 104216 3488 104664 3516
rect 104216 3476 104222 3488
rect 98380 3420 99052 3448
rect 93596 3352 96568 3380
rect 97258 3340 97264 3392
rect 97316 3380 97322 3392
rect 98380 3380 98408 3420
rect 97316 3352 98408 3380
rect 97316 3340 97322 3352
rect 98454 3340 98460 3392
rect 98512 3340 98518 3392
rect 98638 3340 98644 3392
rect 98696 3380 98702 3392
rect 98733 3383 98791 3389
rect 98733 3380 98745 3383
rect 98696 3352 98745 3380
rect 98696 3340 98702 3352
rect 98733 3349 98745 3352
rect 98779 3349 98791 3383
rect 99024 3380 99052 3420
rect 99098 3408 99104 3460
rect 99156 3448 99162 3460
rect 99653 3451 99711 3457
rect 99156 3420 99604 3448
rect 99156 3408 99162 3420
rect 99466 3380 99472 3392
rect 99024 3352 99472 3380
rect 98733 3343 98791 3349
rect 99466 3340 99472 3352
rect 99524 3340 99530 3392
rect 99576 3380 99604 3420
rect 99653 3417 99665 3451
rect 99699 3448 99711 3451
rect 99742 3448 99748 3460
rect 99699 3420 99748 3448
rect 99699 3417 99711 3420
rect 99653 3411 99711 3417
rect 99742 3408 99748 3420
rect 99800 3448 99806 3460
rect 102137 3451 102195 3457
rect 102137 3448 102149 3451
rect 99800 3420 102149 3448
rect 99800 3408 99806 3420
rect 102137 3417 102149 3420
rect 102183 3417 102195 3451
rect 104636 3448 104664 3488
rect 104805 3451 104863 3457
rect 104636 3420 104756 3448
rect 102137 3411 102195 3417
rect 101306 3380 101312 3392
rect 99576 3352 101312 3380
rect 101306 3340 101312 3352
rect 101364 3340 101370 3392
rect 102152 3380 102180 3411
rect 103146 3380 103152 3392
rect 102152 3352 103152 3380
rect 103146 3340 103152 3352
rect 103204 3380 103210 3392
rect 104618 3380 104624 3392
rect 103204 3352 104624 3380
rect 103204 3340 103210 3352
rect 104618 3340 104624 3352
rect 104676 3340 104682 3392
rect 104728 3380 104756 3420
rect 104805 3417 104817 3451
rect 104851 3448 104863 3451
rect 104894 3448 104900 3460
rect 104851 3420 104900 3448
rect 104851 3417 104863 3420
rect 104805 3411 104863 3417
rect 104894 3408 104900 3420
rect 104952 3408 104958 3460
rect 106918 3380 106924 3392
rect 104728 3352 106924 3380
rect 106918 3340 106924 3352
rect 106976 3340 106982 3392
rect 107028 3380 107056 3547
rect 108850 3544 108856 3596
rect 108908 3584 108914 3596
rect 109129 3587 109187 3593
rect 109129 3584 109141 3587
rect 108908 3556 109141 3584
rect 108908 3544 108914 3556
rect 109129 3553 109141 3556
rect 109175 3553 109187 3587
rect 109129 3547 109187 3553
rect 110506 3544 110512 3596
rect 110564 3584 110570 3596
rect 110966 3584 110972 3596
rect 110564 3556 110972 3584
rect 110564 3544 110570 3556
rect 110966 3544 110972 3556
rect 111024 3544 111030 3596
rect 112916 3516 112944 3692
rect 113450 3680 113456 3732
rect 113508 3720 113514 3732
rect 115842 3720 115848 3732
rect 113508 3692 115848 3720
rect 113508 3680 113514 3692
rect 115842 3680 115848 3692
rect 115900 3680 115906 3732
rect 115934 3680 115940 3732
rect 115992 3720 115998 3732
rect 115992 3692 116532 3720
rect 115992 3680 115998 3692
rect 116504 3652 116532 3692
rect 116762 3680 116768 3732
rect 116820 3680 116826 3732
rect 152366 3720 152372 3732
rect 118666 3692 152372 3720
rect 118666 3652 118694 3692
rect 152366 3680 152372 3692
rect 152424 3680 152430 3732
rect 152826 3680 152832 3732
rect 152884 3720 152890 3732
rect 155678 3720 155684 3732
rect 152884 3692 155684 3720
rect 152884 3680 152890 3692
rect 155678 3680 155684 3692
rect 155736 3680 155742 3732
rect 157521 3723 157579 3729
rect 157521 3689 157533 3723
rect 157567 3720 157579 3723
rect 158254 3720 158260 3732
rect 157567 3692 158260 3720
rect 157567 3689 157579 3692
rect 157521 3683 157579 3689
rect 158254 3680 158260 3692
rect 158312 3680 158318 3732
rect 158622 3680 158628 3732
rect 158680 3720 158686 3732
rect 160189 3723 160247 3729
rect 158680 3692 160140 3720
rect 158680 3680 158686 3692
rect 116504 3624 118694 3652
rect 119798 3612 119804 3664
rect 119856 3612 119862 3664
rect 120994 3612 121000 3664
rect 121052 3612 121058 3664
rect 143442 3612 143448 3664
rect 143500 3652 143506 3664
rect 143721 3655 143779 3661
rect 143721 3652 143733 3655
rect 143500 3624 143733 3652
rect 143500 3612 143506 3624
rect 143721 3621 143733 3624
rect 143767 3621 143779 3655
rect 143721 3615 143779 3621
rect 144730 3612 144736 3664
rect 144788 3612 144794 3664
rect 144822 3612 144828 3664
rect 144880 3652 144886 3664
rect 144917 3655 144975 3661
rect 144917 3652 144929 3655
rect 144880 3624 144929 3652
rect 144880 3612 144886 3624
rect 144917 3621 144929 3624
rect 144963 3621 144975 3655
rect 147217 3655 147275 3661
rect 144917 3615 144975 3621
rect 145300 3624 146156 3652
rect 112990 3544 112996 3596
rect 113048 3584 113054 3596
rect 115290 3584 115296 3596
rect 113048 3556 115296 3584
rect 113048 3544 113054 3556
rect 115290 3544 115296 3556
rect 115348 3584 115354 3596
rect 115569 3587 115627 3593
rect 115569 3584 115581 3587
rect 115348 3556 115581 3584
rect 115348 3544 115354 3556
rect 115569 3553 115581 3556
rect 115615 3553 115627 3587
rect 115569 3547 115627 3553
rect 115658 3544 115664 3596
rect 115716 3584 115722 3596
rect 115845 3587 115903 3593
rect 115845 3584 115857 3587
rect 115716 3556 115857 3584
rect 115716 3544 115722 3556
rect 115845 3553 115857 3556
rect 115891 3553 115903 3587
rect 115845 3547 115903 3553
rect 115983 3587 116041 3593
rect 115983 3553 115995 3587
rect 116029 3584 116041 3587
rect 117222 3584 117228 3596
rect 116029 3556 117228 3584
rect 116029 3553 116041 3556
rect 115983 3547 116041 3553
rect 117222 3544 117228 3556
rect 117280 3544 117286 3596
rect 118970 3544 118976 3596
rect 119028 3584 119034 3596
rect 119157 3587 119215 3593
rect 119157 3584 119169 3587
rect 119028 3556 119169 3584
rect 119028 3544 119034 3556
rect 119157 3553 119169 3556
rect 119203 3553 119215 3587
rect 119157 3547 119215 3553
rect 120074 3544 120080 3596
rect 120132 3544 120138 3596
rect 120350 3544 120356 3596
rect 120408 3544 120414 3596
rect 141418 3584 141424 3596
rect 120920 3556 141424 3584
rect 112916 3488 113404 3516
rect 109310 3408 109316 3460
rect 109368 3408 109374 3460
rect 113174 3380 113180 3392
rect 107028 3352 113180 3380
rect 113174 3340 113180 3352
rect 113232 3340 113238 3392
rect 113376 3380 113404 3488
rect 114922 3476 114928 3528
rect 114980 3476 114986 3528
rect 115106 3476 115112 3528
rect 115164 3476 115170 3528
rect 116118 3476 116124 3528
rect 116176 3476 116182 3528
rect 119338 3476 119344 3528
rect 119396 3476 119402 3528
rect 120166 3476 120172 3528
rect 120224 3525 120230 3528
rect 120224 3519 120252 3525
rect 120240 3485 120252 3519
rect 120224 3479 120252 3485
rect 120224 3476 120230 3479
rect 120920 3380 120948 3556
rect 141418 3544 141424 3556
rect 141476 3544 141482 3596
rect 142982 3544 142988 3596
rect 143040 3584 143046 3596
rect 143077 3587 143135 3593
rect 143077 3584 143089 3587
rect 143040 3556 143089 3584
rect 143040 3544 143046 3556
rect 143077 3553 143089 3556
rect 143123 3553 143135 3587
rect 143077 3547 143135 3553
rect 143994 3544 144000 3596
rect 144052 3544 144058 3596
rect 144135 3587 144193 3593
rect 144135 3553 144147 3587
rect 144181 3584 144193 3587
rect 144638 3584 144644 3596
rect 144181 3556 144644 3584
rect 144181 3553 144193 3556
rect 144135 3547 144193 3553
rect 144638 3544 144644 3556
rect 144696 3544 144702 3596
rect 144748 3584 144776 3612
rect 145300 3584 145328 3624
rect 144748 3556 145328 3584
rect 145374 3544 145380 3596
rect 145432 3544 145438 3596
rect 146021 3587 146079 3593
rect 146021 3584 146033 3587
rect 145484 3556 146033 3584
rect 122558 3476 122564 3528
rect 122616 3476 122622 3528
rect 138934 3476 138940 3528
rect 138992 3476 138998 3528
rect 143166 3476 143172 3528
rect 143224 3516 143230 3528
rect 143261 3519 143319 3525
rect 143261 3516 143273 3519
rect 143224 3488 143273 3516
rect 143224 3476 143230 3488
rect 143261 3485 143273 3488
rect 143307 3485 143319 3519
rect 143261 3479 143319 3485
rect 144270 3476 144276 3528
rect 144328 3476 144334 3528
rect 139118 3408 139124 3460
rect 139176 3408 139182 3460
rect 140682 3408 140688 3460
rect 140740 3448 140746 3460
rect 140777 3451 140835 3457
rect 140777 3448 140789 3451
rect 140740 3420 140789 3448
rect 140740 3408 140746 3420
rect 140777 3417 140789 3420
rect 140823 3417 140835 3451
rect 140777 3411 140835 3417
rect 144822 3408 144828 3460
rect 144880 3448 144886 3460
rect 145484 3448 145512 3556
rect 146021 3553 146033 3556
rect 146067 3553 146079 3587
rect 146128 3584 146156 3624
rect 147217 3621 147229 3655
rect 147263 3652 147275 3655
rect 147950 3652 147956 3664
rect 147263 3624 147956 3652
rect 147263 3621 147275 3624
rect 147217 3615 147275 3621
rect 147950 3612 147956 3624
rect 148008 3612 148014 3664
rect 148042 3612 148048 3664
rect 148100 3652 148106 3664
rect 154482 3652 154488 3664
rect 148100 3624 154488 3652
rect 148100 3612 148106 3624
rect 154482 3612 154488 3624
rect 154540 3652 154546 3664
rect 156046 3652 156052 3664
rect 154540 3624 156052 3652
rect 154540 3612 154546 3624
rect 156046 3612 156052 3624
rect 156104 3612 156110 3664
rect 159008 3661 159036 3692
rect 158993 3655 159051 3661
rect 158993 3621 159005 3655
rect 159039 3621 159051 3655
rect 160112 3652 160140 3692
rect 160189 3689 160201 3723
rect 160235 3720 160247 3723
rect 161014 3720 161020 3732
rect 160235 3692 161020 3720
rect 160235 3689 160247 3692
rect 160189 3683 160247 3689
rect 161014 3680 161020 3692
rect 161072 3680 161078 3732
rect 161934 3680 161940 3732
rect 161992 3720 161998 3732
rect 173158 3720 173164 3732
rect 161992 3692 173164 3720
rect 161992 3680 161998 3692
rect 173158 3680 173164 3692
rect 173216 3680 173222 3732
rect 207474 3680 207480 3732
rect 207532 3720 207538 3732
rect 217045 3723 217103 3729
rect 217045 3720 217057 3723
rect 207532 3692 210464 3720
rect 207532 3680 207538 3692
rect 162670 3652 162676 3664
rect 160112 3624 162676 3652
rect 158993 3615 159051 3621
rect 162670 3612 162676 3624
rect 162728 3612 162734 3664
rect 210050 3652 210056 3664
rect 209332 3624 210056 3652
rect 146573 3587 146631 3593
rect 146573 3584 146585 3587
rect 146128 3556 146585 3584
rect 146021 3547 146079 3553
rect 146573 3553 146585 3556
rect 146619 3584 146631 3587
rect 148962 3584 148968 3596
rect 146619 3556 148968 3584
rect 146619 3553 146631 3556
rect 146573 3547 146631 3553
rect 148962 3544 148968 3556
rect 149020 3544 149026 3596
rect 154574 3544 154580 3596
rect 154632 3584 154638 3596
rect 155681 3587 155739 3593
rect 155681 3584 155693 3587
rect 154632 3556 155693 3584
rect 154632 3544 154638 3556
rect 155681 3553 155693 3556
rect 155727 3553 155739 3587
rect 155681 3547 155739 3553
rect 156322 3544 156328 3596
rect 156380 3544 156386 3596
rect 156598 3544 156604 3596
rect 156656 3544 156662 3596
rect 156690 3544 156696 3596
rect 156748 3593 156754 3596
rect 156748 3587 156776 3593
rect 156764 3553 156776 3587
rect 156748 3547 156776 3553
rect 156748 3544 156754 3547
rect 156874 3544 156880 3596
rect 156932 3544 156938 3596
rect 158346 3544 158352 3596
rect 158404 3544 158410 3596
rect 159266 3544 159272 3596
rect 159324 3544 159330 3596
rect 159542 3544 159548 3596
rect 159600 3544 159606 3596
rect 176654 3584 176660 3596
rect 160112 3556 176660 3584
rect 145561 3519 145619 3525
rect 145561 3485 145573 3519
rect 145607 3485 145619 3519
rect 145561 3479 145619 3485
rect 144880 3420 145512 3448
rect 144880 3408 144886 3420
rect 113376 3352 120948 3380
rect 122834 3340 122840 3392
rect 122892 3340 122898 3392
rect 138566 3340 138572 3392
rect 138624 3380 138630 3392
rect 138661 3383 138719 3389
rect 138661 3380 138673 3383
rect 138624 3352 138673 3380
rect 138624 3340 138630 3352
rect 138661 3349 138673 3352
rect 138707 3380 138719 3383
rect 140700 3380 140728 3408
rect 138707 3352 140728 3380
rect 138707 3349 138719 3352
rect 138661 3343 138719 3349
rect 143810 3340 143816 3392
rect 143868 3380 143874 3392
rect 145576 3380 145604 3479
rect 146294 3476 146300 3528
rect 146352 3476 146358 3528
rect 146478 3525 146484 3528
rect 146435 3519 146484 3525
rect 146435 3485 146447 3519
rect 146481 3485 146484 3519
rect 146435 3479 146484 3485
rect 146478 3476 146484 3479
rect 146536 3476 146542 3528
rect 147490 3476 147496 3528
rect 147548 3516 147554 3528
rect 148229 3519 148287 3525
rect 148229 3516 148241 3519
rect 147548 3488 148241 3516
rect 147548 3476 147554 3488
rect 148229 3485 148241 3488
rect 148275 3485 148287 3519
rect 148229 3479 148287 3485
rect 152366 3476 152372 3528
rect 152424 3516 152430 3528
rect 154666 3516 154672 3528
rect 152424 3488 154672 3516
rect 152424 3476 152430 3488
rect 154666 3476 154672 3488
rect 154724 3476 154730 3528
rect 155218 3476 155224 3528
rect 155276 3476 155282 3528
rect 155862 3476 155868 3528
rect 155920 3476 155926 3528
rect 158530 3476 158536 3528
rect 158588 3476 158594 3528
rect 159450 3525 159456 3528
rect 159407 3519 159456 3525
rect 159407 3485 159419 3519
rect 159453 3485 159456 3519
rect 159407 3479 159456 3485
rect 159450 3476 159456 3479
rect 159508 3476 159514 3528
rect 148410 3408 148416 3460
rect 148468 3408 148474 3460
rect 148686 3408 148692 3460
rect 148744 3448 148750 3460
rect 148870 3448 148876 3460
rect 148744 3420 148876 3448
rect 148744 3408 148750 3420
rect 148870 3408 148876 3420
rect 148928 3408 148934 3460
rect 150066 3408 150072 3460
rect 150124 3408 150130 3460
rect 151170 3408 151176 3460
rect 151228 3448 151234 3460
rect 154850 3448 154856 3460
rect 151228 3420 154856 3448
rect 151228 3408 151234 3420
rect 154850 3408 154856 3420
rect 154908 3408 154914 3460
rect 143868 3352 145604 3380
rect 143868 3340 143874 3352
rect 146846 3340 146852 3392
rect 146904 3380 146910 3392
rect 149146 3380 149152 3392
rect 146904 3352 149152 3380
rect 146904 3340 146910 3352
rect 149146 3340 149152 3352
rect 149204 3340 149210 3392
rect 154390 3340 154396 3392
rect 154448 3380 154454 3392
rect 155405 3383 155463 3389
rect 155405 3380 155417 3383
rect 154448 3352 155417 3380
rect 154448 3340 154454 3352
rect 155405 3349 155417 3352
rect 155451 3380 155463 3383
rect 156874 3380 156880 3392
rect 155451 3352 156880 3380
rect 155451 3349 155463 3352
rect 155405 3343 155463 3349
rect 156874 3340 156880 3352
rect 156932 3340 156938 3392
rect 156966 3340 156972 3392
rect 157024 3380 157030 3392
rect 160112 3380 160140 3556
rect 176654 3544 176660 3556
rect 176712 3544 176718 3596
rect 205082 3544 205088 3596
rect 205140 3584 205146 3596
rect 205140 3556 206508 3584
rect 205140 3544 205146 3556
rect 160830 3476 160836 3528
rect 160888 3476 160894 3528
rect 162486 3476 162492 3528
rect 162544 3516 162550 3528
rect 204254 3516 204260 3528
rect 162544 3488 204260 3516
rect 162544 3476 162550 3488
rect 204254 3476 204260 3488
rect 204312 3476 204318 3528
rect 204898 3476 204904 3528
rect 204956 3476 204962 3528
rect 206480 3516 206508 3556
rect 207198 3544 207204 3596
rect 207256 3544 207262 3596
rect 207658 3544 207664 3596
rect 207716 3584 207722 3596
rect 209332 3593 209360 3624
rect 210050 3612 210056 3624
rect 210108 3612 210114 3664
rect 209317 3587 209375 3593
rect 209317 3584 209329 3587
rect 207716 3556 209329 3584
rect 207716 3544 207722 3556
rect 209317 3553 209329 3556
rect 209363 3553 209375 3587
rect 209317 3547 209375 3553
rect 206480 3488 207244 3516
rect 161017 3451 161075 3457
rect 161017 3417 161029 3451
rect 161063 3448 161075 3451
rect 161290 3448 161296 3460
rect 161063 3420 161296 3448
rect 161063 3417 161075 3420
rect 161017 3411 161075 3417
rect 161290 3408 161296 3420
rect 161348 3408 161354 3460
rect 162670 3408 162676 3460
rect 162728 3408 162734 3460
rect 163406 3408 163412 3460
rect 163464 3448 163470 3460
rect 180886 3448 180892 3460
rect 163464 3420 180892 3448
rect 163464 3408 163470 3420
rect 180886 3408 180892 3420
rect 180944 3408 180950 3460
rect 205082 3408 205088 3460
rect 205140 3408 205146 3460
rect 206741 3451 206799 3457
rect 206741 3417 206753 3451
rect 206787 3448 206799 3451
rect 207106 3448 207112 3460
rect 206787 3420 207112 3448
rect 206787 3417 206799 3420
rect 206741 3411 206799 3417
rect 157024 3352 160140 3380
rect 157024 3340 157030 3352
rect 160554 3340 160560 3392
rect 160612 3340 160618 3392
rect 160646 3340 160652 3392
rect 160704 3380 160710 3392
rect 203889 3383 203947 3389
rect 203889 3380 203901 3383
rect 160704 3352 203901 3380
rect 160704 3340 160710 3352
rect 203889 3349 203901 3352
rect 203935 3380 203947 3383
rect 204257 3383 204315 3389
rect 204257 3380 204269 3383
rect 203935 3352 204269 3380
rect 203935 3349 203947 3352
rect 203889 3343 203947 3349
rect 204257 3349 204269 3352
rect 204303 3380 204315 3383
rect 206756 3380 206784 3411
rect 207106 3408 207112 3420
rect 207164 3408 207170 3460
rect 207216 3448 207244 3488
rect 207385 3451 207443 3457
rect 207385 3448 207397 3451
rect 207216 3420 207397 3448
rect 207385 3417 207397 3420
rect 207431 3448 207443 3451
rect 207750 3448 207756 3460
rect 207431 3420 207756 3448
rect 207431 3417 207443 3420
rect 207385 3411 207443 3417
rect 207750 3408 207756 3420
rect 207808 3408 207814 3460
rect 209240 3420 209452 3448
rect 204303 3352 206784 3380
rect 204303 3349 204315 3352
rect 204257 3343 204315 3349
rect 208394 3340 208400 3392
rect 208452 3380 208458 3392
rect 209240 3380 209268 3420
rect 208452 3352 209268 3380
rect 209424 3380 209452 3420
rect 209682 3408 209688 3460
rect 209740 3448 209746 3460
rect 210326 3448 210332 3460
rect 209740 3420 210332 3448
rect 209740 3408 209746 3420
rect 210326 3408 210332 3420
rect 210384 3408 210390 3460
rect 210142 3380 210148 3392
rect 209424 3352 210148 3380
rect 208452 3340 208458 3352
rect 210142 3340 210148 3352
rect 210200 3340 210206 3392
rect 210436 3380 210464 3692
rect 210528 3692 217057 3720
rect 210528 3593 210556 3692
rect 217045 3689 217057 3692
rect 217091 3689 217103 3723
rect 217045 3683 217103 3689
rect 222565 3723 222623 3729
rect 222565 3689 222577 3723
rect 222611 3720 222623 3723
rect 224494 3720 224500 3732
rect 222611 3692 224500 3720
rect 222611 3689 222623 3692
rect 222565 3683 222623 3689
rect 224494 3680 224500 3692
rect 224552 3680 224558 3732
rect 225230 3680 225236 3732
rect 225288 3720 225294 3732
rect 225288 3692 227116 3720
rect 225288 3680 225294 3692
rect 210602 3612 210608 3664
rect 210660 3652 210666 3664
rect 214650 3652 214656 3664
rect 210660 3624 213224 3652
rect 210660 3612 210666 3624
rect 210513 3587 210571 3593
rect 210513 3553 210525 3587
rect 210559 3553 210571 3587
rect 210513 3547 210571 3553
rect 210694 3544 210700 3596
rect 210752 3544 210758 3596
rect 211246 3544 211252 3596
rect 211304 3584 211310 3596
rect 212445 3587 212503 3593
rect 212445 3584 212457 3587
rect 211304 3556 212457 3584
rect 211304 3544 211310 3556
rect 212445 3553 212457 3556
rect 212491 3553 212503 3587
rect 212445 3547 212503 3553
rect 213086 3544 213092 3596
rect 213144 3544 213150 3596
rect 213196 3584 213224 3624
rect 214024 3624 214656 3652
rect 214024 3584 214052 3624
rect 214650 3612 214656 3624
rect 214708 3612 214714 3664
rect 215754 3612 215760 3664
rect 215812 3652 215818 3664
rect 215849 3655 215907 3661
rect 215849 3652 215861 3655
rect 215812 3624 215861 3652
rect 215812 3612 215818 3624
rect 215849 3621 215861 3624
rect 215895 3621 215907 3655
rect 217410 3652 217416 3664
rect 215849 3615 215907 3621
rect 216968 3624 217416 3652
rect 213196 3556 214052 3584
rect 214374 3544 214380 3596
rect 214432 3584 214438 3596
rect 215205 3587 215263 3593
rect 215205 3584 215217 3587
rect 214432 3556 215217 3584
rect 214432 3544 214438 3556
rect 215205 3553 215217 3556
rect 215251 3553 215263 3587
rect 215205 3547 215263 3553
rect 216122 3544 216128 3596
rect 216180 3544 216186 3596
rect 216242 3587 216300 3593
rect 216242 3553 216254 3587
rect 216288 3584 216300 3587
rect 216968 3584 216996 3624
rect 217410 3612 217416 3624
rect 217468 3612 217474 3664
rect 217502 3612 217508 3664
rect 217560 3652 217566 3664
rect 226242 3652 226248 3664
rect 217560 3624 226248 3652
rect 217560 3612 217566 3624
rect 226242 3612 226248 3624
rect 226300 3612 226306 3664
rect 227088 3652 227116 3692
rect 227346 3680 227352 3732
rect 227404 3680 227410 3732
rect 251450 3680 251456 3732
rect 251508 3720 251514 3732
rect 256510 3720 256516 3732
rect 251508 3692 256516 3720
rect 251508 3680 251514 3692
rect 256510 3680 256516 3692
rect 256568 3720 256574 3732
rect 258534 3720 258540 3732
rect 256568 3692 258540 3720
rect 256568 3680 256574 3692
rect 258534 3680 258540 3692
rect 258592 3720 258598 3732
rect 260561 3723 260619 3729
rect 260561 3720 260573 3723
rect 258592 3692 260573 3720
rect 258592 3680 258598 3692
rect 260561 3689 260573 3692
rect 260607 3689 260619 3723
rect 260561 3683 260619 3689
rect 265342 3680 265348 3732
rect 265400 3680 265406 3732
rect 265986 3680 265992 3732
rect 266044 3680 266050 3732
rect 267185 3723 267243 3729
rect 267185 3689 267197 3723
rect 267231 3720 267243 3723
rect 268473 3723 268531 3729
rect 267231 3692 268424 3720
rect 267231 3689 267243 3692
rect 267185 3683 267243 3689
rect 238570 3652 238576 3664
rect 227088 3624 238576 3652
rect 238570 3612 238576 3624
rect 238628 3612 238634 3664
rect 259914 3612 259920 3664
rect 259972 3652 259978 3664
rect 268010 3652 268016 3664
rect 259972 3624 268016 3652
rect 259972 3612 259978 3624
rect 268010 3612 268016 3624
rect 268068 3612 268074 3664
rect 268396 3652 268424 3692
rect 268473 3689 268485 3723
rect 268519 3720 268531 3723
rect 269482 3720 269488 3732
rect 268519 3692 269488 3720
rect 268519 3689 268531 3692
rect 268473 3683 268531 3689
rect 269482 3680 269488 3692
rect 269540 3680 269546 3732
rect 270037 3723 270095 3729
rect 270037 3689 270049 3723
rect 270083 3720 270095 3723
rect 270586 3720 270592 3732
rect 270083 3692 270592 3720
rect 270083 3689 270095 3692
rect 270037 3683 270095 3689
rect 270586 3680 270592 3692
rect 270644 3680 270650 3732
rect 270681 3723 270739 3729
rect 270681 3689 270693 3723
rect 270727 3720 270739 3723
rect 270770 3720 270776 3732
rect 270727 3692 270776 3720
rect 270727 3689 270739 3692
rect 270681 3683 270739 3689
rect 270770 3680 270776 3692
rect 270828 3680 270834 3732
rect 269206 3652 269212 3664
rect 268396 3624 269212 3652
rect 269206 3612 269212 3624
rect 269264 3612 269270 3664
rect 269301 3655 269359 3661
rect 269301 3621 269313 3655
rect 269347 3652 269359 3655
rect 269574 3652 269580 3664
rect 269347 3624 269580 3652
rect 269347 3621 269359 3624
rect 269301 3615 269359 3621
rect 269574 3612 269580 3624
rect 269632 3612 269638 3664
rect 269850 3612 269856 3664
rect 269908 3612 269914 3664
rect 216288 3556 216996 3584
rect 216288 3553 216300 3556
rect 216242 3547 216300 3553
rect 218882 3544 218888 3596
rect 218940 3544 218946 3596
rect 224954 3544 224960 3596
rect 225012 3584 225018 3596
rect 225012 3556 225092 3584
rect 225012 3544 225018 3556
rect 212534 3476 212540 3528
rect 212592 3516 212598 3528
rect 212629 3519 212687 3525
rect 212629 3516 212641 3519
rect 212592 3488 212641 3516
rect 212592 3476 212598 3488
rect 212629 3485 212641 3488
rect 212675 3485 212687 3519
rect 212629 3479 212687 3485
rect 213362 3476 213368 3528
rect 213420 3476 213426 3528
rect 213454 3476 213460 3528
rect 213512 3525 213518 3528
rect 213512 3519 213540 3525
rect 213528 3485 213540 3519
rect 213512 3479 213540 3485
rect 213512 3476 213518 3479
rect 213638 3476 213644 3528
rect 213696 3476 213702 3528
rect 215386 3476 215392 3528
rect 215444 3476 215450 3528
rect 216398 3476 216404 3528
rect 216456 3476 216462 3528
rect 217226 3476 217232 3528
rect 217284 3516 217290 3528
rect 217505 3519 217563 3525
rect 217505 3516 217517 3519
rect 217284 3488 217517 3516
rect 217284 3476 217290 3488
rect 217505 3485 217517 3488
rect 217551 3485 217563 3519
rect 217505 3479 217563 3485
rect 219158 3476 219164 3528
rect 219216 3516 219222 3528
rect 219216 3488 221872 3516
rect 219216 3476 219222 3488
rect 212350 3408 212356 3460
rect 212408 3408 212414 3460
rect 217689 3451 217747 3457
rect 217336 3420 217640 3448
rect 214285 3383 214343 3389
rect 214285 3380 214297 3383
rect 210436 3352 214297 3380
rect 214285 3349 214297 3352
rect 214331 3349 214343 3383
rect 214285 3343 214343 3349
rect 214653 3383 214711 3389
rect 214653 3349 214665 3383
rect 214699 3380 214711 3383
rect 215846 3380 215852 3392
rect 214699 3352 215852 3380
rect 214699 3349 214711 3352
rect 214653 3343 214711 3349
rect 215846 3340 215852 3352
rect 215904 3340 215910 3392
rect 216490 3340 216496 3392
rect 216548 3380 216554 3392
rect 217336 3380 217364 3420
rect 216548 3352 217364 3380
rect 216548 3340 216554 3352
rect 217410 3340 217416 3392
rect 217468 3340 217474 3392
rect 217612 3380 217640 3420
rect 217689 3417 217701 3451
rect 217735 3448 217747 3451
rect 220170 3448 220176 3460
rect 217735 3420 220176 3448
rect 217735 3417 217747 3420
rect 217689 3411 217747 3417
rect 220170 3408 220176 3420
rect 220228 3408 220234 3460
rect 221844 3448 221872 3488
rect 222746 3476 222752 3528
rect 222804 3476 222810 3528
rect 225064 3516 225092 3556
rect 225138 3544 225144 3596
rect 225196 3584 225202 3596
rect 225509 3587 225567 3593
rect 225509 3584 225521 3587
rect 225196 3556 225521 3584
rect 225196 3544 225202 3556
rect 225509 3553 225521 3556
rect 225555 3553 225567 3587
rect 226150 3584 226156 3596
rect 225509 3547 225567 3553
rect 225616 3556 226156 3584
rect 225616 3516 225644 3556
rect 226150 3544 226156 3556
rect 226208 3544 226214 3596
rect 226567 3587 226625 3593
rect 226567 3553 226579 3587
rect 226613 3584 226625 3587
rect 227714 3584 227720 3596
rect 226613 3556 227720 3584
rect 226613 3553 226625 3556
rect 226567 3547 226625 3553
rect 227714 3544 227720 3556
rect 227772 3544 227778 3596
rect 228008 3556 234614 3584
rect 225064 3488 225644 3516
rect 225690 3476 225696 3528
rect 225748 3476 225754 3528
rect 226426 3476 226432 3528
rect 226484 3476 226490 3528
rect 226702 3476 226708 3528
rect 226760 3476 226766 3528
rect 228008 3516 228036 3556
rect 227640 3488 228036 3516
rect 230661 3519 230719 3525
rect 225598 3448 225604 3460
rect 221844 3420 225604 3448
rect 225598 3408 225604 3420
rect 225656 3408 225662 3460
rect 227640 3380 227668 3488
rect 230661 3485 230673 3519
rect 230707 3516 230719 3519
rect 231486 3516 231492 3528
rect 230707 3488 231492 3516
rect 230707 3485 230719 3488
rect 230661 3479 230719 3485
rect 231486 3476 231492 3488
rect 231544 3476 231550 3528
rect 234586 3516 234614 3556
rect 242894 3544 242900 3596
rect 242952 3584 242958 3596
rect 253934 3584 253940 3596
rect 242952 3556 253940 3584
rect 242952 3544 242958 3556
rect 253934 3544 253940 3556
rect 253992 3544 253998 3596
rect 259273 3587 259331 3593
rect 259273 3553 259285 3587
rect 259319 3584 259331 3587
rect 268102 3584 268108 3596
rect 259319 3556 268108 3584
rect 259319 3553 259331 3556
rect 259273 3547 259331 3553
rect 268102 3544 268108 3556
rect 268160 3544 268166 3596
rect 248966 3516 248972 3528
rect 234586 3488 248972 3516
rect 248966 3476 248972 3488
rect 249024 3476 249030 3528
rect 251910 3476 251916 3528
rect 251968 3516 251974 3528
rect 252097 3519 252155 3525
rect 252097 3516 252109 3519
rect 251968 3488 252109 3516
rect 251968 3476 251974 3488
rect 252097 3485 252109 3488
rect 252143 3485 252155 3519
rect 252097 3479 252155 3485
rect 258074 3476 258080 3528
rect 258132 3476 258138 3528
rect 258258 3476 258264 3528
rect 258316 3516 258322 3528
rect 258997 3519 259055 3525
rect 258997 3516 259009 3519
rect 258316 3488 259009 3516
rect 258316 3476 258322 3488
rect 258997 3485 259009 3488
rect 259043 3485 259055 3519
rect 260834 3516 260840 3528
rect 258997 3479 259055 3485
rect 259840 3488 260840 3516
rect 229186 3408 229192 3460
rect 229244 3448 229250 3460
rect 251450 3448 251456 3460
rect 229244 3420 251456 3448
rect 229244 3408 229250 3420
rect 251450 3408 251456 3420
rect 251508 3408 251514 3460
rect 256421 3451 256479 3457
rect 256421 3448 256433 3451
rect 252296 3420 256433 3448
rect 217612 3352 227668 3380
rect 227714 3340 227720 3392
rect 227772 3380 227778 3392
rect 229830 3380 229836 3392
rect 227772 3352 229836 3380
rect 227772 3340 227778 3352
rect 229830 3340 229836 3352
rect 229888 3340 229894 3392
rect 230750 3340 230756 3392
rect 230808 3380 230814 3392
rect 230845 3383 230903 3389
rect 230845 3380 230857 3383
rect 230808 3352 230857 3380
rect 230808 3340 230814 3352
rect 230845 3349 230857 3352
rect 230891 3349 230903 3383
rect 230845 3343 230903 3349
rect 242986 3340 242992 3392
rect 243044 3380 243050 3392
rect 252296 3380 252324 3420
rect 256421 3417 256433 3420
rect 256467 3448 256479 3451
rect 257614 3448 257620 3460
rect 256467 3420 257620 3448
rect 256467 3417 256479 3420
rect 256421 3411 256479 3417
rect 257614 3408 257620 3420
rect 257672 3408 257678 3460
rect 258445 3451 258503 3457
rect 258445 3417 258457 3451
rect 258491 3448 258503 3451
rect 259840 3448 259868 3488
rect 260834 3476 260840 3488
rect 260892 3476 260898 3528
rect 265529 3519 265587 3525
rect 265529 3485 265541 3519
rect 265575 3516 265587 3519
rect 266078 3516 266084 3528
rect 265575 3488 266084 3516
rect 265575 3485 265587 3488
rect 265529 3479 265587 3485
rect 266078 3476 266084 3488
rect 266136 3476 266142 3528
rect 266170 3476 266176 3528
rect 266228 3476 266234 3528
rect 267366 3476 267372 3528
rect 267424 3476 267430 3528
rect 267734 3476 267740 3528
rect 267792 3516 267798 3528
rect 268013 3519 268071 3525
rect 267792 3488 267964 3516
rect 267792 3476 267798 3488
rect 258491 3420 259868 3448
rect 259917 3451 259975 3457
rect 258491 3417 258503 3420
rect 258445 3411 258503 3417
rect 259917 3417 259929 3451
rect 259963 3448 259975 3451
rect 260006 3448 260012 3460
rect 259963 3420 260012 3448
rect 259963 3417 259975 3420
rect 259917 3411 259975 3417
rect 260006 3408 260012 3420
rect 260064 3408 260070 3460
rect 260285 3451 260343 3457
rect 260285 3417 260297 3451
rect 260331 3448 260343 3451
rect 267642 3448 267648 3460
rect 260331 3420 267648 3448
rect 260331 3417 260343 3420
rect 260285 3411 260343 3417
rect 267642 3408 267648 3420
rect 267700 3408 267706 3460
rect 267936 3448 267964 3488
rect 268013 3485 268025 3519
rect 268059 3512 268071 3519
rect 268194 3516 268200 3528
rect 268120 3512 268200 3516
rect 268059 3488 268200 3512
rect 268059 3485 268148 3488
rect 268013 3484 268148 3485
rect 268013 3479 268071 3484
rect 268194 3476 268200 3488
rect 268252 3476 268258 3528
rect 268657 3519 268715 3525
rect 268657 3485 268669 3519
rect 268703 3516 268715 3519
rect 268746 3516 268752 3528
rect 268703 3488 268752 3516
rect 268703 3485 268715 3488
rect 268657 3479 268715 3485
rect 268746 3476 268752 3488
rect 268804 3476 268810 3528
rect 269874 3525 269902 3612
rect 269117 3519 269175 3525
rect 269117 3516 269129 3519
rect 268856 3488 269129 3516
rect 268856 3448 268884 3488
rect 269117 3485 269129 3488
rect 269163 3485 269175 3519
rect 269117 3479 269175 3485
rect 269853 3519 269911 3525
rect 269853 3485 269865 3519
rect 269899 3485 269911 3519
rect 269853 3479 269911 3485
rect 269942 3476 269948 3528
rect 270000 3516 270006 3528
rect 270589 3519 270647 3525
rect 270589 3516 270601 3519
rect 270000 3488 270601 3516
rect 270000 3476 270006 3488
rect 270589 3485 270601 3488
rect 270635 3485 270647 3519
rect 270589 3479 270647 3485
rect 267936 3420 268884 3448
rect 269022 3408 269028 3460
rect 269080 3448 269086 3460
rect 271966 3448 271972 3460
rect 269080 3420 271972 3448
rect 269080 3408 269086 3420
rect 271966 3408 271972 3420
rect 272024 3408 272030 3460
rect 243044 3352 252324 3380
rect 243044 3340 243050 3352
rect 252370 3340 252376 3392
rect 252428 3340 252434 3392
rect 257632 3380 257660 3408
rect 258721 3383 258779 3389
rect 258721 3380 258733 3383
rect 257632 3352 258733 3380
rect 258721 3349 258733 3352
rect 258767 3380 258779 3383
rect 259641 3383 259699 3389
rect 259641 3380 259653 3383
rect 258767 3352 259653 3380
rect 258767 3349 258779 3352
rect 258721 3343 258779 3349
rect 259641 3349 259653 3352
rect 259687 3349 259699 3383
rect 259641 3343 259699 3349
rect 265618 3340 265624 3392
rect 265676 3380 265682 3392
rect 267734 3380 267740 3392
rect 265676 3352 267740 3380
rect 265676 3340 265682 3352
rect 267734 3340 267740 3352
rect 267792 3340 267798 3392
rect 267829 3383 267887 3389
rect 267829 3349 267841 3383
rect 267875 3380 267887 3383
rect 270034 3380 270040 3392
rect 267875 3352 270040 3380
rect 267875 3349 267887 3352
rect 267829 3343 267887 3349
rect 270034 3340 270040 3352
rect 270092 3340 270098 3392
rect 1104 3290 271651 3312
rect 1104 3238 68546 3290
rect 68598 3238 68610 3290
rect 68662 3238 68674 3290
rect 68726 3238 68738 3290
rect 68790 3238 68802 3290
rect 68854 3238 136143 3290
rect 136195 3238 136207 3290
rect 136259 3238 136271 3290
rect 136323 3238 136335 3290
rect 136387 3238 136399 3290
rect 136451 3238 203740 3290
rect 203792 3238 203804 3290
rect 203856 3238 203868 3290
rect 203920 3238 203932 3290
rect 203984 3238 203996 3290
rect 204048 3238 271337 3290
rect 271389 3238 271401 3290
rect 271453 3238 271465 3290
rect 271517 3238 271529 3290
rect 271581 3238 271593 3290
rect 271645 3238 271651 3290
rect 1104 3216 271651 3238
rect 27246 3136 27252 3188
rect 27304 3176 27310 3188
rect 37550 3176 37556 3188
rect 27304 3148 37556 3176
rect 27304 3136 27310 3148
rect 37550 3136 37556 3148
rect 37608 3136 37614 3188
rect 37660 3148 41414 3176
rect 26326 3108 26332 3120
rect 25332 3080 26332 3108
rect 23842 3000 23848 3052
rect 23900 3040 23906 3052
rect 24305 3043 24363 3049
rect 24305 3040 24317 3043
rect 23900 3012 24317 3040
rect 23900 3000 23906 3012
rect 24305 3009 24317 3012
rect 24351 3009 24363 3043
rect 24305 3003 24363 3009
rect 19242 2932 19248 2984
rect 19300 2972 19306 2984
rect 24854 2972 24860 2984
rect 19300 2944 24860 2972
rect 19300 2932 19306 2944
rect 24854 2932 24860 2944
rect 24912 2932 24918 2984
rect 24949 2975 25007 2981
rect 24949 2941 24961 2975
rect 24995 2972 25007 2975
rect 25222 2972 25228 2984
rect 24995 2944 25228 2972
rect 24995 2941 25007 2944
rect 24949 2935 25007 2941
rect 25222 2932 25228 2944
rect 25280 2932 25286 2984
rect 22922 2864 22928 2916
rect 22980 2904 22986 2916
rect 24489 2907 24547 2913
rect 24489 2904 24501 2907
rect 22980 2876 24501 2904
rect 22980 2864 22986 2876
rect 24489 2873 24501 2876
rect 24535 2873 24547 2907
rect 24489 2867 24547 2873
rect 19978 2796 19984 2848
rect 20036 2836 20042 2848
rect 25332 2836 25360 3080
rect 26326 3068 26332 3080
rect 26384 3068 26390 3120
rect 27062 3068 27068 3120
rect 27120 3108 27126 3120
rect 27120 3080 27384 3108
rect 27120 3068 27126 3080
rect 25406 3000 25412 3052
rect 25464 3040 25470 3052
rect 26142 3040 26148 3052
rect 25464 3012 26148 3040
rect 25464 3000 25470 3012
rect 26142 3000 26148 3012
rect 26200 3040 26206 3052
rect 26237 3043 26295 3049
rect 26237 3040 26249 3043
rect 26200 3012 26249 3040
rect 26200 3000 26206 3012
rect 26237 3009 26249 3012
rect 26283 3009 26295 3043
rect 26237 3003 26295 3009
rect 26050 2932 26056 2984
rect 26108 2972 26114 2984
rect 27356 2981 27384 3080
rect 27614 3068 27620 3120
rect 27672 3108 27678 3120
rect 35894 3108 35900 3120
rect 27672 3080 35900 3108
rect 27672 3068 27678 3080
rect 35894 3068 35900 3080
rect 35952 3068 35958 3120
rect 37660 3108 37688 3148
rect 36556 3080 37688 3108
rect 37829 3111 37887 3117
rect 27525 3043 27583 3049
rect 27525 3009 27537 3043
rect 27571 3040 27583 3043
rect 27890 3040 27896 3052
rect 27571 3012 27896 3040
rect 27571 3009 27583 3012
rect 27525 3003 27583 3009
rect 27890 3000 27896 3012
rect 27948 3000 27954 3052
rect 27982 3000 27988 3052
rect 28040 3000 28046 3052
rect 27341 2975 27399 2981
rect 26108 2944 27200 2972
rect 26108 2932 26114 2944
rect 20036 2808 25360 2836
rect 20036 2796 20042 2808
rect 25590 2796 25596 2848
rect 25648 2796 25654 2848
rect 26418 2796 26424 2848
rect 26476 2796 26482 2848
rect 27172 2836 27200 2944
rect 27341 2941 27353 2975
rect 27387 2941 27399 2975
rect 36556 2972 36584 3080
rect 37829 3077 37841 3111
rect 37875 3108 37887 3111
rect 38010 3108 38016 3120
rect 37875 3080 38016 3108
rect 37875 3077 37887 3080
rect 37829 3071 37887 3077
rect 38010 3068 38016 3080
rect 38068 3068 38074 3120
rect 38102 3068 38108 3120
rect 38160 3068 38166 3120
rect 38194 3068 38200 3120
rect 38252 3068 38258 3120
rect 38562 3068 38568 3120
rect 38620 3068 38626 3120
rect 38930 3068 38936 3120
rect 38988 3068 38994 3120
rect 39850 3068 39856 3120
rect 39908 3068 39914 3120
rect 40126 3068 40132 3120
rect 40184 3068 40190 3120
rect 40494 3068 40500 3120
rect 40552 3108 40558 3120
rect 40589 3111 40647 3117
rect 40589 3108 40601 3111
rect 40552 3080 40601 3108
rect 40552 3068 40558 3080
rect 40589 3077 40601 3080
rect 40635 3077 40647 3111
rect 40589 3071 40647 3077
rect 40957 3111 41015 3117
rect 40957 3077 40969 3111
rect 41003 3108 41015 3111
rect 41046 3108 41052 3120
rect 41003 3080 41052 3108
rect 41003 3077 41015 3080
rect 40957 3071 41015 3077
rect 41046 3068 41052 3080
rect 41104 3068 41110 3120
rect 37182 3000 37188 3052
rect 37240 3040 37246 3052
rect 38470 3040 38476 3052
rect 37240 3012 38476 3040
rect 37240 3000 37246 3012
rect 38470 3000 38476 3012
rect 38528 3040 38534 3052
rect 39942 3040 39948 3052
rect 38528 3012 39948 3040
rect 38528 3000 38534 3012
rect 27341 2935 27399 2941
rect 27540 2944 36584 2972
rect 38856 2958 38884 3012
rect 39942 3000 39948 3012
rect 40000 3000 40006 3052
rect 40218 3000 40224 3052
rect 40276 3000 40282 3052
rect 40770 3000 40776 3052
rect 40828 3000 40834 3052
rect 41386 3040 41414 3148
rect 52270 3136 52276 3188
rect 52328 3176 52334 3188
rect 81434 3176 81440 3188
rect 52328 3148 81440 3176
rect 52328 3136 52334 3148
rect 81434 3136 81440 3148
rect 81492 3136 81498 3188
rect 83277 3179 83335 3185
rect 83277 3145 83289 3179
rect 83323 3176 83335 3179
rect 84013 3179 84071 3185
rect 84013 3176 84025 3179
rect 83323 3148 84025 3176
rect 83323 3145 83335 3148
rect 83277 3139 83335 3145
rect 84013 3145 84025 3148
rect 84059 3176 84071 3179
rect 98638 3176 98644 3188
rect 84059 3148 98644 3176
rect 84059 3145 84071 3148
rect 84013 3139 84071 3145
rect 41874 3068 41880 3120
rect 41932 3108 41938 3120
rect 86034 3108 86040 3120
rect 41932 3080 86040 3108
rect 41932 3068 41938 3080
rect 86034 3068 86040 3080
rect 86092 3068 86098 3120
rect 86144 3117 86172 3148
rect 98638 3136 98644 3148
rect 98696 3136 98702 3188
rect 98730 3136 98736 3188
rect 98788 3136 98794 3188
rect 101490 3136 101496 3188
rect 101548 3136 101554 3188
rect 102042 3136 102048 3188
rect 102100 3176 102106 3188
rect 102100 3148 103376 3176
rect 102100 3136 102106 3148
rect 86129 3111 86187 3117
rect 86129 3077 86141 3111
rect 86175 3077 86187 3111
rect 96617 3111 96675 3117
rect 96617 3108 96629 3111
rect 86129 3071 86187 3077
rect 88352 3080 96629 3108
rect 54110 3040 54116 3052
rect 41386 3012 54116 3040
rect 54110 3000 54116 3012
rect 54168 3000 54174 3052
rect 82354 3000 82360 3052
rect 82412 3000 82418 3052
rect 86586 3000 86592 3052
rect 86644 3000 86650 3052
rect 40788 2958 40816 3000
rect 27249 2839 27307 2845
rect 27249 2836 27261 2839
rect 27172 2808 27261 2836
rect 27249 2805 27261 2808
rect 27295 2836 27307 2839
rect 27540 2836 27568 2944
rect 40954 2932 40960 2984
rect 41012 2972 41018 2984
rect 67542 2972 67548 2984
rect 41012 2944 67548 2972
rect 41012 2932 41018 2944
rect 67542 2932 67548 2944
rect 67600 2932 67606 2984
rect 82078 2932 82084 2984
rect 82136 2932 82142 2984
rect 84286 2932 84292 2984
rect 84344 2932 84350 2984
rect 84470 2932 84476 2984
rect 84528 2932 84534 2984
rect 86770 2932 86776 2984
rect 86828 2932 86834 2984
rect 28074 2864 28080 2916
rect 28132 2904 28138 2916
rect 28169 2907 28227 2913
rect 28169 2904 28181 2907
rect 28132 2876 28181 2904
rect 28132 2864 28138 2876
rect 28169 2873 28181 2876
rect 28215 2873 28227 2907
rect 28169 2867 28227 2873
rect 39114 2864 39120 2916
rect 39172 2864 39178 2916
rect 41138 2864 41144 2916
rect 41196 2864 41202 2916
rect 73154 2864 73160 2916
rect 73212 2904 73218 2916
rect 73212 2876 77294 2904
rect 73212 2864 73218 2876
rect 27295 2808 27568 2836
rect 27295 2805 27307 2808
rect 27249 2799 27307 2805
rect 27706 2796 27712 2848
rect 27764 2796 27770 2848
rect 30926 2796 30932 2848
rect 30984 2836 30990 2848
rect 37458 2836 37464 2848
rect 30984 2808 37464 2836
rect 30984 2796 30990 2808
rect 37458 2796 37464 2808
rect 37516 2796 37522 2848
rect 77266 2836 77294 2876
rect 88352 2836 88380 3080
rect 96617 3077 96629 3080
rect 96663 3108 96675 3111
rect 103348 3108 103376 3148
rect 106274 3136 106280 3188
rect 106332 3176 106338 3188
rect 106332 3148 132494 3176
rect 106332 3136 106338 3148
rect 109494 3108 109500 3120
rect 96663 3080 97120 3108
rect 103348 3080 109500 3108
rect 96663 3077 96675 3080
rect 96617 3071 96675 3077
rect 89162 3000 89168 3052
rect 89220 3000 89226 3052
rect 91925 3043 91983 3049
rect 91925 3009 91937 3043
rect 91971 3040 91983 3043
rect 92290 3040 92296 3052
rect 91971 3012 92296 3040
rect 91971 3009 91983 3012
rect 91925 3003 91983 3009
rect 92290 3000 92296 3012
rect 92348 3000 92354 3052
rect 94222 3000 94228 3052
rect 94280 3000 94286 3052
rect 96062 3000 96068 3052
rect 96120 3000 96126 3052
rect 96890 3000 96896 3052
rect 96948 3000 96954 3052
rect 97092 3049 97120 3080
rect 109494 3068 109500 3080
rect 109552 3068 109558 3120
rect 110417 3111 110475 3117
rect 110417 3108 110429 3111
rect 109604 3080 110429 3108
rect 97077 3043 97135 3049
rect 97077 3009 97089 3043
rect 97123 3009 97135 3043
rect 97077 3003 97135 3009
rect 98086 3000 98092 3052
rect 98144 3000 98150 3052
rect 99650 3000 99656 3052
rect 99708 3000 99714 3052
rect 101674 3000 101680 3052
rect 101732 3000 101738 3052
rect 102615 3043 102673 3049
rect 102615 3040 102627 3043
rect 102612 3018 102627 3040
rect 88429 2975 88487 2981
rect 88429 2941 88441 2975
rect 88475 2941 88487 2975
rect 88429 2935 88487 2941
rect 88444 2904 88472 2935
rect 90082 2932 90088 2984
rect 90140 2932 90146 2984
rect 90266 2932 90272 2984
rect 90324 2972 90330 2984
rect 91646 2972 91652 2984
rect 90324 2944 91652 2972
rect 90324 2932 90330 2944
rect 91646 2932 91652 2944
rect 91704 2932 91710 2984
rect 93762 2972 93768 2984
rect 92216 2944 93768 2972
rect 88981 2907 89039 2913
rect 88981 2904 88993 2907
rect 88444 2876 88993 2904
rect 88981 2873 88993 2876
rect 89027 2904 89039 2907
rect 89806 2904 89812 2916
rect 89027 2876 89812 2904
rect 89027 2873 89039 2876
rect 88981 2867 89039 2873
rect 89806 2864 89812 2876
rect 89864 2864 89870 2916
rect 91664 2904 91692 2932
rect 92216 2904 92244 2944
rect 93762 2932 93768 2944
rect 93820 2972 93826 2984
rect 94409 2975 94467 2981
rect 94409 2972 94421 2975
rect 93820 2944 94421 2972
rect 93820 2932 93826 2944
rect 94409 2941 94421 2944
rect 94455 2941 94467 2975
rect 94409 2935 94467 2941
rect 97166 2932 97172 2984
rect 97224 2972 97230 2984
rect 97813 2975 97871 2981
rect 97813 2972 97825 2975
rect 97224 2944 97825 2972
rect 97224 2932 97230 2944
rect 97813 2941 97825 2944
rect 97859 2941 97871 2975
rect 97813 2935 97871 2941
rect 97951 2975 98009 2981
rect 97951 2941 97963 2975
rect 97997 2972 98009 2975
rect 99466 2972 99472 2984
rect 97997 2944 99472 2972
rect 97997 2941 98009 2944
rect 97951 2935 98009 2941
rect 99466 2932 99472 2944
rect 99524 2932 99530 2984
rect 99834 2932 99840 2984
rect 99892 2932 99898 2984
rect 100386 2932 100392 2984
rect 100444 2972 100450 2984
rect 100573 2975 100631 2981
rect 100573 2972 100585 2975
rect 100444 2944 100585 2972
rect 100444 2932 100450 2944
rect 100573 2941 100585 2944
rect 100619 2941 100631 2975
rect 100573 2935 100631 2941
rect 100662 2932 100668 2984
rect 100720 2981 100726 2984
rect 100720 2975 100748 2981
rect 100736 2941 100748 2975
rect 100720 2935 100748 2941
rect 100849 2975 100907 2981
rect 100849 2941 100861 2975
rect 100895 2972 100907 2975
rect 101398 2972 101404 2984
rect 100895 2944 101404 2972
rect 100895 2941 100907 2944
rect 100849 2935 100907 2941
rect 100720 2932 100726 2935
rect 101398 2932 101404 2944
rect 101456 2932 101462 2984
rect 101858 2932 101864 2984
rect 101916 2932 101922 2984
rect 102226 2932 102232 2984
rect 102284 2972 102290 2984
rect 102321 2975 102379 2981
rect 102321 2972 102333 2975
rect 102284 2944 102333 2972
rect 102284 2932 102290 2944
rect 102321 2941 102333 2944
rect 102367 2941 102379 2975
rect 102594 2966 102600 3018
rect 102661 3009 102673 3043
rect 102652 3003 102673 3009
rect 102652 2966 102658 3003
rect 102870 3000 102876 3052
rect 102928 3000 102934 3052
rect 105832 3012 107056 3040
rect 102735 2975 102793 2981
rect 102321 2935 102379 2941
rect 102735 2941 102747 2975
rect 102781 2972 102793 2975
rect 103517 2975 103575 2981
rect 102781 2944 103468 2972
rect 102781 2941 102793 2944
rect 102735 2935 102793 2941
rect 91664 2876 92244 2904
rect 92290 2864 92296 2916
rect 92348 2864 92354 2916
rect 97537 2907 97595 2913
rect 97537 2873 97549 2907
rect 97583 2873 97595 2907
rect 97537 2867 97595 2873
rect 77266 2808 88380 2836
rect 89346 2796 89352 2848
rect 89404 2796 89410 2848
rect 89717 2839 89775 2845
rect 89717 2805 89729 2839
rect 89763 2836 89775 2839
rect 92308 2836 92336 2864
rect 89763 2808 92336 2836
rect 89763 2805 89775 2808
rect 89717 2799 89775 2805
rect 96798 2796 96804 2848
rect 96856 2836 96862 2848
rect 96982 2836 96988 2848
rect 96856 2808 96988 2836
rect 96856 2796 96862 2808
rect 96982 2796 96988 2808
rect 97040 2796 97046 2848
rect 97350 2796 97356 2848
rect 97408 2836 97414 2848
rect 97552 2836 97580 2867
rect 99926 2864 99932 2916
rect 99984 2904 99990 2916
rect 100297 2907 100355 2913
rect 100297 2904 100309 2907
rect 99984 2876 100309 2904
rect 99984 2864 99990 2876
rect 100297 2873 100309 2876
rect 100343 2873 100355 2907
rect 100297 2867 100355 2873
rect 99944 2836 99972 2864
rect 97408 2808 99972 2836
rect 100312 2836 100340 2867
rect 102244 2836 102272 2932
rect 103440 2904 103468 2944
rect 103517 2941 103529 2975
rect 103563 2972 103575 2975
rect 104437 2975 104495 2981
rect 104437 2972 104449 2975
rect 103563 2944 104449 2972
rect 103563 2941 103575 2944
rect 103517 2935 103575 2941
rect 104437 2941 104449 2944
rect 104483 2941 104495 2975
rect 104437 2935 104495 2941
rect 104618 2932 104624 2984
rect 104676 2972 104682 2984
rect 105832 2972 105860 3012
rect 104676 2944 105860 2972
rect 106277 2975 106335 2981
rect 104676 2932 104682 2944
rect 106277 2941 106289 2975
rect 106323 2941 106335 2975
rect 107028 2972 107056 3012
rect 107102 3000 107108 3052
rect 107160 3000 107166 3052
rect 109310 3000 109316 3052
rect 109368 3040 109374 3052
rect 109604 3040 109632 3080
rect 110417 3077 110429 3080
rect 110463 3077 110475 3111
rect 110417 3071 110475 3077
rect 112714 3068 112720 3120
rect 112772 3108 112778 3120
rect 116670 3108 116676 3120
rect 112772 3080 116676 3108
rect 112772 3068 112778 3080
rect 116670 3068 116676 3080
rect 116728 3068 116734 3120
rect 117682 3068 117688 3120
rect 117740 3108 117746 3120
rect 117740 3080 118694 3108
rect 117740 3068 117746 3080
rect 109368 3012 109632 3040
rect 109368 3000 109374 3012
rect 110230 3000 110236 3052
rect 110288 3000 110294 3052
rect 112073 3043 112131 3049
rect 112073 3009 112085 3043
rect 112119 3040 112131 3043
rect 115934 3040 115940 3052
rect 112119 3012 115940 3040
rect 112119 3009 112131 3012
rect 112073 3003 112131 3009
rect 107286 2972 107292 2984
rect 107028 2944 107292 2972
rect 106277 2935 106335 2941
rect 106182 2904 106188 2916
rect 103440 2876 106188 2904
rect 106182 2864 106188 2876
rect 106240 2864 106246 2916
rect 100312 2808 102272 2836
rect 97408 2796 97414 2808
rect 103330 2796 103336 2848
rect 103388 2836 103394 2848
rect 103885 2839 103943 2845
rect 103885 2836 103897 2839
rect 103388 2808 103897 2836
rect 103388 2796 103394 2808
rect 103885 2805 103897 2808
rect 103931 2836 103943 2839
rect 106292 2836 106320 2935
rect 107286 2932 107292 2944
rect 107344 2932 107350 2984
rect 107654 2932 107660 2984
rect 107712 2932 107718 2984
rect 109678 2932 109684 2984
rect 109736 2972 109742 2984
rect 112088 2972 112116 3003
rect 115934 3000 115940 3012
rect 115992 3000 115998 3052
rect 116118 3000 116124 3052
rect 116176 3000 116182 3052
rect 116486 3000 116492 3052
rect 116544 3000 116550 3052
rect 109736 2944 112116 2972
rect 109736 2932 109742 2944
rect 113542 2932 113548 2984
rect 113600 2972 113606 2984
rect 116136 2972 116164 3000
rect 113600 2944 116164 2972
rect 113600 2932 113606 2944
rect 116302 2932 116308 2984
rect 116360 2972 116366 2984
rect 116673 2975 116731 2981
rect 116673 2972 116685 2975
rect 116360 2944 116685 2972
rect 116360 2932 116366 2944
rect 116673 2941 116685 2944
rect 116719 2941 116731 2975
rect 116673 2935 116731 2941
rect 114646 2904 114652 2916
rect 109006 2876 114652 2904
rect 106553 2839 106611 2845
rect 106553 2836 106565 2839
rect 103931 2808 106565 2836
rect 103931 2805 103943 2808
rect 103885 2799 103943 2805
rect 106553 2805 106565 2808
rect 106599 2836 106611 2839
rect 109006 2836 109034 2876
rect 114646 2864 114652 2876
rect 114704 2864 114710 2916
rect 115750 2864 115756 2916
rect 115808 2904 115814 2916
rect 116121 2907 116179 2913
rect 116121 2904 116133 2907
rect 115808 2876 116133 2904
rect 115808 2864 115814 2876
rect 116121 2873 116133 2876
rect 116167 2873 116179 2907
rect 116688 2904 116716 2935
rect 116946 2932 116952 2984
rect 117004 2932 117010 2984
rect 117884 2904 117912 3080
rect 118666 2972 118694 3080
rect 120626 3068 120632 3120
rect 120684 3108 120690 3120
rect 120997 3111 121055 3117
rect 120997 3108 121009 3111
rect 120684 3080 121009 3108
rect 120684 3068 120690 3080
rect 120997 3077 121009 3080
rect 121043 3108 121055 3111
rect 123205 3111 123263 3117
rect 123205 3108 123217 3111
rect 121043 3080 123217 3108
rect 121043 3077 121055 3080
rect 120997 3071 121055 3077
rect 123205 3077 123217 3080
rect 123251 3108 123263 3111
rect 123481 3111 123539 3117
rect 123481 3108 123493 3111
rect 123251 3080 123493 3108
rect 123251 3077 123263 3080
rect 123205 3071 123263 3077
rect 123481 3077 123493 3080
rect 123527 3108 123539 3111
rect 123570 3108 123576 3120
rect 123527 3080 123576 3108
rect 123527 3077 123539 3080
rect 123481 3071 123539 3077
rect 123570 3068 123576 3080
rect 123628 3068 123634 3120
rect 120258 3000 120264 3052
rect 120316 3040 120322 3052
rect 121365 3043 121423 3049
rect 121365 3040 121377 3043
rect 120316 3012 121377 3040
rect 120316 3000 120322 3012
rect 121365 3009 121377 3012
rect 121411 3009 121423 3043
rect 121365 3003 121423 3009
rect 121549 2975 121607 2981
rect 121549 2972 121561 2975
rect 118666 2944 121561 2972
rect 121549 2941 121561 2944
rect 121595 2972 121607 2975
rect 121914 2972 121920 2984
rect 121595 2944 121920 2972
rect 121595 2941 121607 2944
rect 121549 2935 121607 2941
rect 121914 2932 121920 2944
rect 121972 2932 121978 2984
rect 116688 2876 117912 2904
rect 116121 2867 116179 2873
rect 106599 2808 109034 2836
rect 116136 2836 116164 2867
rect 116946 2836 116952 2848
rect 116136 2808 116952 2836
rect 106599 2805 106611 2808
rect 106553 2799 106611 2805
rect 116946 2796 116952 2808
rect 117004 2836 117010 2848
rect 118697 2839 118755 2845
rect 118697 2836 118709 2839
rect 117004 2808 118709 2836
rect 117004 2796 117010 2808
rect 118697 2805 118709 2808
rect 118743 2836 118755 2839
rect 124306 2836 124312 2848
rect 118743 2808 124312 2836
rect 118743 2805 118755 2808
rect 118697 2799 118755 2805
rect 124306 2796 124312 2808
rect 124364 2796 124370 2848
rect 132466 2836 132494 3148
rect 138934 3136 138940 3188
rect 138992 3176 138998 3188
rect 139581 3179 139639 3185
rect 139581 3176 139593 3179
rect 138992 3148 139593 3176
rect 138992 3136 138998 3148
rect 139581 3145 139593 3148
rect 139627 3145 139639 3179
rect 139581 3139 139639 3145
rect 141786 3136 141792 3188
rect 141844 3176 141850 3188
rect 144641 3179 144699 3185
rect 144641 3176 144653 3179
rect 141844 3148 144653 3176
rect 141844 3136 141850 3148
rect 144641 3145 144653 3148
rect 144687 3145 144699 3179
rect 144641 3139 144699 3145
rect 144822 3136 144828 3188
rect 144880 3176 144886 3188
rect 144880 3148 147352 3176
rect 144880 3136 144886 3148
rect 140685 3111 140743 3117
rect 140685 3108 140697 3111
rect 139504 3080 140697 3108
rect 137738 3000 137744 3052
rect 137796 3000 137802 3052
rect 138658 3000 138664 3052
rect 138716 3000 138722 3052
rect 137922 2932 137928 2984
rect 137980 2932 137986 2984
rect 138750 2932 138756 2984
rect 138808 2981 138814 2984
rect 138808 2975 138836 2981
rect 138824 2941 138836 2975
rect 138808 2935 138836 2941
rect 138808 2932 138814 2935
rect 138934 2932 138940 2984
rect 138992 2932 138998 2984
rect 139118 2932 139124 2984
rect 139176 2972 139182 2984
rect 139504 2972 139532 3080
rect 140685 3077 140697 3080
rect 140731 3108 140743 3111
rect 142154 3108 142160 3120
rect 140731 3080 142160 3108
rect 140731 3077 140743 3080
rect 140685 3071 140743 3077
rect 142154 3068 142160 3080
rect 142212 3068 142218 3120
rect 147324 3108 147352 3148
rect 147490 3136 147496 3188
rect 147548 3136 147554 3188
rect 148134 3136 148140 3188
rect 148192 3176 148198 3188
rect 148192 3148 149744 3176
rect 148192 3136 148198 3148
rect 148042 3108 148048 3120
rect 147324 3080 148048 3108
rect 148042 3068 148048 3080
rect 148100 3068 148106 3120
rect 141878 3000 141884 3052
rect 141936 3040 141942 3052
rect 142985 3043 143043 3049
rect 142985 3040 142997 3043
rect 141936 3012 142997 3040
rect 141936 3000 141942 3012
rect 142985 3009 142997 3012
rect 143031 3009 143043 3043
rect 142985 3003 143043 3009
rect 143718 3000 143724 3052
rect 143776 3000 143782 3052
rect 145837 3043 145895 3049
rect 145837 3040 145849 3043
rect 144564 3012 145849 3040
rect 139176 2944 139532 2972
rect 140501 2975 140559 2981
rect 139176 2932 139182 2944
rect 140501 2941 140513 2975
rect 140547 2941 140559 2975
rect 140501 2935 140559 2941
rect 140961 2975 141019 2981
rect 140961 2941 140973 2975
rect 141007 2941 141019 2975
rect 140961 2935 141019 2941
rect 138382 2864 138388 2916
rect 138440 2864 138446 2916
rect 140516 2904 140544 2935
rect 140774 2904 140780 2916
rect 140516 2876 140780 2904
rect 140774 2864 140780 2876
rect 140832 2864 140838 2916
rect 139857 2839 139915 2845
rect 139857 2836 139869 2839
rect 132466 2808 139869 2836
rect 139857 2805 139869 2808
rect 139903 2836 139915 2839
rect 140976 2836 141004 2935
rect 142706 2932 142712 2984
rect 142764 2972 142770 2984
rect 142801 2975 142859 2981
rect 142801 2972 142813 2975
rect 142764 2944 142813 2972
rect 142764 2932 142770 2944
rect 142801 2941 142813 2944
rect 142847 2941 142859 2975
rect 142801 2935 142859 2941
rect 143442 2932 143448 2984
rect 143500 2932 143506 2984
rect 143902 2981 143908 2984
rect 143859 2975 143908 2981
rect 143859 2941 143871 2975
rect 143905 2941 143908 2975
rect 143859 2935 143908 2941
rect 143902 2932 143908 2935
rect 143960 2932 143966 2984
rect 143994 2932 144000 2984
rect 144052 2932 144058 2984
rect 144362 2932 144368 2984
rect 144420 2972 144426 2984
rect 144564 2972 144592 3012
rect 145837 3009 145849 3012
rect 145883 3009 145895 3043
rect 145837 3003 145895 3009
rect 146570 3000 146576 3052
rect 146628 3000 146634 3052
rect 146846 3000 146852 3052
rect 146904 3000 146910 3052
rect 147766 3000 147772 3052
rect 147824 3040 147830 3052
rect 147953 3043 148011 3049
rect 147953 3040 147965 3043
rect 147824 3012 147965 3040
rect 147824 3000 147830 3012
rect 147953 3009 147965 3012
rect 147999 3009 148011 3043
rect 147953 3003 148011 3009
rect 148870 3000 148876 3052
rect 148928 3000 148934 3052
rect 149146 3000 149152 3052
rect 149204 3000 149210 3052
rect 144420 2944 144592 2972
rect 144420 2932 144426 2944
rect 145558 2932 145564 2984
rect 145616 2972 145622 2984
rect 146754 2981 146760 2984
rect 145653 2975 145711 2981
rect 145653 2972 145665 2975
rect 145616 2944 145665 2972
rect 145616 2932 145622 2944
rect 145653 2941 145665 2944
rect 145699 2941 145711 2975
rect 145653 2935 145711 2941
rect 146711 2975 146760 2981
rect 146711 2941 146723 2975
rect 146757 2941 146760 2975
rect 146711 2935 146760 2941
rect 146754 2932 146760 2935
rect 146812 2932 146818 2984
rect 148134 2932 148140 2984
rect 148192 2932 148198 2984
rect 148597 2975 148655 2981
rect 148597 2941 148609 2975
rect 148643 2972 148655 2975
rect 148686 2972 148692 2984
rect 148643 2944 148692 2972
rect 148643 2941 148655 2944
rect 148597 2935 148655 2941
rect 142617 2839 142675 2845
rect 142617 2836 142629 2839
rect 139903 2808 142629 2836
rect 139903 2805 139915 2808
rect 139857 2799 139915 2805
rect 142617 2805 142629 2808
rect 142663 2836 142675 2839
rect 142706 2836 142712 2848
rect 142663 2808 142712 2836
rect 142663 2805 142675 2808
rect 142617 2799 142675 2805
rect 142706 2796 142712 2808
rect 142764 2796 142770 2848
rect 143460 2836 143488 2932
rect 146297 2907 146355 2913
rect 146297 2873 146309 2907
rect 146343 2873 146355 2907
rect 146297 2867 146355 2873
rect 147416 2876 147674 2904
rect 144822 2836 144828 2848
rect 143460 2808 144828 2836
rect 144822 2796 144828 2808
rect 144880 2796 144886 2848
rect 146312 2836 146340 2867
rect 147416 2836 147444 2876
rect 146312 2808 147444 2836
rect 147646 2836 147674 2876
rect 148612 2836 148640 2935
rect 148686 2932 148692 2944
rect 148744 2932 148750 2984
rect 148962 2932 148968 2984
rect 149020 2981 149026 2984
rect 149020 2975 149048 2981
rect 149036 2941 149048 2975
rect 149020 2935 149048 2941
rect 149020 2932 149026 2935
rect 149716 2904 149744 3148
rect 150986 3136 150992 3188
rect 151044 3176 151050 3188
rect 151044 3148 195974 3176
rect 151044 3136 151050 3148
rect 152918 3068 152924 3120
rect 152976 3108 152982 3120
rect 156138 3108 156144 3120
rect 152976 3080 156144 3108
rect 152976 3068 152982 3080
rect 155954 3000 155960 3052
rect 156012 3000 156018 3052
rect 156064 3040 156092 3080
rect 156138 3068 156144 3080
rect 156196 3068 156202 3120
rect 157797 3111 157855 3117
rect 157797 3077 157809 3111
rect 157843 3108 157855 3111
rect 157886 3108 157892 3120
rect 157843 3080 157892 3108
rect 157843 3077 157855 3080
rect 157797 3071 157855 3077
rect 157886 3068 157892 3080
rect 157944 3068 157950 3120
rect 159729 3111 159787 3117
rect 159729 3077 159741 3111
rect 159775 3108 159787 3111
rect 160830 3108 160836 3120
rect 159775 3080 160836 3108
rect 159775 3077 159787 3080
rect 159729 3071 159787 3077
rect 160830 3068 160836 3080
rect 160888 3068 160894 3120
rect 162670 3108 162676 3120
rect 161032 3080 162676 3108
rect 156064 3012 156276 3040
rect 149793 2975 149851 2981
rect 149793 2941 149805 2975
rect 149839 2972 149851 2975
rect 150805 2975 150863 2981
rect 150805 2972 150817 2975
rect 149839 2944 150817 2972
rect 149839 2941 149851 2944
rect 149793 2935 149851 2941
rect 150805 2941 150817 2944
rect 150851 2941 150863 2975
rect 150805 2935 150863 2941
rect 150989 2975 151047 2981
rect 150989 2941 151001 2975
rect 151035 2941 151047 2975
rect 151265 2975 151323 2981
rect 151265 2972 151277 2975
rect 150989 2935 151047 2941
rect 151188 2944 151277 2972
rect 151004 2904 151032 2935
rect 149716 2876 151032 2904
rect 147646 2808 148640 2836
rect 149238 2796 149244 2848
rect 149296 2836 149302 2848
rect 151188 2836 151216 2944
rect 151265 2941 151277 2944
rect 151311 2941 151323 2975
rect 151265 2935 151323 2941
rect 156138 2932 156144 2984
rect 156196 2932 156202 2984
rect 156248 2972 156276 3012
rect 156874 3000 156880 3052
rect 156932 3000 156938 3052
rect 156966 3000 156972 3052
rect 157024 3049 157030 3052
rect 157024 3043 157052 3049
rect 157040 3009 157052 3043
rect 157024 3003 157052 3009
rect 157812 3012 158208 3040
rect 157024 3000 157030 3003
rect 157153 2975 157211 2981
rect 157153 2972 157165 2975
rect 156248 2944 157165 2972
rect 157153 2941 157165 2944
rect 157199 2972 157211 2975
rect 157812 2972 157840 3012
rect 157199 2944 157840 2972
rect 157889 2975 157947 2981
rect 157199 2941 157211 2944
rect 157153 2935 157211 2941
rect 157889 2941 157901 2975
rect 157935 2972 157947 2975
rect 157978 2972 157984 2984
rect 157935 2944 157984 2972
rect 157935 2941 157947 2944
rect 157889 2935 157947 2941
rect 157978 2932 157984 2944
rect 158036 2932 158042 2984
rect 158073 2975 158131 2981
rect 158073 2941 158085 2975
rect 158119 2941 158131 2975
rect 158180 2972 158208 3012
rect 158806 3000 158812 3052
rect 158864 3000 158870 3052
rect 158898 3000 158904 3052
rect 158956 3049 158962 3052
rect 158956 3043 158984 3049
rect 158972 3009 158984 3043
rect 158956 3003 158984 3009
rect 158956 3000 158962 3003
rect 160186 3000 160192 3052
rect 160244 3040 160250 3052
rect 160554 3040 160560 3052
rect 160244 3012 160560 3040
rect 160244 3000 160250 3012
rect 160554 3000 160560 3012
rect 160612 3040 160618 3052
rect 161032 3040 161060 3080
rect 162670 3068 162676 3080
rect 162728 3108 162734 3120
rect 175918 3108 175924 3120
rect 162728 3080 175924 3108
rect 162728 3068 162734 3080
rect 175918 3068 175924 3080
rect 175976 3068 175982 3120
rect 195946 3108 195974 3148
rect 204898 3136 204904 3188
rect 204956 3176 204962 3188
rect 211893 3179 211951 3185
rect 211893 3176 211905 3179
rect 204956 3148 211905 3176
rect 204956 3136 204962 3148
rect 211893 3145 211905 3148
rect 211939 3145 211951 3179
rect 211893 3139 211951 3145
rect 213362 3136 213368 3188
rect 213420 3176 213426 3188
rect 213914 3176 213920 3188
rect 213420 3148 213920 3176
rect 213420 3136 213426 3148
rect 213914 3136 213920 3148
rect 213972 3136 213978 3188
rect 214466 3136 214472 3188
rect 214524 3136 214530 3188
rect 214837 3179 214895 3185
rect 214837 3145 214849 3179
rect 214883 3176 214895 3179
rect 216030 3176 216036 3188
rect 214883 3148 216036 3176
rect 214883 3145 214895 3148
rect 214837 3139 214895 3145
rect 216030 3136 216036 3148
rect 216088 3136 216094 3188
rect 217226 3136 217232 3188
rect 217284 3136 217290 3188
rect 218698 3136 218704 3188
rect 218756 3136 218762 3188
rect 223853 3179 223911 3185
rect 218808 3148 221688 3176
rect 207934 3108 207940 3120
rect 195946 3080 207940 3108
rect 207934 3068 207940 3080
rect 207992 3068 207998 3120
rect 218054 3068 218060 3120
rect 218112 3108 218118 3120
rect 218808 3108 218836 3148
rect 218112 3080 218836 3108
rect 218112 3068 218118 3080
rect 218882 3068 218888 3120
rect 218940 3108 218946 3120
rect 221660 3108 221688 3148
rect 223853 3145 223865 3179
rect 223899 3176 223911 3179
rect 225690 3176 225696 3188
rect 223899 3148 225696 3176
rect 223899 3145 223911 3148
rect 223853 3139 223911 3145
rect 225690 3136 225696 3148
rect 225748 3136 225754 3188
rect 226242 3136 226248 3188
rect 226300 3176 226306 3188
rect 246206 3176 246212 3188
rect 226300 3148 246212 3176
rect 226300 3136 226306 3148
rect 246206 3136 246212 3148
rect 246264 3136 246270 3188
rect 252370 3136 252376 3188
rect 252428 3176 252434 3188
rect 262214 3176 262220 3188
rect 252428 3148 262220 3176
rect 252428 3136 252434 3148
rect 262214 3136 262220 3148
rect 262272 3136 262278 3188
rect 264054 3136 264060 3188
rect 264112 3176 264118 3188
rect 268470 3176 268476 3188
rect 264112 3148 268476 3176
rect 264112 3136 264118 3148
rect 268470 3136 268476 3148
rect 268528 3136 268534 3188
rect 268565 3179 268623 3185
rect 268565 3145 268577 3179
rect 268611 3176 268623 3179
rect 269298 3176 269304 3188
rect 268611 3148 269304 3176
rect 268611 3145 268623 3148
rect 268565 3139 268623 3145
rect 269298 3136 269304 3148
rect 269356 3136 269362 3188
rect 269942 3176 269948 3188
rect 269408 3148 269948 3176
rect 225969 3111 226027 3117
rect 225969 3108 225981 3111
rect 218940 3080 221596 3108
rect 221660 3080 225981 3108
rect 218940 3068 218946 3080
rect 160612 3012 161060 3040
rect 161201 3043 161259 3049
rect 160612 3000 160618 3012
rect 161201 3009 161213 3043
rect 161247 3040 161259 3043
rect 162026 3040 162032 3052
rect 161247 3012 162032 3040
rect 161247 3009 161259 3012
rect 161201 3003 161259 3009
rect 162026 3000 162032 3012
rect 162084 3000 162090 3052
rect 162946 3000 162952 3052
rect 163004 3000 163010 3052
rect 206005 3043 206063 3049
rect 206005 3009 206017 3043
rect 206051 3040 206063 3043
rect 207198 3040 207204 3052
rect 206051 3012 207204 3040
rect 206051 3009 206063 3012
rect 206005 3003 206063 3009
rect 159085 2975 159143 2981
rect 159085 2972 159097 2975
rect 158180 2944 159097 2972
rect 158073 2935 158131 2941
rect 159085 2941 159097 2944
rect 159131 2972 159143 2975
rect 159131 2944 159588 2972
rect 159131 2941 159143 2944
rect 159085 2935 159143 2941
rect 156598 2864 156604 2916
rect 156656 2864 156662 2916
rect 158088 2904 158116 2935
rect 159560 2916 159588 2944
rect 161290 2932 161296 2984
rect 161348 2972 161354 2984
rect 161569 2975 161627 2981
rect 161569 2972 161581 2975
rect 161348 2944 161581 2972
rect 161348 2932 161354 2944
rect 161569 2941 161581 2944
rect 161615 2941 161627 2975
rect 161569 2935 161627 2941
rect 167730 2932 167736 2984
rect 167788 2932 167794 2984
rect 202322 2932 202328 2984
rect 202380 2932 202386 2984
rect 204165 2975 204223 2981
rect 204165 2941 204177 2975
rect 204211 2972 204223 2975
rect 204349 2975 204407 2981
rect 204211 2944 204300 2972
rect 204211 2941 204223 2944
rect 204165 2935 204223 2941
rect 157720 2876 158116 2904
rect 158533 2907 158591 2913
rect 153102 2836 153108 2848
rect 149296 2808 153108 2836
rect 149296 2796 149302 2808
rect 153102 2796 153108 2808
rect 153160 2796 153166 2848
rect 156046 2796 156052 2848
rect 156104 2836 156110 2848
rect 157720 2836 157748 2876
rect 158533 2873 158545 2907
rect 158579 2904 158591 2907
rect 158622 2904 158628 2916
rect 158579 2876 158628 2904
rect 158579 2873 158591 2876
rect 158533 2867 158591 2873
rect 158622 2864 158628 2876
rect 158680 2864 158686 2916
rect 159542 2864 159548 2916
rect 159600 2864 159606 2916
rect 203794 2864 203800 2916
rect 203852 2864 203858 2916
rect 156104 2808 157748 2836
rect 156104 2796 156110 2808
rect 158346 2796 158352 2848
rect 158404 2836 158410 2848
rect 160646 2836 160652 2848
rect 158404 2808 160652 2836
rect 158404 2796 158410 2808
rect 160646 2796 160652 2808
rect 160704 2796 160710 2848
rect 163130 2796 163136 2848
rect 163188 2796 163194 2848
rect 204272 2836 204300 2944
rect 204349 2941 204361 2975
rect 204395 2972 204407 2975
rect 205082 2972 205088 2984
rect 204395 2944 205088 2972
rect 204395 2941 204407 2944
rect 204349 2935 204407 2941
rect 205082 2932 205088 2944
rect 205140 2932 205146 2984
rect 204438 2864 204444 2916
rect 204496 2904 204502 2916
rect 206020 2904 206048 3003
rect 207198 3000 207204 3012
rect 207256 3000 207262 3052
rect 207382 3000 207388 3052
rect 207440 3040 207446 3052
rect 207753 3043 207811 3049
rect 207753 3040 207765 3043
rect 207440 3012 207765 3040
rect 207440 3000 207446 3012
rect 207753 3009 207765 3012
rect 207799 3009 207811 3043
rect 207753 3003 207811 3009
rect 208670 3000 208676 3052
rect 208728 3000 208734 3052
rect 210970 3000 210976 3052
rect 211028 3000 211034 3052
rect 211062 3000 211068 3052
rect 211120 3049 211126 3052
rect 211120 3043 211148 3049
rect 211136 3009 211148 3043
rect 211120 3003 211148 3009
rect 211120 3000 211126 3003
rect 212166 3000 212172 3052
rect 212224 3040 212230 3052
rect 212629 3043 212687 3049
rect 212629 3040 212641 3043
rect 212224 3012 212641 3040
rect 212224 3000 212230 3012
rect 212629 3009 212641 3012
rect 212675 3009 212687 3043
rect 212629 3003 212687 3009
rect 213546 3000 213552 3052
rect 213604 3000 213610 3052
rect 213730 3049 213736 3052
rect 213687 3043 213736 3049
rect 213687 3009 213699 3043
rect 213733 3009 213736 3043
rect 213687 3003 213736 3009
rect 213730 3000 213736 3003
rect 213788 3000 213794 3052
rect 215573 3043 215631 3049
rect 215573 3040 215585 3043
rect 215266 3012 215585 3040
rect 206370 2932 206376 2984
rect 206428 2972 206434 2984
rect 207937 2975 207995 2981
rect 207937 2972 207949 2975
rect 206428 2944 207949 2972
rect 206428 2932 206434 2944
rect 207937 2941 207949 2944
rect 207983 2941 207995 2975
rect 207937 2935 207995 2941
rect 208394 2932 208400 2984
rect 208452 2932 208458 2984
rect 208854 2981 208860 2984
rect 208811 2975 208860 2981
rect 208811 2941 208823 2975
rect 208857 2941 208860 2975
rect 208811 2935 208860 2941
rect 208854 2932 208860 2935
rect 208912 2932 208918 2984
rect 208949 2975 209007 2981
rect 208949 2941 208961 2975
rect 208995 2972 209007 2975
rect 208995 2944 209544 2972
rect 208995 2941 209007 2944
rect 208949 2935 209007 2941
rect 204496 2876 206048 2904
rect 209516 2904 209544 2944
rect 209590 2932 209596 2984
rect 209648 2972 209654 2984
rect 210053 2975 210111 2981
rect 210053 2972 210065 2975
rect 209648 2944 210065 2972
rect 209648 2932 209654 2944
rect 210053 2941 210065 2944
rect 210099 2941 210111 2975
rect 210053 2935 210111 2941
rect 210234 2932 210240 2984
rect 210292 2932 210298 2984
rect 211246 2972 211252 2984
rect 210620 2944 211252 2972
rect 209516 2876 209774 2904
rect 204496 2864 204502 2876
rect 209593 2839 209651 2845
rect 209593 2836 209605 2839
rect 204272 2808 209605 2836
rect 209593 2805 209605 2808
rect 209639 2805 209651 2839
rect 209746 2836 209774 2876
rect 210620 2836 210648 2944
rect 211246 2932 211252 2944
rect 211304 2972 211310 2984
rect 211430 2972 211436 2984
rect 211304 2944 211436 2972
rect 211304 2932 211310 2944
rect 211430 2932 211436 2944
rect 211488 2972 211494 2984
rect 211488 2944 211660 2972
rect 211488 2932 211494 2944
rect 210697 2907 210755 2913
rect 210697 2873 210709 2907
rect 210743 2873 210755 2907
rect 211632 2904 211660 2944
rect 212810 2932 212816 2984
rect 212868 2932 212874 2984
rect 213825 2975 213883 2981
rect 213825 2972 213837 2975
rect 213196 2944 213837 2972
rect 213196 2904 213224 2944
rect 213825 2941 213837 2944
rect 213871 2972 213883 2975
rect 213871 2944 214328 2972
rect 213871 2941 213883 2944
rect 213825 2935 213883 2941
rect 211632 2876 213224 2904
rect 213273 2907 213331 2913
rect 210697 2867 210755 2873
rect 213273 2873 213285 2907
rect 213319 2873 213331 2907
rect 214300 2904 214328 2944
rect 214374 2932 214380 2984
rect 214432 2972 214438 2984
rect 215266 2972 215294 3012
rect 215573 3009 215585 3012
rect 215619 3009 215631 3043
rect 215573 3003 215631 3009
rect 216306 3000 216312 3052
rect 216364 3000 216370 3052
rect 216582 3000 216588 3052
rect 216640 3000 216646 3052
rect 221568 3049 221596 3080
rect 225969 3077 225981 3080
rect 226015 3077 226027 3111
rect 225969 3071 226027 3077
rect 226058 3068 226064 3120
rect 226116 3108 226122 3120
rect 226794 3108 226800 3120
rect 226116 3080 226800 3108
rect 226116 3068 226122 3080
rect 226794 3068 226800 3080
rect 226852 3068 226858 3120
rect 226978 3068 226984 3120
rect 227036 3108 227042 3120
rect 230382 3108 230388 3120
rect 227036 3080 230388 3108
rect 227036 3068 227042 3080
rect 230382 3068 230388 3080
rect 230440 3068 230446 3120
rect 259730 3068 259736 3120
rect 259788 3108 259794 3120
rect 259825 3111 259883 3117
rect 259825 3108 259837 3111
rect 259788 3080 259837 3108
rect 259788 3068 259794 3080
rect 259825 3077 259837 3080
rect 259871 3077 259883 3111
rect 259825 3071 259883 3077
rect 259914 3068 259920 3120
rect 259972 3108 259978 3120
rect 269408 3108 269436 3148
rect 269942 3136 269948 3148
rect 270000 3136 270006 3188
rect 271138 3136 271144 3188
rect 271196 3176 271202 3188
rect 271966 3176 271972 3188
rect 271196 3148 271972 3176
rect 271196 3136 271202 3148
rect 271966 3136 271972 3148
rect 272024 3136 272030 3188
rect 272058 3108 272064 3120
rect 259972 3080 269436 3108
rect 269776 3080 272064 3108
rect 259972 3068 259978 3080
rect 217965 3043 218023 3049
rect 217965 3009 217977 3043
rect 218011 3040 218023 3043
rect 221553 3043 221611 3049
rect 218011 3012 219112 3040
rect 218011 3009 218023 3012
rect 217965 3003 218023 3009
rect 219084 2984 219112 3012
rect 221553 3009 221565 3043
rect 221599 3009 221611 3043
rect 221553 3003 221611 3009
rect 222197 3043 222255 3049
rect 222197 3009 222209 3043
rect 222243 3040 222255 3043
rect 222933 3043 222991 3049
rect 222933 3040 222945 3043
rect 222243 3012 222945 3040
rect 222243 3009 222255 3012
rect 222197 3003 222255 3009
rect 222933 3009 222945 3012
rect 222979 3009 222991 3043
rect 222933 3003 222991 3009
rect 223206 3000 223212 3052
rect 223264 3000 223270 3052
rect 223298 3000 223304 3052
rect 223356 3040 223362 3052
rect 224037 3043 224095 3049
rect 224037 3040 224049 3043
rect 223356 3012 224049 3040
rect 223356 3000 223362 3012
rect 224037 3009 224049 3012
rect 224083 3009 224095 3043
rect 224037 3003 224095 3009
rect 226886 3000 226892 3052
rect 226944 3040 226950 3052
rect 227073 3043 227131 3049
rect 227073 3040 227085 3043
rect 226944 3012 227085 3040
rect 226944 3000 226950 3012
rect 227073 3009 227085 3012
rect 227119 3009 227131 3043
rect 227073 3003 227131 3009
rect 228082 3000 228088 3052
rect 228140 3000 228146 3052
rect 242526 3040 242532 3052
rect 234586 3012 242532 3040
rect 214432 2944 215294 2972
rect 215389 2975 215447 2981
rect 214432 2932 214438 2944
rect 215389 2941 215401 2975
rect 215435 2972 215447 2975
rect 215662 2972 215668 2984
rect 215435 2944 215668 2972
rect 215435 2941 215447 2944
rect 215389 2935 215447 2941
rect 215662 2932 215668 2944
rect 215720 2932 215726 2984
rect 215754 2932 215760 2984
rect 215812 2972 215818 2984
rect 216490 2981 216496 2984
rect 216033 2975 216091 2981
rect 216033 2972 216045 2975
rect 215812 2944 216045 2972
rect 215812 2932 215818 2944
rect 216033 2941 216045 2944
rect 216079 2941 216091 2975
rect 216033 2935 216091 2941
rect 216447 2975 216496 2981
rect 216447 2941 216459 2975
rect 216493 2941 216496 2975
rect 216447 2935 216496 2941
rect 216490 2932 216496 2935
rect 216548 2932 216554 2984
rect 216766 2932 216772 2984
rect 216824 2972 216830 2984
rect 217781 2975 217839 2981
rect 217781 2972 217793 2975
rect 216824 2944 217793 2972
rect 216824 2932 216830 2944
rect 217781 2941 217793 2944
rect 217827 2941 217839 2975
rect 217781 2935 217839 2941
rect 218146 2932 218152 2984
rect 218204 2972 218210 2984
rect 218885 2975 218943 2981
rect 218885 2972 218897 2975
rect 218204 2944 218897 2972
rect 218204 2932 218210 2944
rect 218885 2941 218897 2944
rect 218931 2941 218943 2975
rect 218885 2935 218943 2941
rect 219066 2932 219072 2984
rect 219124 2972 219130 2984
rect 220998 2972 221004 2984
rect 219124 2944 221004 2972
rect 219124 2932 219130 2944
rect 220998 2932 221004 2944
rect 221056 2972 221062 2984
rect 221737 2975 221795 2981
rect 221737 2972 221749 2975
rect 221056 2944 221749 2972
rect 221056 2932 221062 2944
rect 221737 2941 221749 2944
rect 221783 2972 221795 2975
rect 223574 2972 223580 2984
rect 221783 2944 223580 2972
rect 221783 2941 221795 2944
rect 221737 2935 221795 2941
rect 223574 2932 223580 2944
rect 223632 2972 223638 2984
rect 226058 2972 226064 2984
rect 223632 2944 226064 2972
rect 223632 2932 223638 2944
rect 226058 2932 226064 2944
rect 226116 2932 226122 2984
rect 226613 2975 226671 2981
rect 226613 2941 226625 2975
rect 226659 2972 226671 2975
rect 227622 2972 227628 2984
rect 226659 2944 227628 2972
rect 226659 2941 226671 2944
rect 226613 2935 226671 2941
rect 227622 2932 227628 2944
rect 227680 2932 227686 2984
rect 234586 2972 234614 3012
rect 242526 3000 242532 3012
rect 242584 3000 242590 3052
rect 257617 3043 257675 3049
rect 257617 3009 257629 3043
rect 257663 3040 257675 3043
rect 257982 3040 257988 3052
rect 257663 3012 257988 3040
rect 257663 3009 257675 3012
rect 257617 3003 257675 3009
rect 257982 3000 257988 3012
rect 258040 3000 258046 3052
rect 258994 3000 259000 3052
rect 259052 3000 259058 3052
rect 266173 3043 266231 3049
rect 266173 3009 266185 3043
rect 266219 3040 266231 3043
rect 266262 3040 266268 3052
rect 266219 3012 266268 3040
rect 266219 3009 266231 3012
rect 266173 3003 266231 3009
rect 266262 3000 266268 3012
rect 266320 3000 266326 3052
rect 266814 3000 266820 3052
rect 266872 3000 266878 3052
rect 267458 3000 267464 3052
rect 267516 3000 267522 3052
rect 268105 3043 268163 3049
rect 268105 3009 268117 3043
rect 268151 3040 268163 3043
rect 268654 3040 268660 3052
rect 268151 3012 268660 3040
rect 268151 3009 268163 3012
rect 268105 3003 268163 3009
rect 268654 3000 268660 3012
rect 268712 3000 268718 3052
rect 268749 3043 268807 3049
rect 268749 3009 268761 3043
rect 268795 3040 268807 3043
rect 269776 3040 269804 3080
rect 272058 3068 272064 3080
rect 272116 3068 272122 3120
rect 268795 3012 269804 3040
rect 268795 3009 268807 3012
rect 268749 3003 268807 3009
rect 269850 3000 269856 3052
rect 269908 3000 269914 3052
rect 270957 3043 271015 3049
rect 270957 3009 270969 3043
rect 271003 3040 271015 3043
rect 271874 3040 271880 3052
rect 271003 3012 271880 3040
rect 271003 3009 271015 3012
rect 270957 3003 271015 3009
rect 271874 3000 271880 3012
rect 271932 3000 271938 3052
rect 229756 2944 234614 2972
rect 214300 2876 216168 2904
rect 213273 2867 213331 2873
rect 209746 2808 210648 2836
rect 210712 2836 210740 2867
rect 210786 2836 210792 2848
rect 210712 2808 210792 2836
rect 209593 2799 209651 2805
rect 210786 2796 210792 2808
rect 210844 2836 210850 2848
rect 213288 2836 213316 2867
rect 215754 2836 215760 2848
rect 210844 2808 215760 2836
rect 210844 2796 210850 2808
rect 215754 2796 215760 2808
rect 215812 2796 215818 2848
rect 216140 2836 216168 2876
rect 217410 2864 217416 2916
rect 217468 2904 217474 2916
rect 229756 2904 229784 2944
rect 235810 2932 235816 2984
rect 235868 2932 235874 2984
rect 236086 2932 236092 2984
rect 236144 2972 236150 2984
rect 255314 2972 255320 2984
rect 236144 2944 255320 2972
rect 236144 2932 236150 2944
rect 255314 2932 255320 2944
rect 255372 2932 255378 2984
rect 262398 2932 262404 2984
rect 262456 2972 262462 2984
rect 262456 2944 267320 2972
rect 262456 2932 262462 2944
rect 217468 2876 229784 2904
rect 217468 2864 217474 2876
rect 229830 2864 229836 2916
rect 229888 2904 229894 2916
rect 246482 2904 246488 2916
rect 229888 2876 246488 2904
rect 229888 2864 229894 2876
rect 246482 2864 246488 2876
rect 246540 2864 246546 2916
rect 260101 2907 260159 2913
rect 260101 2873 260113 2907
rect 260147 2904 260159 2907
rect 267182 2904 267188 2916
rect 260147 2876 267188 2904
rect 260147 2873 260159 2876
rect 260101 2867 260159 2873
rect 267182 2864 267188 2876
rect 267240 2864 267246 2916
rect 267292 2913 267320 2944
rect 268286 2932 268292 2984
rect 268344 2972 268350 2984
rect 268344 2944 270816 2972
rect 268344 2932 268350 2944
rect 267277 2907 267335 2913
rect 267277 2873 267289 2907
rect 267323 2873 267335 2907
rect 267277 2867 267335 2873
rect 267921 2907 267979 2913
rect 267921 2873 267933 2907
rect 267967 2904 267979 2907
rect 269114 2904 269120 2916
rect 267967 2876 269120 2904
rect 267967 2873 267979 2876
rect 267921 2867 267979 2873
rect 269114 2864 269120 2876
rect 269172 2864 269178 2916
rect 270788 2913 270816 2944
rect 270773 2907 270831 2913
rect 270773 2873 270785 2907
rect 270819 2873 270831 2907
rect 270773 2867 270831 2873
rect 216582 2836 216588 2848
rect 216140 2808 216588 2836
rect 216582 2796 216588 2808
rect 216640 2796 216646 2848
rect 217778 2796 217784 2848
rect 217836 2836 217842 2848
rect 218149 2839 218207 2845
rect 218149 2836 218161 2839
rect 217836 2808 218161 2836
rect 217836 2796 217842 2808
rect 218149 2805 218161 2808
rect 218195 2805 218207 2839
rect 218149 2799 218207 2805
rect 219434 2796 219440 2848
rect 219492 2796 219498 2848
rect 223482 2796 223488 2848
rect 223540 2836 223546 2848
rect 226518 2836 226524 2848
rect 223540 2808 226524 2836
rect 223540 2796 223546 2808
rect 226518 2796 226524 2808
rect 226576 2796 226582 2848
rect 227254 2796 227260 2848
rect 227312 2796 227318 2848
rect 228266 2796 228272 2848
rect 228324 2796 228330 2848
rect 231670 2796 231676 2848
rect 231728 2836 231734 2848
rect 238662 2836 238668 2848
rect 231728 2808 238668 2836
rect 231728 2796 231734 2808
rect 238662 2796 238668 2808
rect 238720 2796 238726 2848
rect 257801 2839 257859 2845
rect 257801 2805 257813 2839
rect 257847 2836 257859 2839
rect 258074 2836 258080 2848
rect 257847 2808 258080 2836
rect 257847 2805 257859 2808
rect 257801 2799 257859 2805
rect 258074 2796 258080 2808
rect 258132 2796 258138 2848
rect 259178 2796 259184 2848
rect 259236 2796 259242 2848
rect 265526 2796 265532 2848
rect 265584 2796 265590 2848
rect 266630 2796 266636 2848
rect 266688 2796 266694 2848
rect 266814 2796 266820 2848
rect 266872 2836 266878 2848
rect 268470 2836 268476 2848
rect 266872 2808 268476 2836
rect 266872 2796 266878 2808
rect 268470 2796 268476 2808
rect 268528 2796 268534 2848
rect 270037 2839 270095 2845
rect 270037 2805 270049 2839
rect 270083 2836 270095 2839
rect 270494 2836 270500 2848
rect 270083 2808 270500 2836
rect 270083 2805 270095 2808
rect 270037 2799 270095 2805
rect 270494 2796 270500 2808
rect 270552 2796 270558 2848
rect 1104 2746 271492 2768
rect 1104 2694 34748 2746
rect 34800 2694 34812 2746
rect 34864 2694 34876 2746
rect 34928 2694 34940 2746
rect 34992 2694 35004 2746
rect 35056 2694 102345 2746
rect 102397 2694 102409 2746
rect 102461 2694 102473 2746
rect 102525 2694 102537 2746
rect 102589 2694 102601 2746
rect 102653 2694 169942 2746
rect 169994 2694 170006 2746
rect 170058 2694 170070 2746
rect 170122 2694 170134 2746
rect 170186 2694 170198 2746
rect 170250 2694 237539 2746
rect 237591 2694 237603 2746
rect 237655 2694 237667 2746
rect 237719 2694 237731 2746
rect 237783 2694 237795 2746
rect 237847 2694 271492 2746
rect 1104 2672 271492 2694
rect 23474 2592 23480 2644
rect 23532 2632 23538 2644
rect 23937 2635 23995 2641
rect 23937 2632 23949 2635
rect 23532 2604 23949 2632
rect 23532 2592 23538 2604
rect 23937 2601 23949 2604
rect 23983 2601 23995 2635
rect 23937 2595 23995 2601
rect 25225 2635 25283 2641
rect 25225 2601 25237 2635
rect 25271 2632 25283 2635
rect 25774 2632 25780 2644
rect 25271 2604 25780 2632
rect 25271 2601 25283 2604
rect 25225 2595 25283 2601
rect 25774 2592 25780 2604
rect 25832 2592 25838 2644
rect 26234 2592 26240 2644
rect 26292 2592 26298 2644
rect 26510 2592 26516 2644
rect 26568 2632 26574 2644
rect 27065 2635 27123 2641
rect 27065 2632 27077 2635
rect 26568 2604 27077 2632
rect 26568 2592 26574 2604
rect 27065 2601 27077 2604
rect 27111 2601 27123 2635
rect 27065 2595 27123 2601
rect 27982 2592 27988 2644
rect 28040 2632 28046 2644
rect 28077 2635 28135 2641
rect 28077 2632 28089 2635
rect 28040 2604 28089 2632
rect 28040 2592 28046 2604
rect 28077 2601 28089 2604
rect 28123 2601 28135 2635
rect 28077 2595 28135 2601
rect 58621 2635 58679 2641
rect 58621 2601 58633 2635
rect 58667 2632 58679 2635
rect 58894 2632 58900 2644
rect 58667 2604 58900 2632
rect 58667 2601 58679 2604
rect 58621 2595 58679 2601
rect 58894 2592 58900 2604
rect 58952 2592 58958 2644
rect 60734 2592 60740 2644
rect 60792 2632 60798 2644
rect 60829 2635 60887 2641
rect 60829 2632 60841 2635
rect 60792 2604 60841 2632
rect 60792 2592 60798 2604
rect 60829 2601 60841 2604
rect 60875 2601 60887 2635
rect 60829 2595 60887 2601
rect 85390 2592 85396 2644
rect 85448 2632 85454 2644
rect 85761 2635 85819 2641
rect 85761 2632 85773 2635
rect 85448 2604 85773 2632
rect 85448 2592 85454 2604
rect 85761 2601 85773 2604
rect 85807 2632 85819 2635
rect 85807 2604 98316 2632
rect 85807 2601 85819 2604
rect 85761 2595 85819 2601
rect 4798 2524 4804 2576
rect 4856 2564 4862 2576
rect 23566 2564 23572 2576
rect 4856 2536 23572 2564
rect 4856 2524 4862 2536
rect 23566 2524 23572 2536
rect 23624 2524 23630 2576
rect 25130 2524 25136 2576
rect 25188 2564 25194 2576
rect 33134 2564 33140 2576
rect 25188 2536 33140 2564
rect 25188 2524 25194 2536
rect 33134 2524 33140 2536
rect 33192 2524 33198 2576
rect 70854 2524 70860 2576
rect 70912 2564 70918 2576
rect 96890 2564 96896 2576
rect 70912 2536 96660 2564
rect 70912 2524 70918 2536
rect 1857 2499 1915 2505
rect 1857 2465 1869 2499
rect 1903 2496 1915 2499
rect 36630 2496 36636 2508
rect 1903 2468 36636 2496
rect 1903 2465 1915 2468
rect 1857 2459 1915 2465
rect 36630 2456 36636 2468
rect 36688 2456 36694 2508
rect 37182 2456 37188 2508
rect 37240 2456 37246 2508
rect 53742 2456 53748 2508
rect 53800 2456 53806 2508
rect 53852 2468 78168 2496
rect 1578 2388 1584 2440
rect 1636 2388 1642 2440
rect 23750 2388 23756 2440
rect 23808 2388 23814 2440
rect 24946 2388 24952 2440
rect 25004 2388 25010 2440
rect 25038 2388 25044 2440
rect 25096 2388 25102 2440
rect 25498 2388 25504 2440
rect 25556 2388 25562 2440
rect 25593 2431 25651 2437
rect 25593 2397 25605 2431
rect 25639 2428 25651 2431
rect 25682 2428 25688 2440
rect 25639 2400 25688 2428
rect 25639 2397 25651 2400
rect 25593 2391 25651 2397
rect 25682 2388 25688 2400
rect 25740 2388 25746 2440
rect 25869 2431 25927 2437
rect 25869 2397 25881 2431
rect 25915 2397 25927 2431
rect 25869 2391 25927 2397
rect 26053 2431 26111 2437
rect 26053 2397 26065 2431
rect 26099 2428 26111 2431
rect 26142 2428 26148 2440
rect 26099 2400 26148 2428
rect 26099 2397 26111 2400
rect 26053 2391 26111 2397
rect 2590 2320 2596 2372
rect 2648 2360 2654 2372
rect 24765 2363 24823 2369
rect 2648 2332 22094 2360
rect 2648 2320 2654 2332
rect 22066 2292 22094 2332
rect 24765 2329 24777 2363
rect 24811 2360 24823 2363
rect 25516 2360 25544 2388
rect 25884 2360 25912 2391
rect 26142 2388 26148 2400
rect 26200 2388 26206 2440
rect 26786 2388 26792 2440
rect 26844 2388 26850 2440
rect 26881 2431 26939 2437
rect 26881 2397 26893 2431
rect 26927 2397 26939 2431
rect 26881 2391 26939 2397
rect 24811 2332 25912 2360
rect 26160 2360 26188 2388
rect 26896 2360 26924 2391
rect 27338 2388 27344 2440
rect 27396 2428 27402 2440
rect 27433 2431 27491 2437
rect 27433 2428 27445 2431
rect 27396 2400 27445 2428
rect 27396 2388 27402 2400
rect 27433 2397 27445 2400
rect 27479 2428 27491 2431
rect 27801 2431 27859 2437
rect 27801 2428 27813 2431
rect 27479 2400 27813 2428
rect 27479 2397 27491 2400
rect 27433 2391 27491 2397
rect 27801 2397 27813 2400
rect 27847 2397 27859 2431
rect 27801 2391 27859 2397
rect 27816 2360 27844 2391
rect 27890 2388 27896 2440
rect 27948 2388 27954 2440
rect 28534 2388 28540 2440
rect 28592 2388 28598 2440
rect 31938 2388 31944 2440
rect 31996 2428 32002 2440
rect 32217 2431 32275 2437
rect 32217 2428 32229 2431
rect 31996 2400 32229 2428
rect 31996 2388 32002 2400
rect 32217 2397 32229 2400
rect 32263 2397 32275 2431
rect 32217 2391 32275 2397
rect 32401 2431 32459 2437
rect 32401 2397 32413 2431
rect 32447 2428 32459 2431
rect 32490 2428 32496 2440
rect 32447 2400 32496 2428
rect 32447 2397 32459 2400
rect 32401 2391 32459 2397
rect 32490 2388 32496 2400
rect 32548 2428 32554 2440
rect 38654 2428 38660 2440
rect 32548 2400 38660 2428
rect 32548 2388 32554 2400
rect 38654 2388 38660 2400
rect 38712 2388 38718 2440
rect 53466 2388 53472 2440
rect 53524 2428 53530 2440
rect 53852 2428 53880 2468
rect 53524 2400 53880 2428
rect 53929 2431 53987 2437
rect 53524 2388 53530 2400
rect 53929 2397 53941 2431
rect 53975 2428 53987 2431
rect 54018 2428 54024 2440
rect 53975 2400 54024 2428
rect 53975 2397 53987 2400
rect 53929 2391 53987 2397
rect 54018 2388 54024 2400
rect 54076 2388 54082 2440
rect 54202 2388 54208 2440
rect 54260 2428 54266 2440
rect 54665 2431 54723 2437
rect 54665 2428 54677 2431
rect 54260 2400 54677 2428
rect 54260 2388 54266 2400
rect 54665 2397 54677 2400
rect 54711 2397 54723 2431
rect 54665 2391 54723 2397
rect 55030 2388 55036 2440
rect 55088 2428 55094 2440
rect 55493 2431 55551 2437
rect 55493 2428 55505 2431
rect 55088 2400 55505 2428
rect 55088 2388 55094 2400
rect 55493 2397 55505 2400
rect 55539 2397 55551 2431
rect 55493 2391 55551 2397
rect 57514 2388 57520 2440
rect 57572 2428 57578 2440
rect 57609 2431 57667 2437
rect 57609 2428 57621 2431
rect 57572 2400 57621 2428
rect 57572 2388 57578 2400
rect 57609 2397 57621 2400
rect 57655 2397 57667 2431
rect 57609 2391 57667 2397
rect 59173 2431 59231 2437
rect 59173 2397 59185 2431
rect 59219 2428 59231 2431
rect 59262 2428 59268 2440
rect 59219 2400 59268 2428
rect 59219 2397 59231 2400
rect 59173 2391 59231 2397
rect 59262 2388 59268 2400
rect 59320 2388 59326 2440
rect 59998 2388 60004 2440
rect 60056 2428 60062 2440
rect 60645 2431 60703 2437
rect 60645 2428 60657 2431
rect 60056 2400 60657 2428
rect 60056 2388 60062 2400
rect 60645 2397 60657 2400
rect 60691 2397 60703 2431
rect 60645 2391 60703 2397
rect 62666 2388 62672 2440
rect 62724 2428 62730 2440
rect 62761 2431 62819 2437
rect 62761 2428 62773 2431
rect 62724 2400 62773 2428
rect 62724 2388 62730 2400
rect 62761 2397 62773 2400
rect 62807 2397 62819 2431
rect 62761 2391 62819 2397
rect 65242 2388 65248 2440
rect 65300 2428 65306 2440
rect 65797 2431 65855 2437
rect 65797 2428 65809 2431
rect 65300 2400 65809 2428
rect 65300 2388 65306 2400
rect 65797 2397 65809 2400
rect 65843 2397 65855 2431
rect 65797 2391 65855 2397
rect 71314 2388 71320 2440
rect 71372 2388 71378 2440
rect 71593 2431 71651 2437
rect 71593 2397 71605 2431
rect 71639 2428 71651 2431
rect 73154 2428 73160 2440
rect 71639 2400 73160 2428
rect 71639 2397 71651 2400
rect 71593 2391 71651 2397
rect 73154 2388 73160 2400
rect 73212 2388 73218 2440
rect 73522 2388 73528 2440
rect 73580 2388 73586 2440
rect 73798 2388 73804 2440
rect 73856 2388 73862 2440
rect 76466 2388 76472 2440
rect 76524 2388 76530 2440
rect 76742 2388 76748 2440
rect 76800 2388 76806 2440
rect 77938 2388 77944 2440
rect 77996 2388 78002 2440
rect 78140 2428 78168 2468
rect 78214 2456 78220 2508
rect 78272 2456 78278 2508
rect 87966 2496 87972 2508
rect 78324 2468 85344 2496
rect 78324 2428 78352 2468
rect 78140 2400 78352 2428
rect 79410 2388 79416 2440
rect 79468 2388 79474 2440
rect 79689 2431 79747 2437
rect 79689 2397 79701 2431
rect 79735 2428 79747 2431
rect 79962 2428 79968 2440
rect 79735 2400 79968 2428
rect 79735 2397 79747 2400
rect 79689 2391 79747 2397
rect 79962 2388 79968 2400
rect 80020 2388 80026 2440
rect 82081 2431 82139 2437
rect 82081 2397 82093 2431
rect 82127 2397 82139 2431
rect 82081 2391 82139 2397
rect 35618 2360 35624 2372
rect 26160 2332 27752 2360
rect 27816 2332 35624 2360
rect 24811 2329 24823 2332
rect 24765 2323 24823 2329
rect 27246 2292 27252 2304
rect 22066 2264 27252 2292
rect 27246 2252 27252 2264
rect 27304 2252 27310 2304
rect 27724 2292 27752 2332
rect 35618 2320 35624 2332
rect 35676 2320 35682 2372
rect 36446 2320 36452 2372
rect 36504 2360 36510 2372
rect 36504 2332 37044 2360
rect 36504 2320 36510 2332
rect 27890 2292 27896 2304
rect 27724 2264 27896 2292
rect 27890 2252 27896 2264
rect 27948 2252 27954 2304
rect 28718 2252 28724 2304
rect 28776 2252 28782 2304
rect 32306 2252 32312 2304
rect 32364 2292 32370 2304
rect 32585 2295 32643 2301
rect 32585 2292 32597 2295
rect 32364 2264 32597 2292
rect 32364 2252 32370 2264
rect 32585 2261 32597 2264
rect 32631 2261 32643 2295
rect 32585 2255 32643 2261
rect 33042 2252 33048 2304
rect 33100 2252 33106 2304
rect 36722 2252 36728 2304
rect 36780 2292 36786 2304
rect 36909 2295 36967 2301
rect 36909 2292 36921 2295
rect 36780 2264 36921 2292
rect 36780 2252 36786 2264
rect 36909 2261 36921 2264
rect 36955 2261 36967 2295
rect 37016 2292 37044 2332
rect 37090 2320 37096 2372
rect 37148 2360 37154 2372
rect 37185 2363 37243 2369
rect 37185 2360 37197 2363
rect 37148 2332 37197 2360
rect 37148 2320 37154 2332
rect 37185 2329 37197 2332
rect 37231 2329 37243 2363
rect 37185 2323 37243 2329
rect 37274 2320 37280 2372
rect 37332 2320 37338 2372
rect 37645 2363 37703 2369
rect 37645 2329 37657 2363
rect 37691 2329 37703 2363
rect 37645 2323 37703 2329
rect 37660 2292 37688 2323
rect 40034 2320 40040 2372
rect 40092 2360 40098 2372
rect 82096 2360 82124 2391
rect 82354 2388 82360 2440
rect 82412 2388 82418 2440
rect 83553 2431 83611 2437
rect 83553 2428 83565 2431
rect 83108 2400 83565 2428
rect 82998 2360 83004 2372
rect 40092 2332 74534 2360
rect 82096 2332 83004 2360
rect 40092 2320 40098 2332
rect 37016 2264 37688 2292
rect 36909 2255 36967 2261
rect 37734 2252 37740 2304
rect 37792 2292 37798 2304
rect 38013 2295 38071 2301
rect 38013 2292 38025 2295
rect 37792 2264 38025 2292
rect 37792 2252 37798 2264
rect 38013 2261 38025 2264
rect 38059 2261 38071 2295
rect 38013 2255 38071 2261
rect 38194 2252 38200 2304
rect 38252 2252 38258 2304
rect 53834 2252 53840 2304
rect 53892 2292 53898 2304
rect 54113 2295 54171 2301
rect 54113 2292 54125 2295
rect 53892 2264 54125 2292
rect 53892 2252 53898 2264
rect 54113 2261 54125 2264
rect 54159 2261 54171 2295
rect 54113 2255 54171 2261
rect 54846 2252 54852 2304
rect 54904 2252 54910 2304
rect 55674 2252 55680 2304
rect 55732 2252 55738 2304
rect 57790 2252 57796 2304
rect 57848 2252 57854 2304
rect 59354 2252 59360 2304
rect 59412 2252 59418 2304
rect 62942 2252 62948 2304
rect 63000 2252 63006 2304
rect 65610 2252 65616 2304
rect 65668 2292 65674 2304
rect 65981 2295 66039 2301
rect 65981 2292 65993 2295
rect 65668 2264 65993 2292
rect 65668 2252 65674 2264
rect 65981 2261 65993 2264
rect 66027 2261 66039 2295
rect 65981 2255 66039 2261
rect 66622 2252 66628 2304
rect 66680 2252 66686 2304
rect 74506 2292 74534 2332
rect 82998 2320 83004 2332
rect 83056 2320 83062 2372
rect 83108 2292 83136 2400
rect 83553 2397 83565 2400
rect 83599 2397 83611 2431
rect 85316 2428 85344 2468
rect 85500 2468 87972 2496
rect 85500 2428 85528 2468
rect 87966 2456 87972 2468
rect 88024 2456 88030 2508
rect 88061 2499 88119 2505
rect 88061 2465 88073 2499
rect 88107 2496 88119 2499
rect 90177 2499 90235 2505
rect 90177 2496 90189 2499
rect 88107 2468 90189 2496
rect 88107 2465 88119 2468
rect 88061 2459 88119 2465
rect 90177 2465 90189 2468
rect 90223 2496 90235 2499
rect 90545 2499 90603 2505
rect 90545 2496 90557 2499
rect 90223 2468 90557 2496
rect 90223 2465 90235 2468
rect 90177 2459 90235 2465
rect 90545 2465 90557 2468
rect 90591 2496 90603 2499
rect 96338 2496 96344 2508
rect 90591 2468 96344 2496
rect 90591 2465 90603 2468
rect 90545 2459 90603 2465
rect 96338 2456 96344 2468
rect 96396 2456 96402 2508
rect 85316 2400 85528 2428
rect 87417 2431 87475 2437
rect 83553 2391 83611 2397
rect 87417 2397 87429 2431
rect 87463 2397 87475 2431
rect 87417 2391 87475 2397
rect 83734 2320 83740 2372
rect 83792 2360 83798 2372
rect 84010 2360 84016 2372
rect 83792 2332 84016 2360
rect 83792 2320 83798 2332
rect 84010 2320 84016 2332
rect 84068 2320 84074 2372
rect 85390 2360 85396 2372
rect 84166 2332 85396 2360
rect 74506 2264 83136 2292
rect 83277 2295 83335 2301
rect 83277 2261 83289 2295
rect 83323 2292 83335 2295
rect 84166 2292 84194 2332
rect 85390 2320 85396 2332
rect 85448 2320 85454 2372
rect 87432 2360 87460 2391
rect 88334 2388 88340 2440
rect 88392 2388 88398 2440
rect 89898 2388 89904 2440
rect 89956 2428 89962 2440
rect 90637 2431 90695 2437
rect 90637 2428 90649 2431
rect 89956 2400 90649 2428
rect 89956 2388 89962 2400
rect 90637 2397 90649 2400
rect 90683 2397 90695 2431
rect 90637 2391 90695 2397
rect 91094 2388 91100 2440
rect 91152 2428 91158 2440
rect 91557 2431 91615 2437
rect 91557 2428 91569 2431
rect 91152 2400 91569 2428
rect 91152 2388 91158 2400
rect 91557 2397 91569 2400
rect 91603 2397 91615 2431
rect 91557 2391 91615 2397
rect 92750 2388 92756 2440
rect 92808 2428 92814 2440
rect 92845 2431 92903 2437
rect 92845 2428 92857 2431
rect 92808 2400 92857 2428
rect 92808 2388 92814 2400
rect 92845 2397 92857 2400
rect 92891 2397 92903 2431
rect 92845 2391 92903 2397
rect 93670 2388 93676 2440
rect 93728 2388 93734 2440
rect 94406 2388 94412 2440
rect 94464 2388 94470 2440
rect 95145 2431 95203 2437
rect 95145 2397 95157 2431
rect 95191 2428 95203 2431
rect 95418 2428 95424 2440
rect 95191 2400 95424 2428
rect 95191 2397 95203 2400
rect 95145 2391 95203 2397
rect 95418 2388 95424 2400
rect 95476 2388 95482 2440
rect 95881 2431 95939 2437
rect 95881 2397 95893 2431
rect 95927 2428 95939 2431
rect 96246 2428 96252 2440
rect 95927 2400 96252 2428
rect 95927 2397 95939 2400
rect 95881 2391 95939 2397
rect 96246 2388 96252 2400
rect 96304 2388 96310 2440
rect 96632 2428 96660 2536
rect 96724 2536 96896 2564
rect 96724 2505 96752 2536
rect 96890 2524 96896 2536
rect 96948 2524 96954 2576
rect 97350 2524 97356 2576
rect 97408 2524 97414 2576
rect 96709 2499 96767 2505
rect 96709 2465 96721 2499
rect 96755 2465 96767 2499
rect 96709 2459 96767 2465
rect 97442 2456 97448 2508
rect 97500 2496 97506 2508
rect 97746 2499 97804 2505
rect 97746 2496 97758 2499
rect 97500 2468 97758 2496
rect 97500 2456 97506 2468
rect 97746 2465 97758 2468
rect 97792 2465 97804 2499
rect 97746 2459 97804 2465
rect 96893 2431 96951 2437
rect 96893 2428 96905 2431
rect 96632 2400 96905 2428
rect 96893 2397 96905 2400
rect 96939 2397 96951 2431
rect 96893 2391 96951 2397
rect 97626 2388 97632 2440
rect 97684 2388 97690 2440
rect 97902 2422 97908 2474
rect 97960 2422 97966 2474
rect 98086 2456 98092 2508
rect 98144 2496 98150 2508
rect 98288 2496 98316 2604
rect 98546 2592 98552 2644
rect 98604 2592 98610 2644
rect 98822 2592 98828 2644
rect 98880 2632 98886 2644
rect 98880 2604 105216 2632
rect 98880 2592 98886 2604
rect 98638 2524 98644 2576
rect 98696 2564 98702 2576
rect 103330 2564 103336 2576
rect 98696 2536 103336 2564
rect 98696 2524 98702 2536
rect 103330 2524 103336 2536
rect 103388 2524 103394 2576
rect 104069 2567 104127 2573
rect 104069 2533 104081 2567
rect 104115 2564 104127 2567
rect 104158 2564 104164 2576
rect 104115 2536 104164 2564
rect 104115 2533 104127 2536
rect 104069 2527 104127 2533
rect 104158 2524 104164 2536
rect 104216 2524 104222 2576
rect 105188 2564 105216 2604
rect 105262 2592 105268 2644
rect 105320 2592 105326 2644
rect 107654 2632 107660 2644
rect 106246 2604 107660 2632
rect 106246 2564 106274 2604
rect 107654 2592 107660 2604
rect 107712 2632 107718 2644
rect 149146 2632 149152 2644
rect 107712 2604 149152 2632
rect 107712 2592 107718 2604
rect 149146 2592 149152 2604
rect 149204 2592 149210 2644
rect 156874 2632 156880 2644
rect 154546 2604 156880 2632
rect 143718 2564 143724 2576
rect 105188 2536 106274 2564
rect 142080 2536 143724 2564
rect 98144 2468 98316 2496
rect 98144 2456 98150 2468
rect 98454 2456 98460 2508
rect 98512 2496 98518 2508
rect 99377 2499 99435 2505
rect 99377 2496 99389 2499
rect 98512 2468 99389 2496
rect 98512 2456 98518 2468
rect 99377 2465 99389 2468
rect 99423 2465 99435 2499
rect 99377 2459 99435 2465
rect 99561 2499 99619 2505
rect 99561 2465 99573 2499
rect 99607 2496 99619 2499
rect 99742 2496 99748 2508
rect 99607 2468 99748 2496
rect 99607 2465 99619 2468
rect 99561 2459 99619 2465
rect 99742 2456 99748 2468
rect 99800 2456 99806 2508
rect 103422 2456 103428 2508
rect 103480 2456 103486 2508
rect 104342 2456 104348 2508
rect 104400 2456 104406 2508
rect 104483 2499 104541 2505
rect 104483 2465 104495 2499
rect 104529 2496 104541 2499
rect 107470 2496 107476 2508
rect 104529 2468 107476 2496
rect 104529 2465 104541 2468
rect 104483 2459 104541 2465
rect 107470 2456 107476 2468
rect 107528 2456 107534 2508
rect 107930 2456 107936 2508
rect 107988 2496 107994 2508
rect 108485 2499 108543 2505
rect 108485 2496 108497 2499
rect 107988 2468 108497 2496
rect 107988 2456 107994 2468
rect 108485 2465 108497 2468
rect 108531 2465 108543 2499
rect 108485 2459 108543 2465
rect 109034 2456 109040 2508
rect 109092 2456 109098 2508
rect 139118 2456 139124 2508
rect 139176 2456 139182 2508
rect 141142 2456 141148 2508
rect 141200 2496 141206 2508
rect 142080 2496 142108 2536
rect 143718 2524 143724 2536
rect 143776 2524 143782 2576
rect 144917 2567 144975 2573
rect 144917 2533 144929 2567
rect 144963 2564 144975 2567
rect 145650 2564 145656 2576
rect 144963 2536 145656 2564
rect 144963 2533 144975 2536
rect 144917 2527 144975 2533
rect 145650 2524 145656 2536
rect 145708 2524 145714 2576
rect 148870 2524 148876 2576
rect 148928 2524 148934 2576
rect 150636 2536 153332 2564
rect 141200 2468 142108 2496
rect 143077 2499 143135 2505
rect 141200 2456 141206 2468
rect 143077 2465 143089 2499
rect 143123 2496 143135 2499
rect 143166 2496 143172 2508
rect 143123 2468 143172 2496
rect 143123 2465 143135 2468
rect 143077 2459 143135 2465
rect 143166 2456 143172 2468
rect 143224 2456 143230 2508
rect 143997 2499 144055 2505
rect 143997 2465 144009 2499
rect 144043 2496 144055 2499
rect 144454 2496 144460 2508
rect 144043 2468 144460 2496
rect 144043 2465 144055 2468
rect 143997 2459 144055 2465
rect 144454 2456 144460 2468
rect 144512 2456 144518 2508
rect 146202 2456 146208 2508
rect 146260 2496 146266 2508
rect 148229 2499 148287 2505
rect 148229 2496 148241 2499
rect 146260 2468 148241 2496
rect 146260 2456 146266 2468
rect 148229 2465 148241 2468
rect 148275 2465 148287 2499
rect 148229 2459 148287 2465
rect 149146 2456 149152 2508
rect 149204 2456 149210 2508
rect 149287 2499 149345 2505
rect 149287 2465 149299 2499
rect 149333 2496 149345 2499
rect 150636 2496 150664 2536
rect 149333 2468 150664 2496
rect 150713 2499 150771 2505
rect 149333 2465 149345 2468
rect 149287 2459 149345 2465
rect 150713 2465 150725 2499
rect 150759 2496 150771 2499
rect 150986 2496 150992 2508
rect 150759 2468 150992 2496
rect 150759 2465 150771 2468
rect 150713 2459 150771 2465
rect 150986 2456 150992 2468
rect 151044 2456 151050 2508
rect 152366 2456 152372 2508
rect 152424 2456 152430 2508
rect 153304 2496 153332 2536
rect 154546 2496 154574 2604
rect 156874 2592 156880 2604
rect 156932 2592 156938 2644
rect 156966 2592 156972 2644
rect 157024 2632 157030 2644
rect 157150 2632 157156 2644
rect 157024 2604 157156 2632
rect 157024 2592 157030 2604
rect 157150 2592 157156 2604
rect 157208 2592 157214 2644
rect 157334 2592 157340 2644
rect 157392 2632 157398 2644
rect 157889 2635 157947 2641
rect 157889 2632 157901 2635
rect 157392 2604 157901 2632
rect 157392 2592 157398 2604
rect 157889 2601 157901 2604
rect 157935 2601 157947 2635
rect 157889 2595 157947 2601
rect 160094 2592 160100 2644
rect 160152 2632 160158 2644
rect 160557 2635 160615 2641
rect 160557 2632 160569 2635
rect 160152 2604 160569 2632
rect 160152 2592 160158 2604
rect 160557 2601 160569 2604
rect 160603 2601 160615 2635
rect 160557 2595 160615 2601
rect 160738 2592 160744 2644
rect 160796 2632 160802 2644
rect 161293 2635 161351 2641
rect 161293 2632 161305 2635
rect 160796 2604 161305 2632
rect 160796 2592 160802 2604
rect 161293 2601 161305 2604
rect 161339 2632 161351 2635
rect 161382 2632 161388 2644
rect 161339 2604 161388 2632
rect 161339 2601 161351 2604
rect 161293 2595 161351 2601
rect 161382 2592 161388 2604
rect 161440 2592 161446 2644
rect 176654 2592 176660 2644
rect 176712 2632 176718 2644
rect 176712 2604 187280 2632
rect 176712 2592 176718 2604
rect 155037 2567 155095 2573
rect 155037 2533 155049 2567
rect 155083 2564 155095 2567
rect 155126 2564 155132 2576
rect 155083 2536 155132 2564
rect 155083 2533 155095 2536
rect 155037 2527 155095 2533
rect 155126 2524 155132 2536
rect 155184 2524 155190 2576
rect 159450 2524 159456 2576
rect 159508 2564 159514 2576
rect 159508 2536 187096 2564
rect 159508 2524 159514 2536
rect 153304 2468 154574 2496
rect 156874 2456 156880 2508
rect 156932 2496 156938 2508
rect 179877 2499 179935 2505
rect 179877 2496 179889 2499
rect 156932 2468 179889 2496
rect 156932 2456 156938 2468
rect 179877 2465 179889 2468
rect 179923 2465 179935 2499
rect 179877 2459 179935 2465
rect 103609 2431 103667 2437
rect 103609 2428 103621 2431
rect 97905 2397 97917 2422
rect 97951 2397 97963 2422
rect 97905 2391 97963 2397
rect 101140 2400 103621 2428
rect 88521 2363 88579 2369
rect 87432 2332 88472 2360
rect 83323 2264 84194 2292
rect 83323 2261 83335 2264
rect 83277 2255 83335 2261
rect 87598 2252 87604 2304
rect 87656 2252 87662 2304
rect 88444 2292 88472 2332
rect 88521 2329 88533 2363
rect 88567 2360 88579 2363
rect 89530 2360 89536 2372
rect 88567 2332 89536 2360
rect 88567 2329 88579 2332
rect 88521 2323 88579 2329
rect 89530 2320 89536 2332
rect 89588 2360 89594 2372
rect 89588 2332 89714 2360
rect 89588 2320 89594 2332
rect 89254 2292 89260 2304
rect 88444 2264 89260 2292
rect 89254 2252 89260 2264
rect 89312 2252 89318 2304
rect 89686 2292 89714 2332
rect 91002 2320 91008 2372
rect 91060 2360 91066 2372
rect 91060 2332 96200 2360
rect 91060 2320 91066 2332
rect 90266 2292 90272 2304
rect 89686 2264 90272 2292
rect 90266 2252 90272 2264
rect 90324 2252 90330 2304
rect 90818 2252 90824 2304
rect 90876 2252 90882 2304
rect 91738 2252 91744 2304
rect 91796 2252 91802 2304
rect 93026 2252 93032 2304
rect 93084 2252 93090 2304
rect 93854 2252 93860 2304
rect 93912 2252 93918 2304
rect 94590 2252 94596 2304
rect 94648 2252 94654 2304
rect 95326 2252 95332 2304
rect 95384 2252 95390 2304
rect 96062 2252 96068 2304
rect 96120 2252 96126 2304
rect 96172 2292 96200 2332
rect 98380 2332 99144 2360
rect 98380 2292 98408 2332
rect 96172 2264 98408 2292
rect 99006 2252 99012 2304
rect 99064 2252 99070 2304
rect 99116 2292 99144 2332
rect 99190 2320 99196 2372
rect 99248 2360 99254 2372
rect 101140 2360 101168 2400
rect 103609 2397 103621 2400
rect 103655 2397 103667 2431
rect 103609 2391 103667 2397
rect 104618 2388 104624 2440
rect 104676 2388 104682 2440
rect 122006 2388 122012 2440
rect 122064 2428 122070 2440
rect 122469 2431 122527 2437
rect 122469 2428 122481 2431
rect 122064 2400 122481 2428
rect 122064 2388 122070 2400
rect 122469 2397 122481 2400
rect 122515 2397 122527 2431
rect 122469 2391 122527 2397
rect 124490 2388 124496 2440
rect 124548 2428 124554 2440
rect 124585 2431 124643 2437
rect 124585 2428 124597 2431
rect 124548 2400 124597 2428
rect 124548 2388 124554 2400
rect 124585 2397 124597 2400
rect 124631 2397 124643 2431
rect 124585 2391 124643 2397
rect 126149 2431 126207 2437
rect 126149 2397 126161 2431
rect 126195 2428 126207 2431
rect 126238 2428 126244 2440
rect 126195 2400 126244 2428
rect 126195 2397 126207 2400
rect 126149 2391 126207 2397
rect 126238 2388 126244 2400
rect 126296 2388 126302 2440
rect 127621 2431 127679 2437
rect 127621 2397 127633 2431
rect 127667 2428 127679 2431
rect 127894 2428 127900 2440
rect 127667 2400 127900 2428
rect 127667 2397 127679 2400
rect 127621 2391 127679 2397
rect 127894 2388 127900 2400
rect 127952 2388 127958 2440
rect 128357 2431 128415 2437
rect 128357 2397 128369 2431
rect 128403 2428 128415 2431
rect 128630 2428 128636 2440
rect 128403 2400 128636 2428
rect 128403 2397 128415 2400
rect 128357 2391 128415 2397
rect 128630 2388 128636 2400
rect 128688 2388 128694 2440
rect 129642 2388 129648 2440
rect 129700 2428 129706 2440
rect 129829 2431 129887 2437
rect 129829 2428 129841 2431
rect 129700 2400 129841 2428
rect 129700 2388 129706 2400
rect 129829 2397 129841 2400
rect 129875 2397 129887 2431
rect 129829 2391 129887 2397
rect 131393 2431 131451 2437
rect 131393 2397 131405 2431
rect 131439 2428 131451 2431
rect 131666 2428 131672 2440
rect 131439 2400 131672 2428
rect 131439 2397 131451 2400
rect 131393 2391 131451 2397
rect 131666 2388 131672 2400
rect 131724 2388 131730 2440
rect 132773 2431 132831 2437
rect 132773 2397 132785 2431
rect 132819 2428 132831 2431
rect 133322 2428 133328 2440
rect 132819 2400 133328 2428
rect 132819 2397 132831 2400
rect 132773 2391 132831 2397
rect 133322 2388 133328 2400
rect 133380 2388 133386 2440
rect 133509 2431 133567 2437
rect 133509 2397 133521 2431
rect 133555 2428 133567 2431
rect 133598 2428 133604 2440
rect 133555 2400 133604 2428
rect 133555 2397 133567 2400
rect 133509 2391 133567 2397
rect 133598 2388 133604 2400
rect 133656 2388 133662 2440
rect 134245 2431 134303 2437
rect 134245 2397 134257 2431
rect 134291 2428 134303 2431
rect 134334 2428 134340 2440
rect 134291 2400 134340 2428
rect 134291 2397 134303 2400
rect 134245 2391 134303 2397
rect 134334 2388 134340 2400
rect 134392 2388 134398 2440
rect 138937 2431 138995 2437
rect 138937 2397 138949 2431
rect 138983 2397 138995 2431
rect 138937 2391 138995 2397
rect 99248 2332 101168 2360
rect 99248 2320 99254 2332
rect 101214 2320 101220 2372
rect 101272 2320 101278 2372
rect 107286 2320 107292 2372
rect 107344 2360 107350 2372
rect 108669 2363 108727 2369
rect 108669 2360 108681 2363
rect 107344 2332 108681 2360
rect 107344 2320 107350 2332
rect 108669 2329 108681 2332
rect 108715 2360 108727 2363
rect 109310 2360 109316 2372
rect 108715 2332 109316 2360
rect 108715 2329 108727 2332
rect 108669 2323 108727 2329
rect 109310 2320 109316 2332
rect 109368 2320 109374 2372
rect 133230 2320 133236 2372
rect 133288 2360 133294 2372
rect 138952 2360 138980 2391
rect 142798 2388 142804 2440
rect 142856 2428 142862 2440
rect 144178 2437 144184 2440
rect 143261 2431 143319 2437
rect 143261 2428 143273 2431
rect 142856 2400 143273 2428
rect 142856 2388 142862 2400
rect 143261 2397 143273 2400
rect 143307 2397 143319 2431
rect 143261 2391 143319 2397
rect 144135 2431 144184 2437
rect 144135 2397 144147 2431
rect 144181 2397 144184 2431
rect 144135 2391 144184 2397
rect 144178 2388 144184 2391
rect 144236 2388 144242 2440
rect 144270 2388 144276 2440
rect 144328 2388 144334 2440
rect 147766 2388 147772 2440
rect 147824 2428 147830 2440
rect 148413 2431 148471 2437
rect 148413 2428 148425 2431
rect 147824 2400 148425 2428
rect 147824 2388 147830 2400
rect 148413 2397 148425 2400
rect 148459 2397 148471 2431
rect 148413 2391 148471 2397
rect 149422 2388 149428 2440
rect 149480 2388 149486 2440
rect 150069 2431 150127 2437
rect 150069 2397 150081 2431
rect 150115 2428 150127 2431
rect 150529 2431 150587 2437
rect 150529 2428 150541 2431
rect 150115 2400 150541 2428
rect 150115 2397 150127 2400
rect 150069 2391 150127 2397
rect 150529 2397 150541 2400
rect 150575 2397 150587 2431
rect 150529 2391 150587 2397
rect 155218 2388 155224 2440
rect 155276 2388 155282 2440
rect 156598 2437 156604 2440
rect 156555 2431 156604 2437
rect 156555 2430 156567 2431
rect 156524 2400 156567 2430
rect 156555 2397 156567 2400
rect 156601 2397 156604 2431
rect 156555 2391 156604 2397
rect 156598 2388 156604 2391
rect 156656 2388 156662 2440
rect 157334 2388 157340 2440
rect 157392 2388 157398 2440
rect 157702 2388 157708 2440
rect 157760 2388 157766 2440
rect 157794 2388 157800 2440
rect 157852 2428 157858 2440
rect 157852 2400 158576 2428
rect 157852 2388 157858 2400
rect 158548 2372 158576 2400
rect 158622 2388 158628 2440
rect 158680 2388 158686 2440
rect 159910 2388 159916 2440
rect 159968 2388 159974 2440
rect 160002 2388 160008 2440
rect 160060 2428 160066 2440
rect 160097 2431 160155 2437
rect 160097 2428 160109 2431
rect 160060 2400 160109 2428
rect 160060 2388 160066 2400
rect 160097 2397 160109 2400
rect 160143 2397 160155 2431
rect 160097 2391 160155 2397
rect 160370 2388 160376 2440
rect 160428 2388 160434 2440
rect 160741 2431 160799 2437
rect 160741 2397 160753 2431
rect 160787 2397 160799 2431
rect 160741 2391 160799 2397
rect 161569 2431 161627 2437
rect 161569 2397 161581 2431
rect 161615 2428 161627 2431
rect 162302 2428 162308 2440
rect 161615 2400 162308 2428
rect 161615 2397 161627 2400
rect 161569 2391 161627 2397
rect 139946 2360 139952 2372
rect 133288 2332 138014 2360
rect 138952 2332 139952 2360
rect 133288 2320 133294 2332
rect 103514 2292 103520 2304
rect 99116 2264 103520 2292
rect 103514 2252 103520 2264
rect 103572 2252 103578 2304
rect 104618 2252 104624 2304
rect 104676 2292 104682 2304
rect 108390 2292 108396 2304
rect 104676 2264 108396 2292
rect 104676 2252 104682 2264
rect 108390 2252 108396 2264
rect 108448 2252 108454 2304
rect 122650 2252 122656 2304
rect 122708 2252 122714 2304
rect 124766 2252 124772 2304
rect 124824 2252 124830 2304
rect 126330 2252 126336 2304
rect 126388 2252 126394 2304
rect 127802 2252 127808 2304
rect 127860 2252 127866 2304
rect 128354 2252 128360 2304
rect 128412 2292 128418 2304
rect 128541 2295 128599 2301
rect 128541 2292 128553 2295
rect 128412 2264 128553 2292
rect 128412 2252 128418 2264
rect 128541 2261 128553 2264
rect 128587 2261 128599 2295
rect 128541 2255 128599 2261
rect 130010 2252 130016 2304
rect 130068 2252 130074 2304
rect 131574 2252 131580 2304
rect 131632 2252 131638 2304
rect 132954 2252 132960 2304
rect 133012 2252 133018 2304
rect 133690 2252 133696 2304
rect 133748 2252 133754 2304
rect 134426 2252 134432 2304
rect 134484 2252 134490 2304
rect 134978 2252 134984 2304
rect 135036 2252 135042 2304
rect 137986 2292 138014 2332
rect 139946 2320 139952 2332
rect 140004 2320 140010 2372
rect 140777 2363 140835 2369
rect 140777 2329 140789 2363
rect 140823 2329 140835 2363
rect 140777 2323 140835 2329
rect 138661 2295 138719 2301
rect 138661 2292 138673 2295
rect 137986 2264 138673 2292
rect 138661 2261 138673 2264
rect 138707 2292 138719 2295
rect 140792 2292 140820 2323
rect 155770 2320 155776 2372
rect 155828 2360 155834 2372
rect 156874 2360 156880 2372
rect 155828 2332 156880 2360
rect 155828 2320 155834 2332
rect 156874 2320 156880 2332
rect 156932 2360 156938 2372
rect 156969 2363 157027 2369
rect 156969 2360 156981 2363
rect 156932 2332 156981 2360
rect 156932 2320 156938 2332
rect 156969 2329 156981 2332
rect 157015 2329 157027 2363
rect 158162 2360 158168 2372
rect 156969 2323 157027 2329
rect 157306 2332 158168 2360
rect 141145 2295 141203 2301
rect 141145 2292 141157 2295
rect 138707 2264 141157 2292
rect 138707 2261 138719 2264
rect 138661 2255 138719 2261
rect 141145 2261 141157 2264
rect 141191 2292 141203 2295
rect 141326 2292 141332 2304
rect 141191 2264 141332 2292
rect 141191 2261 141203 2264
rect 141145 2255 141203 2261
rect 141326 2252 141332 2264
rect 141384 2252 141390 2304
rect 148962 2252 148968 2304
rect 149020 2292 149026 2304
rect 156322 2292 156328 2304
rect 149020 2264 156328 2292
rect 149020 2252 149026 2264
rect 156322 2252 156328 2264
rect 156380 2252 156386 2304
rect 156506 2252 156512 2304
rect 156564 2292 156570 2304
rect 157306 2292 157334 2332
rect 158162 2320 158168 2332
rect 158220 2320 158226 2372
rect 158530 2320 158536 2372
rect 158588 2360 158594 2372
rect 159085 2363 159143 2369
rect 159085 2360 159097 2363
rect 158588 2332 159097 2360
rect 158588 2320 158594 2332
rect 159085 2329 159097 2332
rect 159131 2329 159143 2363
rect 159085 2323 159143 2329
rect 160281 2363 160339 2369
rect 160281 2329 160293 2363
rect 160327 2360 160339 2363
rect 160756 2360 160784 2391
rect 162302 2388 162308 2400
rect 162360 2388 162366 2440
rect 163685 2431 163743 2437
rect 163685 2397 163697 2431
rect 163731 2428 163743 2431
rect 163958 2428 163964 2440
rect 163731 2400 163964 2428
rect 163731 2397 163743 2400
rect 163685 2391 163743 2397
rect 163958 2388 163964 2400
rect 164016 2388 164022 2440
rect 164418 2388 164424 2440
rect 164476 2388 164482 2440
rect 165157 2431 165215 2437
rect 165157 2397 165169 2431
rect 165203 2428 165215 2431
rect 165614 2428 165620 2440
rect 165203 2400 165620 2428
rect 165203 2397 165215 2400
rect 165157 2391 165215 2397
rect 165614 2388 165620 2400
rect 165672 2388 165678 2440
rect 165890 2388 165896 2440
rect 165948 2388 165954 2440
rect 166629 2431 166687 2437
rect 166629 2397 166641 2431
rect 166675 2428 166687 2431
rect 167454 2428 167460 2440
rect 166675 2400 167460 2428
rect 166675 2397 166687 2400
rect 166629 2391 166687 2397
rect 167454 2388 167460 2400
rect 167512 2388 167518 2440
rect 167730 2388 167736 2440
rect 167788 2388 167794 2440
rect 167822 2388 167828 2440
rect 167880 2388 167886 2440
rect 176654 2388 176660 2440
rect 176712 2388 176718 2440
rect 176930 2388 176936 2440
rect 176988 2388 176994 2440
rect 179598 2388 179604 2440
rect 179656 2388 179662 2440
rect 186958 2388 186964 2440
rect 187016 2388 187022 2440
rect 187068 2428 187096 2536
rect 187252 2505 187280 2604
rect 190454 2592 190460 2644
rect 190512 2632 190518 2644
rect 190549 2635 190607 2641
rect 190549 2632 190561 2635
rect 190512 2604 190561 2632
rect 190512 2592 190518 2604
rect 190549 2601 190561 2604
rect 190595 2601 190607 2635
rect 190549 2595 190607 2601
rect 191834 2592 191840 2644
rect 191892 2632 191898 2644
rect 192021 2635 192079 2641
rect 192021 2632 192033 2635
rect 191892 2604 192033 2632
rect 191892 2592 191898 2604
rect 192021 2601 192033 2604
rect 192067 2601 192079 2635
rect 192021 2595 192079 2601
rect 202874 2592 202880 2644
rect 202932 2632 202938 2644
rect 202969 2635 203027 2641
rect 202969 2632 202981 2635
rect 202932 2604 202981 2632
rect 202932 2592 202938 2604
rect 202969 2601 202981 2604
rect 203015 2601 203027 2635
rect 211893 2635 211951 2641
rect 211893 2632 211905 2635
rect 202969 2595 203027 2601
rect 204916 2604 211905 2632
rect 187237 2499 187295 2505
rect 187237 2465 187249 2499
rect 187283 2465 187295 2499
rect 187237 2459 187295 2465
rect 201957 2499 202015 2505
rect 201957 2465 201969 2499
rect 202003 2496 202015 2499
rect 202598 2496 202604 2508
rect 202003 2468 202604 2496
rect 202003 2465 202015 2468
rect 201957 2459 202015 2465
rect 202598 2456 202604 2468
rect 202656 2456 202662 2508
rect 204916 2505 204944 2604
rect 211893 2601 211905 2604
rect 211939 2601 211951 2635
rect 211893 2595 211951 2601
rect 213178 2592 213184 2644
rect 213236 2632 213242 2644
rect 221918 2632 221924 2644
rect 213236 2604 221924 2632
rect 213236 2592 213242 2604
rect 221918 2592 221924 2604
rect 221976 2632 221982 2644
rect 224129 2635 224187 2641
rect 224129 2632 224141 2635
rect 221976 2604 224141 2632
rect 221976 2592 221982 2604
rect 224129 2601 224141 2604
rect 224175 2632 224187 2635
rect 224497 2635 224555 2641
rect 224497 2632 224509 2635
rect 224175 2604 224509 2632
rect 224175 2601 224187 2604
rect 224129 2595 224187 2601
rect 224497 2601 224509 2604
rect 224543 2601 224555 2635
rect 224497 2595 224555 2601
rect 224954 2592 224960 2644
rect 225012 2632 225018 2644
rect 225877 2635 225935 2641
rect 225877 2632 225889 2635
rect 225012 2604 225889 2632
rect 225012 2592 225018 2604
rect 225877 2601 225889 2604
rect 225923 2601 225935 2635
rect 225877 2595 225935 2601
rect 226242 2592 226248 2644
rect 226300 2632 226306 2644
rect 227165 2635 227223 2641
rect 227165 2632 227177 2635
rect 226300 2604 227177 2632
rect 226300 2592 226306 2604
rect 227165 2601 227177 2604
rect 227211 2601 227223 2635
rect 227165 2595 227223 2601
rect 227990 2592 227996 2644
rect 228048 2632 228054 2644
rect 231670 2632 231676 2644
rect 228048 2604 231676 2632
rect 228048 2592 228054 2604
rect 231670 2592 231676 2604
rect 231728 2592 231734 2644
rect 235994 2592 236000 2644
rect 236052 2592 236058 2644
rect 236730 2592 236736 2644
rect 236788 2632 236794 2644
rect 242802 2632 242808 2644
rect 236788 2604 242808 2632
rect 236788 2592 236794 2604
rect 242802 2592 242808 2604
rect 242860 2592 242866 2644
rect 258074 2592 258080 2644
rect 258132 2632 258138 2644
rect 266446 2632 266452 2644
rect 258132 2604 266452 2632
rect 258132 2592 258138 2604
rect 266446 2592 266452 2604
rect 266504 2592 266510 2644
rect 267093 2635 267151 2641
rect 267093 2601 267105 2635
rect 267139 2632 267151 2635
rect 268378 2632 268384 2644
rect 267139 2604 268384 2632
rect 267139 2601 267151 2604
rect 267093 2595 267151 2601
rect 268378 2592 268384 2604
rect 268436 2592 268442 2644
rect 210142 2524 210148 2576
rect 210200 2564 210206 2576
rect 210697 2567 210755 2573
rect 210697 2564 210709 2567
rect 210200 2536 210709 2564
rect 210200 2524 210206 2536
rect 210697 2533 210709 2536
rect 210743 2564 210755 2567
rect 210786 2564 210792 2576
rect 210743 2536 210792 2564
rect 210743 2533 210755 2536
rect 210697 2527 210755 2533
rect 210786 2524 210792 2536
rect 210844 2524 210850 2576
rect 213730 2524 213736 2576
rect 213788 2564 213794 2576
rect 243679 2567 243737 2573
rect 243679 2564 243691 2567
rect 213788 2536 221621 2564
rect 213788 2524 213794 2536
rect 204901 2499 204959 2505
rect 204901 2465 204913 2499
rect 204947 2465 204959 2499
rect 204901 2459 204959 2465
rect 205082 2456 205088 2508
rect 205140 2456 205146 2508
rect 205358 2456 205364 2508
rect 205416 2456 205422 2508
rect 208118 2456 208124 2508
rect 208176 2496 208182 2508
rect 210053 2499 210111 2505
rect 210053 2496 210065 2499
rect 208176 2468 210065 2496
rect 208176 2456 208182 2468
rect 210053 2465 210065 2468
rect 210099 2465 210111 2499
rect 210053 2459 210111 2465
rect 210973 2499 211031 2505
rect 210973 2465 210985 2499
rect 211019 2496 211031 2499
rect 216122 2496 216128 2508
rect 211019 2468 211936 2496
rect 211019 2465 211031 2468
rect 210973 2459 211031 2465
rect 189718 2428 189724 2440
rect 187068 2400 189724 2428
rect 189718 2388 189724 2400
rect 189776 2388 189782 2440
rect 190362 2388 190368 2440
rect 190420 2388 190426 2440
rect 191101 2431 191159 2437
rect 191101 2397 191113 2431
rect 191147 2428 191159 2431
rect 191374 2428 191380 2440
rect 191147 2400 191380 2428
rect 191147 2397 191159 2400
rect 191101 2391 191159 2397
rect 191374 2388 191380 2400
rect 191432 2388 191438 2440
rect 191837 2431 191895 2437
rect 191837 2397 191849 2431
rect 191883 2428 191895 2431
rect 192386 2428 192392 2440
rect 191883 2400 192392 2428
rect 191883 2397 191895 2400
rect 191837 2391 191895 2397
rect 192386 2388 192392 2400
rect 192444 2388 192450 2440
rect 194873 2431 194931 2437
rect 194873 2397 194885 2431
rect 194919 2428 194931 2431
rect 195698 2428 195704 2440
rect 194919 2400 195704 2428
rect 194919 2397 194931 2400
rect 194873 2391 194931 2397
rect 195698 2388 195704 2400
rect 195756 2388 195762 2440
rect 196250 2388 196256 2440
rect 196308 2388 196314 2440
rect 197170 2388 197176 2440
rect 197228 2388 197234 2440
rect 197262 2388 197268 2440
rect 197320 2388 197326 2440
rect 198369 2431 198427 2437
rect 198369 2397 198381 2431
rect 198415 2428 198427 2431
rect 199194 2428 199200 2440
rect 198415 2400 199200 2428
rect 198415 2397 198427 2400
rect 198369 2391 198427 2397
rect 199194 2388 199200 2400
rect 199252 2388 199258 2440
rect 199749 2431 199807 2437
rect 199749 2397 199761 2431
rect 199795 2428 199807 2431
rect 200850 2428 200856 2440
rect 199795 2400 200856 2428
rect 199795 2397 199807 2400
rect 199749 2391 199807 2397
rect 200850 2388 200856 2400
rect 200908 2388 200914 2440
rect 201218 2388 201224 2440
rect 201276 2388 201282 2440
rect 201310 2388 201316 2440
rect 201368 2428 201374 2440
rect 202141 2431 202199 2437
rect 202141 2428 202153 2431
rect 201368 2400 202153 2428
rect 201368 2388 201374 2400
rect 202141 2397 202153 2400
rect 202187 2397 202199 2431
rect 202141 2391 202199 2397
rect 202325 2431 202383 2437
rect 202325 2397 202337 2431
rect 202371 2428 202383 2431
rect 202785 2431 202843 2437
rect 202785 2428 202797 2431
rect 202371 2400 202797 2428
rect 202371 2397 202383 2400
rect 202325 2391 202383 2397
rect 202785 2397 202797 2400
rect 202831 2397 202843 2431
rect 202785 2391 202843 2397
rect 209958 2388 209964 2440
rect 210016 2428 210022 2440
rect 210237 2431 210295 2437
rect 210237 2428 210249 2431
rect 210016 2400 210249 2428
rect 210016 2388 210022 2400
rect 210237 2397 210249 2400
rect 210283 2397 210295 2431
rect 210237 2391 210295 2397
rect 211062 2388 211068 2440
rect 211120 2437 211126 2440
rect 211120 2431 211148 2437
rect 211136 2397 211148 2431
rect 211120 2391 211148 2397
rect 211120 2388 211126 2391
rect 211246 2388 211252 2440
rect 211304 2388 211310 2440
rect 211908 2428 211936 2468
rect 212460 2468 216128 2496
rect 212460 2428 212488 2468
rect 216122 2456 216128 2468
rect 216180 2456 216186 2508
rect 216217 2499 216275 2505
rect 216217 2465 216229 2499
rect 216263 2496 216275 2499
rect 216263 2468 217548 2496
rect 216263 2465 216275 2468
rect 216217 2459 216275 2465
rect 211908 2400 212488 2428
rect 214098 2388 214104 2440
rect 214156 2428 214162 2440
rect 217520 2437 217548 2468
rect 218606 2456 218612 2508
rect 218664 2496 218670 2508
rect 219529 2499 219587 2505
rect 219529 2496 219541 2499
rect 218664 2468 219541 2496
rect 218664 2456 218670 2468
rect 219529 2465 219541 2468
rect 219575 2465 219587 2499
rect 219529 2459 219587 2465
rect 220998 2456 221004 2508
rect 221056 2456 221062 2508
rect 221593 2496 221621 2536
rect 221752 2536 243691 2564
rect 221752 2496 221780 2536
rect 243679 2533 243691 2536
rect 243725 2533 243737 2567
rect 243679 2527 243737 2533
rect 255314 2524 255320 2576
rect 255372 2564 255378 2576
rect 269022 2564 269028 2576
rect 255372 2536 269028 2564
rect 255372 2524 255378 2536
rect 269022 2524 269028 2536
rect 269080 2524 269086 2576
rect 221593 2468 221780 2496
rect 221918 2456 221924 2508
rect 221976 2456 221982 2508
rect 222105 2499 222163 2505
rect 222105 2465 222117 2499
rect 222151 2496 222163 2499
rect 223209 2499 223267 2505
rect 222151 2468 223160 2496
rect 222151 2465 222163 2468
rect 222105 2459 222163 2465
rect 216033 2431 216091 2437
rect 216033 2428 216045 2431
rect 214156 2400 216045 2428
rect 214156 2388 214162 2400
rect 216033 2397 216045 2400
rect 216079 2397 216091 2431
rect 216033 2391 216091 2397
rect 217321 2431 217379 2437
rect 217321 2397 217333 2431
rect 217367 2397 217379 2431
rect 217321 2391 217379 2397
rect 217505 2431 217563 2437
rect 217505 2397 217517 2431
rect 217551 2428 217563 2431
rect 218054 2428 218060 2440
rect 217551 2400 218060 2428
rect 217551 2397 217563 2400
rect 217505 2391 217563 2397
rect 160327 2332 160784 2360
rect 160327 2329 160339 2332
rect 160281 2323 160339 2329
rect 161658 2320 161664 2372
rect 161716 2360 161722 2372
rect 167546 2360 167552 2372
rect 161716 2332 167552 2360
rect 161716 2320 161722 2332
rect 167546 2320 167552 2332
rect 167604 2320 167610 2372
rect 168190 2320 168196 2372
rect 168248 2360 168254 2372
rect 174722 2360 174728 2372
rect 168248 2332 174728 2360
rect 168248 2320 168254 2332
rect 174722 2320 174728 2332
rect 174780 2320 174786 2372
rect 216953 2363 217011 2369
rect 216953 2360 216965 2363
rect 215266 2332 216965 2360
rect 156564 2264 157334 2292
rect 156564 2252 156570 2264
rect 157426 2252 157432 2304
rect 157484 2292 157490 2304
rect 157521 2295 157579 2301
rect 157521 2292 157533 2295
rect 157484 2264 157533 2292
rect 157484 2252 157490 2264
rect 157521 2261 157533 2264
rect 157567 2261 157579 2295
rect 157521 2255 157579 2261
rect 160922 2252 160928 2304
rect 160980 2252 160986 2304
rect 161750 2252 161756 2304
rect 161808 2252 161814 2304
rect 162118 2252 162124 2304
rect 162176 2292 162182 2304
rect 162486 2292 162492 2304
rect 162176 2264 162492 2292
rect 162176 2252 162182 2264
rect 162486 2252 162492 2264
rect 162544 2252 162550 2304
rect 163866 2252 163872 2304
rect 163924 2252 163930 2304
rect 164234 2252 164240 2304
rect 164292 2292 164298 2304
rect 164605 2295 164663 2301
rect 164605 2292 164617 2295
rect 164292 2264 164617 2292
rect 164292 2252 164298 2264
rect 164605 2261 164617 2264
rect 164651 2261 164663 2295
rect 164605 2255 164663 2261
rect 165338 2252 165344 2304
rect 165396 2252 165402 2304
rect 166074 2252 166080 2304
rect 166132 2252 166138 2304
rect 166810 2252 166816 2304
rect 166868 2252 166874 2304
rect 168006 2252 168012 2304
rect 168064 2252 168070 2304
rect 173802 2252 173808 2304
rect 173860 2292 173866 2304
rect 183554 2292 183560 2304
rect 173860 2264 183560 2292
rect 173860 2252 173866 2264
rect 183554 2252 183560 2264
rect 183612 2252 183618 2304
rect 191282 2252 191288 2304
rect 191340 2252 191346 2304
rect 194686 2252 194692 2304
rect 194744 2292 194750 2304
rect 195057 2295 195115 2301
rect 195057 2292 195069 2295
rect 194744 2264 195069 2292
rect 194744 2252 194750 2264
rect 195057 2261 195069 2264
rect 195103 2261 195115 2295
rect 195057 2255 195115 2261
rect 195974 2252 195980 2304
rect 196032 2292 196038 2304
rect 196437 2295 196495 2301
rect 196437 2292 196449 2295
rect 196032 2264 196449 2292
rect 196032 2252 196038 2264
rect 196437 2261 196449 2264
rect 196483 2261 196495 2295
rect 196437 2255 196495 2261
rect 197446 2252 197452 2304
rect 197504 2252 197510 2304
rect 198550 2252 198556 2304
rect 198608 2252 198614 2304
rect 199930 2252 199936 2304
rect 199988 2252 199994 2304
rect 201402 2252 201408 2304
rect 201460 2252 201466 2304
rect 204254 2252 204260 2304
rect 204312 2292 204318 2304
rect 205358 2292 205364 2304
rect 204312 2264 205364 2292
rect 204312 2252 204318 2264
rect 205358 2252 205364 2264
rect 205416 2292 205422 2304
rect 207014 2292 207020 2304
rect 205416 2264 207020 2292
rect 205416 2252 205422 2264
rect 207014 2252 207020 2264
rect 207072 2252 207078 2304
rect 207106 2252 207112 2304
rect 207164 2292 207170 2304
rect 213178 2292 213184 2304
rect 207164 2264 213184 2292
rect 207164 2252 207170 2264
rect 213178 2252 213184 2264
rect 213236 2252 213242 2304
rect 213270 2252 213276 2304
rect 213328 2292 213334 2304
rect 215266 2292 215294 2332
rect 216953 2329 216965 2332
rect 216999 2360 217011 2363
rect 217336 2360 217364 2391
rect 218054 2388 218060 2400
rect 218112 2428 218118 2440
rect 218793 2431 218851 2437
rect 218793 2428 218805 2431
rect 218112 2400 218805 2428
rect 218112 2388 218118 2400
rect 218793 2397 218805 2400
rect 218839 2428 218851 2431
rect 219066 2428 219072 2440
rect 218839 2400 219072 2428
rect 218839 2397 218851 2400
rect 218793 2391 218851 2397
rect 219066 2388 219072 2400
rect 219124 2388 219130 2440
rect 220817 2431 220875 2437
rect 220817 2397 220829 2431
rect 220863 2397 220875 2431
rect 220817 2391 220875 2397
rect 218241 2363 218299 2369
rect 218241 2360 218253 2363
rect 216999 2332 218253 2360
rect 216999 2329 217011 2332
rect 216953 2323 217011 2329
rect 218241 2329 218253 2332
rect 218287 2329 218299 2363
rect 218241 2323 218299 2329
rect 219253 2363 219311 2369
rect 219253 2329 219265 2363
rect 219299 2360 219311 2363
rect 220722 2360 220728 2372
rect 219299 2332 220728 2360
rect 219299 2329 219311 2332
rect 219253 2323 219311 2329
rect 220722 2320 220728 2332
rect 220780 2320 220786 2372
rect 213328 2264 215294 2292
rect 213328 2252 213334 2264
rect 216398 2252 216404 2304
rect 216456 2292 216462 2304
rect 216677 2295 216735 2301
rect 216677 2292 216689 2295
rect 216456 2264 216689 2292
rect 216456 2252 216462 2264
rect 216677 2261 216689 2264
rect 216723 2261 216735 2295
rect 216677 2255 216735 2261
rect 217965 2295 218023 2301
rect 217965 2261 217977 2295
rect 218011 2292 218023 2295
rect 218146 2292 218152 2304
rect 218011 2264 218152 2292
rect 218011 2261 218023 2264
rect 217965 2255 218023 2261
rect 218146 2252 218152 2264
rect 218204 2252 218210 2304
rect 219802 2252 219808 2304
rect 219860 2292 219866 2304
rect 220449 2295 220507 2301
rect 220449 2292 220461 2295
rect 219860 2264 220461 2292
rect 219860 2252 219866 2264
rect 220449 2261 220461 2264
rect 220495 2292 220507 2295
rect 220832 2292 220860 2391
rect 221366 2388 221372 2440
rect 221424 2428 221430 2440
rect 222841 2431 222899 2437
rect 222841 2428 222853 2431
rect 221424 2400 222853 2428
rect 221424 2388 221430 2400
rect 222841 2397 222853 2400
rect 222887 2397 222899 2431
rect 222841 2391 222899 2397
rect 223022 2388 223028 2440
rect 223080 2388 223086 2440
rect 223132 2428 223160 2468
rect 223209 2465 223221 2499
rect 223255 2496 223267 2499
rect 223574 2496 223580 2508
rect 223255 2468 223580 2496
rect 223255 2465 223267 2468
rect 223209 2459 223267 2465
rect 223574 2456 223580 2468
rect 223632 2456 223638 2508
rect 246669 2499 246727 2505
rect 246669 2496 246681 2499
rect 224926 2468 246681 2496
rect 223666 2428 223672 2440
rect 223132 2400 223672 2428
rect 223666 2388 223672 2400
rect 223724 2388 223730 2440
rect 224926 2428 224954 2468
rect 246669 2465 246681 2468
rect 246715 2465 246727 2499
rect 246669 2459 246727 2465
rect 258718 2456 258724 2508
rect 258776 2496 258782 2508
rect 258905 2499 258963 2505
rect 258905 2496 258917 2499
rect 258776 2468 258917 2496
rect 258776 2456 258782 2468
rect 258905 2465 258917 2468
rect 258951 2465 258963 2499
rect 270126 2496 270132 2508
rect 258905 2459 258963 2465
rect 269132 2468 270132 2496
rect 223776 2400 224954 2428
rect 221642 2320 221648 2372
rect 221700 2360 221706 2372
rect 223776 2360 223804 2400
rect 225322 2388 225328 2440
rect 225380 2388 225386 2440
rect 225693 2431 225751 2437
rect 225693 2397 225705 2431
rect 225739 2428 225751 2431
rect 226150 2428 226156 2440
rect 225739 2400 226156 2428
rect 225739 2397 225751 2400
rect 225693 2391 225751 2397
rect 226150 2388 226156 2400
rect 226208 2388 226214 2440
rect 226242 2388 226248 2440
rect 226300 2388 226306 2440
rect 226978 2388 226984 2440
rect 227036 2388 227042 2440
rect 227622 2388 227628 2440
rect 227680 2428 227686 2440
rect 227901 2431 227959 2437
rect 227901 2428 227913 2431
rect 227680 2400 227913 2428
rect 227680 2388 227686 2400
rect 227901 2397 227913 2400
rect 227947 2397 227959 2431
rect 227901 2391 227959 2397
rect 228177 2431 228235 2437
rect 228177 2397 228189 2431
rect 228223 2428 228235 2431
rect 228358 2428 228364 2440
rect 228223 2400 228364 2428
rect 228223 2397 228235 2400
rect 228177 2391 228235 2397
rect 228358 2388 228364 2400
rect 228416 2388 228422 2440
rect 228818 2388 228824 2440
rect 228876 2388 228882 2440
rect 231121 2431 231179 2437
rect 231121 2397 231133 2431
rect 231167 2428 231179 2431
rect 231762 2428 231768 2440
rect 231167 2400 231768 2428
rect 231167 2397 231179 2400
rect 231121 2391 231179 2397
rect 231762 2388 231768 2400
rect 231820 2388 231826 2440
rect 231854 2388 231860 2440
rect 231912 2388 231918 2440
rect 232590 2388 232596 2440
rect 232648 2388 232654 2440
rect 235813 2431 235871 2437
rect 235813 2397 235825 2431
rect 235859 2428 235871 2431
rect 236086 2428 236092 2440
rect 235859 2400 236092 2428
rect 235859 2397 235871 2400
rect 235813 2391 235871 2397
rect 236086 2388 236092 2400
rect 236144 2388 236150 2440
rect 236546 2388 236552 2440
rect 236604 2388 236610 2440
rect 243446 2388 243452 2440
rect 243504 2388 243510 2440
rect 246390 2388 246396 2440
rect 246448 2388 246454 2440
rect 256694 2388 256700 2440
rect 256752 2388 256758 2440
rect 256970 2388 256976 2440
rect 257028 2388 257034 2440
rect 259086 2388 259092 2440
rect 259144 2388 259150 2440
rect 259273 2431 259331 2437
rect 259273 2397 259285 2431
rect 259319 2428 259331 2431
rect 259733 2431 259791 2437
rect 259733 2428 259745 2431
rect 259319 2400 259745 2428
rect 259319 2397 259331 2400
rect 259273 2391 259331 2397
rect 259733 2397 259745 2400
rect 259779 2397 259791 2431
rect 259733 2391 259791 2397
rect 261570 2388 261576 2440
rect 261628 2388 261634 2440
rect 263962 2388 263968 2440
rect 264020 2388 264026 2440
rect 264149 2431 264207 2437
rect 264149 2397 264161 2431
rect 264195 2428 264207 2431
rect 264238 2428 264244 2440
rect 264195 2400 264244 2428
rect 264195 2397 264207 2400
rect 264149 2391 264207 2397
rect 264238 2388 264244 2400
rect 264296 2388 264302 2440
rect 264333 2431 264391 2437
rect 264333 2397 264345 2431
rect 264379 2428 264391 2431
rect 264793 2431 264851 2437
rect 264793 2428 264805 2431
rect 264379 2400 264805 2428
rect 264379 2397 264391 2400
rect 264333 2391 264391 2397
rect 264793 2397 264805 2400
rect 264839 2397 264851 2431
rect 264793 2391 264851 2397
rect 267274 2390 267280 2442
rect 267332 2390 267338 2442
rect 267921 2431 267979 2437
rect 267921 2397 267933 2431
rect 267967 2397 267979 2431
rect 267921 2391 267979 2397
rect 221700 2332 223804 2360
rect 221700 2320 221706 2332
rect 224034 2320 224040 2372
rect 224092 2360 224098 2372
rect 224092 2332 225552 2360
rect 224092 2320 224098 2332
rect 221366 2292 221372 2304
rect 220495 2264 221372 2292
rect 220495 2261 220507 2264
rect 220449 2255 220507 2261
rect 221366 2252 221372 2264
rect 221424 2252 221430 2304
rect 221461 2295 221519 2301
rect 221461 2261 221473 2295
rect 221507 2292 221519 2295
rect 222470 2292 222476 2304
rect 221507 2264 222476 2292
rect 221507 2261 221519 2264
rect 221461 2255 221519 2261
rect 222470 2252 222476 2264
rect 222528 2252 222534 2304
rect 222562 2252 222568 2304
rect 222620 2252 222626 2304
rect 223669 2295 223727 2301
rect 223669 2261 223681 2295
rect 223715 2292 223727 2295
rect 223758 2292 223764 2304
rect 223715 2264 223764 2292
rect 223715 2261 223727 2264
rect 223669 2255 223727 2261
rect 223758 2252 223764 2264
rect 223816 2252 223822 2304
rect 224218 2252 224224 2304
rect 224276 2292 224282 2304
rect 225524 2301 225552 2332
rect 227806 2320 227812 2372
rect 227864 2360 227870 2372
rect 237190 2360 237196 2372
rect 227864 2332 237196 2360
rect 227864 2320 227870 2332
rect 237190 2320 237196 2332
rect 237248 2320 237254 2372
rect 258074 2320 258080 2372
rect 258132 2320 258138 2372
rect 264422 2320 264428 2372
rect 264480 2360 264486 2372
rect 267936 2360 267964 2391
rect 268562 2388 268568 2440
rect 268620 2388 268626 2440
rect 269132 2437 269160 2468
rect 270126 2456 270132 2468
rect 270184 2456 270190 2508
rect 269117 2431 269175 2437
rect 269117 2397 269129 2431
rect 269163 2397 269175 2431
rect 269117 2391 269175 2397
rect 269206 2388 269212 2440
rect 269264 2388 269270 2440
rect 269666 2388 269672 2440
rect 269724 2428 269730 2440
rect 269853 2431 269911 2437
rect 269853 2428 269865 2431
rect 269724 2400 269865 2428
rect 269724 2388 269730 2400
rect 269853 2397 269865 2400
rect 269899 2397 269911 2431
rect 269853 2391 269911 2397
rect 270494 2388 270500 2440
rect 270552 2428 270558 2440
rect 270589 2431 270647 2437
rect 270589 2428 270601 2431
rect 270552 2400 270601 2428
rect 270552 2388 270558 2400
rect 270589 2397 270601 2400
rect 270635 2397 270647 2431
rect 270589 2391 270647 2397
rect 268838 2360 268844 2372
rect 264480 2332 267780 2360
rect 267936 2332 268844 2360
rect 264480 2320 264486 2332
rect 224957 2295 225015 2301
rect 224957 2292 224969 2295
rect 224276 2264 224969 2292
rect 224276 2252 224282 2264
rect 224957 2261 224969 2264
rect 225003 2261 225015 2295
rect 224957 2255 225015 2261
rect 225509 2295 225567 2301
rect 225509 2261 225521 2295
rect 225555 2261 225567 2295
rect 225509 2255 225567 2261
rect 225598 2252 225604 2304
rect 225656 2292 225662 2304
rect 226429 2295 226487 2301
rect 226429 2292 226441 2295
rect 225656 2264 226441 2292
rect 225656 2252 225662 2264
rect 226429 2261 226441 2264
rect 226475 2261 226487 2295
rect 226429 2255 226487 2261
rect 226702 2252 226708 2304
rect 226760 2292 226766 2304
rect 227162 2292 227168 2304
rect 226760 2264 227168 2292
rect 226760 2252 226766 2264
rect 227162 2252 227168 2264
rect 227220 2252 227226 2304
rect 228450 2252 228456 2304
rect 228508 2292 228514 2304
rect 229005 2295 229063 2301
rect 229005 2292 229017 2295
rect 228508 2264 229017 2292
rect 228508 2252 228514 2264
rect 229005 2261 229017 2264
rect 229051 2261 229063 2295
rect 229005 2255 229063 2261
rect 231302 2252 231308 2304
rect 231360 2252 231366 2304
rect 232038 2252 232044 2304
rect 232096 2252 232102 2304
rect 232774 2252 232780 2304
rect 232832 2252 232838 2304
rect 236730 2252 236736 2304
rect 236788 2252 236794 2304
rect 244274 2252 244280 2304
rect 244332 2292 244338 2304
rect 255406 2292 255412 2304
rect 244332 2264 255412 2292
rect 244332 2252 244338 2264
rect 255406 2252 255412 2264
rect 255464 2252 255470 2304
rect 257706 2252 257712 2304
rect 257764 2292 257770 2304
rect 257890 2292 257896 2304
rect 257764 2264 257896 2292
rect 257764 2252 257770 2264
rect 257890 2252 257896 2264
rect 257948 2292 257954 2304
rect 258169 2295 258227 2301
rect 258169 2292 258181 2295
rect 257948 2264 258181 2292
rect 257948 2252 257954 2264
rect 258169 2261 258181 2264
rect 258215 2261 258227 2295
rect 258169 2255 258227 2261
rect 259914 2252 259920 2304
rect 259972 2252 259978 2304
rect 261757 2295 261815 2301
rect 261757 2261 261769 2295
rect 261803 2292 261815 2295
rect 261846 2292 261852 2304
rect 261803 2264 261852 2292
rect 261803 2261 261815 2264
rect 261757 2255 261815 2261
rect 261846 2252 261852 2264
rect 261904 2252 261910 2304
rect 264974 2252 264980 2304
rect 265032 2252 265038 2304
rect 265989 2295 266047 2301
rect 265989 2261 266001 2295
rect 266035 2292 266047 2295
rect 267550 2292 267556 2304
rect 266035 2264 267556 2292
rect 266035 2261 266047 2264
rect 265989 2255 266047 2261
rect 267550 2252 267556 2264
rect 267608 2252 267614 2304
rect 267752 2301 267780 2332
rect 268838 2320 268844 2332
rect 268896 2320 268902 2372
rect 267737 2295 267795 2301
rect 267737 2261 267749 2295
rect 267783 2261 267795 2295
rect 267737 2255 267795 2261
rect 268194 2252 268200 2304
rect 268252 2292 268258 2304
rect 268381 2295 268439 2301
rect 268381 2292 268393 2295
rect 268252 2264 268393 2292
rect 268252 2252 268258 2264
rect 268381 2261 268393 2264
rect 268427 2261 268439 2295
rect 268381 2255 268439 2261
rect 269393 2295 269451 2301
rect 269393 2261 269405 2295
rect 269439 2292 269451 2295
rect 269942 2292 269948 2304
rect 269439 2264 269948 2292
rect 269439 2261 269451 2264
rect 269393 2255 269451 2261
rect 269942 2252 269948 2264
rect 270000 2252 270006 2304
rect 270034 2252 270040 2304
rect 270092 2252 270098 2304
rect 270770 2252 270776 2304
rect 270828 2252 270834 2304
rect 1104 2202 271651 2224
rect 1104 2150 68546 2202
rect 68598 2150 68610 2202
rect 68662 2150 68674 2202
rect 68726 2150 68738 2202
rect 68790 2150 68802 2202
rect 68854 2150 136143 2202
rect 136195 2150 136207 2202
rect 136259 2150 136271 2202
rect 136323 2150 136335 2202
rect 136387 2150 136399 2202
rect 136451 2150 203740 2202
rect 203792 2150 203804 2202
rect 203856 2150 203868 2202
rect 203920 2150 203932 2202
rect 203984 2150 203996 2202
rect 204048 2150 271337 2202
rect 271389 2150 271401 2202
rect 271453 2150 271465 2202
rect 271517 2150 271529 2202
rect 271581 2150 271593 2202
rect 271645 2150 271651 2202
rect 1104 2128 271651 2150
rect 6917 2091 6975 2097
rect 6917 2057 6929 2091
rect 6963 2088 6975 2091
rect 6963 2060 22094 2088
rect 6963 2057 6975 2060
rect 6917 2051 6975 2057
rect 9214 1980 9220 2032
rect 9272 1980 9278 2032
rect 17126 1980 17132 2032
rect 17184 1980 17190 2032
rect 22066 2020 22094 2060
rect 23842 2048 23848 2100
rect 23900 2048 23906 2100
rect 26326 2048 26332 2100
rect 26384 2048 26390 2100
rect 26528 2060 57468 2088
rect 25130 2020 25136 2032
rect 22066 1992 25136 2020
rect 25130 1980 25136 1992
rect 25188 1980 25194 2032
rect 25225 2023 25283 2029
rect 25225 1989 25237 2023
rect 25271 2020 25283 2023
rect 25590 2020 25596 2032
rect 25271 1992 25596 2020
rect 25271 1989 25283 1992
rect 25225 1983 25283 1989
rect 25590 1980 25596 1992
rect 25648 1980 25654 2032
rect 26237 2023 26295 2029
rect 26237 1989 26249 2023
rect 26283 2020 26295 2023
rect 26418 2020 26424 2032
rect 26283 1992 26424 2020
rect 26283 1989 26295 1992
rect 26237 1983 26295 1989
rect 26418 1980 26424 1992
rect 26476 1980 26482 2032
rect 2590 1912 2596 1964
rect 2648 1912 2654 1964
rect 4798 1912 4804 1964
rect 4856 1912 4862 1964
rect 6822 1912 6828 1964
rect 6880 1912 6886 1964
rect 7558 1912 7564 1964
rect 7616 1912 7622 1964
rect 9030 1912 9036 1964
rect 9088 1912 9094 1964
rect 14366 1912 14372 1964
rect 14424 1912 14430 1964
rect 15654 1912 15660 1964
rect 15712 1912 15718 1964
rect 15838 1912 15844 1964
rect 15896 1912 15902 1964
rect 16574 1912 16580 1964
rect 16632 1952 16638 1964
rect 16945 1955 17003 1961
rect 16945 1952 16957 1955
rect 16632 1924 16957 1952
rect 16632 1912 16638 1924
rect 16945 1921 16957 1924
rect 16991 1921 17003 1955
rect 16945 1915 17003 1921
rect 23566 1912 23572 1964
rect 23624 1912 23630 1964
rect 23661 1955 23719 1961
rect 23661 1921 23673 1955
rect 23707 1921 23719 1955
rect 23661 1915 23719 1921
rect 2314 1844 2320 1896
rect 2372 1844 2378 1896
rect 4522 1844 4528 1896
rect 4580 1844 4586 1896
rect 14090 1844 14096 1896
rect 14148 1844 14154 1896
rect 23676 1884 23704 1915
rect 23934 1912 23940 1964
rect 23992 1952 23998 1964
rect 24305 1955 24363 1961
rect 24305 1952 24317 1955
rect 23992 1924 24317 1952
rect 23992 1912 23998 1924
rect 24305 1921 24317 1924
rect 24351 1921 24363 1955
rect 24305 1915 24363 1921
rect 24489 1955 24547 1961
rect 24489 1921 24501 1955
rect 24535 1921 24547 1955
rect 24489 1915 24547 1921
rect 24504 1884 24532 1915
rect 24946 1912 24952 1964
rect 25004 1952 25010 1964
rect 25682 1952 25688 1964
rect 25004 1924 25688 1952
rect 25004 1912 25010 1924
rect 25682 1912 25688 1924
rect 25740 1952 25746 1964
rect 26528 1952 26556 2060
rect 27249 2023 27307 2029
rect 27249 1989 27261 2023
rect 27295 2020 27307 2023
rect 27706 2020 27712 2032
rect 27295 1992 27712 2020
rect 27295 1989 27307 1992
rect 27249 1983 27307 1989
rect 27706 1980 27712 1992
rect 27764 1980 27770 2032
rect 27890 1980 27896 2032
rect 27948 2020 27954 2032
rect 33042 2020 33048 2032
rect 27948 1992 31616 2020
rect 27948 1980 27954 1992
rect 25740 1924 26556 1952
rect 25740 1912 25746 1924
rect 28442 1912 28448 1964
rect 28500 1952 28506 1964
rect 28828 1961 28856 1992
rect 28629 1955 28687 1961
rect 28629 1952 28641 1955
rect 28500 1924 28641 1952
rect 28500 1912 28506 1924
rect 28629 1921 28641 1924
rect 28675 1921 28687 1955
rect 28629 1915 28687 1921
rect 28813 1955 28871 1961
rect 28813 1921 28825 1955
rect 28859 1921 28871 1955
rect 28813 1915 28871 1921
rect 29546 1912 29552 1964
rect 29604 1912 29610 1964
rect 29656 1961 29684 1992
rect 29641 1955 29699 1961
rect 29641 1921 29653 1955
rect 29687 1921 29699 1955
rect 29641 1915 29699 1921
rect 30374 1912 30380 1964
rect 30432 1912 30438 1964
rect 30576 1961 30604 1992
rect 30561 1955 30619 1961
rect 30561 1921 30573 1955
rect 30607 1921 30619 1955
rect 30561 1915 30619 1921
rect 31202 1912 31208 1964
rect 31260 1952 31266 1964
rect 31588 1961 31616 1992
rect 32416 1992 33048 2020
rect 32416 1961 32444 1992
rect 33042 1980 33048 1992
rect 33100 1980 33106 2032
rect 35526 1980 35532 2032
rect 35584 1980 35590 2032
rect 35802 1980 35808 2032
rect 35860 1980 35866 2032
rect 36265 2023 36323 2029
rect 36265 1989 36277 2023
rect 36311 2020 36323 2023
rect 36354 2020 36360 2032
rect 36311 1992 36360 2020
rect 36311 1989 36323 1992
rect 36265 1983 36323 1989
rect 36354 1980 36360 1992
rect 36412 1980 36418 2032
rect 36630 1980 36636 2032
rect 36688 1980 36694 2032
rect 37274 1980 37280 2032
rect 37332 2020 37338 2032
rect 37332 1992 38332 2020
rect 37332 1980 37338 1992
rect 31389 1955 31447 1961
rect 31389 1952 31401 1955
rect 31260 1924 31401 1952
rect 31260 1912 31266 1924
rect 31389 1921 31401 1924
rect 31435 1921 31447 1955
rect 31389 1915 31447 1921
rect 31573 1955 31631 1961
rect 31573 1921 31585 1955
rect 31619 1952 31631 1955
rect 32401 1955 32459 1961
rect 31619 1924 31754 1952
rect 31619 1921 31631 1924
rect 31573 1915 31631 1921
rect 25038 1884 25044 1896
rect 23676 1856 25044 1884
rect 25038 1844 25044 1856
rect 25096 1844 25102 1896
rect 25130 1844 25136 1896
rect 25188 1884 25194 1896
rect 31018 1884 31024 1896
rect 25188 1856 31024 1884
rect 25188 1844 25194 1856
rect 31018 1844 31024 1856
rect 31076 1844 31082 1896
rect 31726 1884 31754 1924
rect 32401 1921 32413 1955
rect 32447 1921 32459 1955
rect 32401 1915 32459 1921
rect 32490 1912 32496 1964
rect 32548 1912 32554 1964
rect 32677 1955 32735 1961
rect 32677 1921 32689 1955
rect 32723 1952 32735 1955
rect 33137 1955 33195 1961
rect 33137 1952 33149 1955
rect 32723 1924 33149 1952
rect 32723 1921 32735 1924
rect 32677 1915 32735 1921
rect 33137 1921 33149 1924
rect 33183 1921 33195 1955
rect 33137 1915 33195 1921
rect 35897 1955 35955 1961
rect 35897 1921 35909 1955
rect 35943 1952 35955 1955
rect 37292 1952 37320 1980
rect 38304 1964 38332 1992
rect 38654 1980 38660 2032
rect 38712 2020 38718 2032
rect 39025 2023 39083 2029
rect 39025 2020 39037 2023
rect 38712 1992 39037 2020
rect 38712 1980 38718 1992
rect 39025 1989 39037 1992
rect 39071 1989 39083 2023
rect 39025 1983 39083 1989
rect 39298 1980 39304 2032
rect 39356 1980 39362 2032
rect 39758 1980 39764 2032
rect 39816 1980 39822 2032
rect 40034 2020 40040 2032
rect 39868 1992 40040 2020
rect 35943 1924 37320 1952
rect 35943 1921 35955 1924
rect 35897 1915 35955 1921
rect 38102 1912 38108 1964
rect 38160 1912 38166 1964
rect 38286 1912 38292 1964
rect 38344 1952 38350 1964
rect 39393 1955 39451 1961
rect 39393 1952 39405 1955
rect 38344 1924 39405 1952
rect 38344 1912 38350 1924
rect 39393 1921 39405 1924
rect 39439 1952 39451 1955
rect 39868 1952 39896 1992
rect 40034 1980 40040 1992
rect 40092 1980 40098 2032
rect 40126 1980 40132 2032
rect 40184 1980 40190 2032
rect 54202 1980 54208 2032
rect 54260 1980 54266 2032
rect 55030 1980 55036 2032
rect 55088 1980 55094 2032
rect 57440 2020 57468 2060
rect 57514 2048 57520 2100
rect 57572 2048 57578 2100
rect 58526 2048 58532 2100
rect 58584 2048 58590 2100
rect 59262 2048 59268 2100
rect 59320 2048 59326 2100
rect 62666 2048 62672 2100
rect 62724 2048 62730 2100
rect 65242 2048 65248 2100
rect 65300 2048 65306 2100
rect 91002 2088 91008 2100
rect 76024 2060 91008 2088
rect 58544 2020 58572 2048
rect 55324 1992 57376 2020
rect 57440 1992 58572 2020
rect 39439 1924 39896 1952
rect 39439 1921 39451 1924
rect 39393 1915 39451 1921
rect 39942 1912 39948 1964
rect 40000 1912 40006 1964
rect 45462 1912 45468 1964
rect 45520 1912 45526 1964
rect 50614 1912 50620 1964
rect 50672 1912 50678 1964
rect 52914 1912 52920 1964
rect 52972 1912 52978 1964
rect 54018 1912 54024 1964
rect 54076 1952 54082 1964
rect 54849 1955 54907 1961
rect 55324 1958 55352 1992
rect 54849 1952 54861 1955
rect 54076 1924 54861 1952
rect 54076 1912 54082 1924
rect 54849 1921 54861 1924
rect 54895 1952 54907 1955
rect 55232 1952 55352 1958
rect 54895 1930 55352 1952
rect 54895 1924 55260 1930
rect 54895 1921 54907 1924
rect 54849 1915 54907 1921
rect 55398 1912 55404 1964
rect 55456 1952 55462 1964
rect 55692 1961 55720 1992
rect 55493 1955 55551 1961
rect 55493 1952 55505 1955
rect 55456 1924 55505 1952
rect 55456 1912 55462 1924
rect 55493 1921 55505 1924
rect 55539 1921 55551 1955
rect 55493 1915 55551 1921
rect 55677 1955 55735 1961
rect 55677 1921 55689 1955
rect 55723 1921 55735 1955
rect 55677 1915 55735 1921
rect 56318 1912 56324 1964
rect 56376 1912 56382 1964
rect 56520 1961 56548 1992
rect 56505 1955 56563 1961
rect 56505 1921 56517 1955
rect 56551 1921 56563 1955
rect 56505 1915 56563 1921
rect 57146 1912 57152 1964
rect 57204 1912 57210 1964
rect 57348 1961 57376 1992
rect 57333 1955 57391 1961
rect 57333 1921 57345 1955
rect 57379 1952 57391 1955
rect 58069 1955 58127 1961
rect 58069 1952 58081 1955
rect 57379 1924 58081 1952
rect 57379 1921 57391 1924
rect 57333 1915 57391 1921
rect 58069 1921 58081 1924
rect 58115 1952 58127 1955
rect 59081 1955 59139 1961
rect 59081 1952 59093 1955
rect 58115 1924 59093 1952
rect 58115 1921 58127 1924
rect 58069 1915 58127 1921
rect 59081 1921 59093 1924
rect 59127 1921 59139 1955
rect 59081 1915 59139 1921
rect 32508 1884 32536 1912
rect 37182 1884 37188 1896
rect 31726 1856 32536 1884
rect 36570 1856 37188 1884
rect 37182 1844 37188 1856
rect 37240 1844 37246 1896
rect 39960 1870 39988 1912
rect 53466 1844 53472 1896
rect 53524 1884 53530 1896
rect 53837 1887 53895 1893
rect 53837 1884 53849 1887
rect 53524 1856 53849 1884
rect 53524 1844 53530 1856
rect 53837 1853 53849 1856
rect 53883 1853 53895 1887
rect 53837 1847 53895 1853
rect 54386 1844 54392 1896
rect 54444 1884 54450 1896
rect 54665 1887 54723 1893
rect 54665 1884 54677 1887
rect 54444 1856 54677 1884
rect 54444 1844 54450 1856
rect 54665 1853 54677 1856
rect 54711 1853 54723 1887
rect 54665 1847 54723 1853
rect 57885 1887 57943 1893
rect 57885 1853 57897 1887
rect 57931 1884 57943 1887
rect 58526 1884 58532 1896
rect 57931 1856 58532 1884
rect 57931 1853 57943 1856
rect 57885 1847 57943 1853
rect 58526 1844 58532 1856
rect 58584 1844 58590 1896
rect 58894 1844 58900 1896
rect 58952 1844 58958 1896
rect 59096 1884 59124 1915
rect 59814 1912 59820 1964
rect 59872 1912 59878 1964
rect 60001 1955 60059 1961
rect 60001 1921 60013 1955
rect 60047 1921 60059 1955
rect 60001 1915 60059 1921
rect 59906 1884 59912 1896
rect 59096 1856 59912 1884
rect 59906 1844 59912 1856
rect 59964 1884 59970 1896
rect 60016 1884 60044 1915
rect 60642 1912 60648 1964
rect 60700 1912 60706 1964
rect 60829 1955 60887 1961
rect 60829 1921 60841 1955
rect 60875 1921 60887 1955
rect 60829 1915 60887 1921
rect 60844 1884 60872 1915
rect 61562 1912 61568 1964
rect 61620 1912 61626 1964
rect 61657 1955 61715 1961
rect 61657 1921 61669 1955
rect 61703 1921 61715 1955
rect 61657 1915 61715 1921
rect 61672 1884 61700 1915
rect 62390 1912 62396 1964
rect 62448 1912 62454 1964
rect 62485 1955 62543 1961
rect 62485 1921 62497 1955
rect 62531 1921 62543 1955
rect 62485 1915 62543 1921
rect 62500 1884 62528 1915
rect 63218 1912 63224 1964
rect 63276 1912 63282 1964
rect 63405 1955 63463 1961
rect 63405 1921 63417 1955
rect 63451 1921 63463 1955
rect 63405 1915 63463 1921
rect 63420 1884 63448 1915
rect 64046 1912 64052 1964
rect 64104 1912 64110 1964
rect 64233 1955 64291 1961
rect 64233 1921 64245 1955
rect 64279 1952 64291 1955
rect 65061 1955 65119 1961
rect 65061 1952 65073 1955
rect 64279 1924 65073 1952
rect 64279 1921 64291 1924
rect 64233 1915 64291 1921
rect 65061 1921 65073 1924
rect 65107 1921 65119 1955
rect 65061 1915 65119 1921
rect 64248 1884 64276 1915
rect 59964 1856 64276 1884
rect 59964 1844 59970 1856
rect 64874 1844 64880 1896
rect 64932 1844 64938 1896
rect 65076 1884 65104 1915
rect 65702 1912 65708 1964
rect 65760 1912 65766 1964
rect 65889 1955 65947 1961
rect 65889 1921 65901 1955
rect 65935 1921 65947 1955
rect 65889 1915 65947 1921
rect 65904 1884 65932 1915
rect 66622 1912 66628 1964
rect 66680 1912 66686 1964
rect 66714 1912 66720 1964
rect 66772 1912 66778 1964
rect 66901 1955 66959 1961
rect 66901 1921 66913 1955
rect 66947 1952 66959 1955
rect 67361 1955 67419 1961
rect 67361 1952 67373 1955
rect 66947 1924 67373 1952
rect 66947 1921 66959 1924
rect 66901 1915 66959 1921
rect 67361 1921 67373 1924
rect 67407 1921 67419 1955
rect 67361 1915 67419 1921
rect 70854 1912 70860 1964
rect 70912 1912 70918 1964
rect 72326 1912 72332 1964
rect 72384 1912 72390 1964
rect 76024 1961 76052 2060
rect 91002 2048 91008 2060
rect 91060 2048 91066 2100
rect 91094 2048 91100 2100
rect 91152 2048 91158 2100
rect 92750 2048 92756 2100
rect 92808 2048 92814 2100
rect 93670 2048 93676 2100
rect 93728 2088 93734 2100
rect 94501 2091 94559 2097
rect 94501 2088 94513 2091
rect 93728 2060 94513 2088
rect 93728 2048 93734 2060
rect 94501 2057 94513 2060
rect 94547 2057 94559 2091
rect 94501 2051 94559 2057
rect 95418 2048 95424 2100
rect 95476 2048 95482 2100
rect 96246 2048 96252 2100
rect 96304 2048 96310 2100
rect 96338 2048 96344 2100
rect 96396 2088 96402 2100
rect 98638 2088 98644 2100
rect 96396 2060 98644 2088
rect 96396 2048 96402 2060
rect 98638 2048 98644 2060
rect 98696 2048 98702 2100
rect 100662 2048 100668 2100
rect 100720 2048 100726 2100
rect 100754 2048 100760 2100
rect 100812 2088 100818 2100
rect 102045 2091 102103 2097
rect 102045 2088 102057 2091
rect 100812 2060 102057 2088
rect 100812 2048 100818 2060
rect 102045 2057 102057 2060
rect 102091 2057 102103 2091
rect 102045 2051 102103 2057
rect 106550 2048 106556 2100
rect 106608 2088 106614 2100
rect 112073 2091 112131 2097
rect 112073 2088 112085 2091
rect 106608 2060 112085 2088
rect 106608 2048 106614 2060
rect 112073 2057 112085 2060
rect 112119 2057 112131 2091
rect 112073 2051 112131 2057
rect 116394 2048 116400 2100
rect 116452 2088 116458 2100
rect 117225 2091 117283 2097
rect 117225 2088 117237 2091
rect 116452 2060 117237 2088
rect 116452 2048 116458 2060
rect 117225 2057 117237 2060
rect 117271 2057 117283 2091
rect 117225 2051 117283 2057
rect 122006 2048 122012 2100
rect 122064 2048 122070 2100
rect 124490 2048 124496 2100
rect 124548 2048 124554 2100
rect 126238 2048 126244 2100
rect 126296 2048 126302 2100
rect 127894 2048 127900 2100
rect 127952 2048 127958 2100
rect 129642 2048 129648 2100
rect 129700 2048 129706 2100
rect 131666 2048 131672 2100
rect 131724 2048 131730 2100
rect 149885 2091 149943 2097
rect 132466 2060 147674 2088
rect 99374 2020 99380 2032
rect 77496 1992 99380 2020
rect 77496 1961 77524 1992
rect 99374 1980 99380 1992
rect 99432 1980 99438 2032
rect 99469 2023 99527 2029
rect 99469 1989 99481 2023
rect 99515 2020 99527 2023
rect 100202 2020 100208 2032
rect 99515 1992 100208 2020
rect 99515 1989 99527 1992
rect 99469 1983 99527 1989
rect 100202 1980 100208 1992
rect 100260 1980 100266 2032
rect 100680 2020 100708 2048
rect 121178 2020 121184 2032
rect 100680 1992 103836 2020
rect 76009 1955 76067 1961
rect 76009 1921 76021 1955
rect 76055 1921 76067 1955
rect 76009 1915 76067 1921
rect 77481 1955 77539 1961
rect 77481 1921 77493 1955
rect 77527 1921 77539 1955
rect 77481 1915 77539 1921
rect 80146 1912 80152 1964
rect 80204 1912 80210 1964
rect 82449 1955 82507 1961
rect 82449 1921 82461 1955
rect 82495 1952 82507 1955
rect 83734 1952 83740 1964
rect 82495 1924 83740 1952
rect 82495 1921 82507 1924
rect 82449 1915 82507 1921
rect 83734 1912 83740 1924
rect 83792 1912 83798 1964
rect 86402 1912 86408 1964
rect 86460 1912 86466 1964
rect 87785 1955 87843 1961
rect 87785 1921 87797 1955
rect 87831 1952 87843 1955
rect 88058 1952 88064 1964
rect 87831 1924 88064 1952
rect 87831 1921 87843 1924
rect 87785 1915 87843 1921
rect 88058 1912 88064 1924
rect 88116 1912 88122 1964
rect 88245 1955 88303 1961
rect 88245 1921 88257 1955
rect 88291 1921 88303 1955
rect 88245 1915 88303 1921
rect 88429 1955 88487 1961
rect 88429 1921 88441 1955
rect 88475 1952 88487 1955
rect 89162 1952 89168 1964
rect 88475 1924 89168 1952
rect 88475 1921 88487 1924
rect 88429 1915 88487 1921
rect 66732 1884 66760 1912
rect 65076 1856 66760 1884
rect 70578 1844 70584 1896
rect 70636 1844 70642 1896
rect 72050 1844 72056 1896
rect 72108 1844 72114 1896
rect 74258 1844 74264 1896
rect 74316 1844 74322 1896
rect 74537 1887 74595 1893
rect 74537 1853 74549 1887
rect 74583 1853 74595 1887
rect 74537 1847 74595 1853
rect 7745 1819 7803 1825
rect 7745 1785 7757 1819
rect 7791 1816 7803 1819
rect 7791 1788 22094 1816
rect 7791 1785 7803 1788
rect 7745 1779 7803 1785
rect 22066 1748 22094 1788
rect 22186 1776 22192 1828
rect 22244 1816 22250 1828
rect 25409 1819 25467 1825
rect 25409 1816 25421 1819
rect 22244 1788 25421 1816
rect 22244 1776 22250 1788
rect 25409 1785 25421 1788
rect 25455 1785 25467 1819
rect 25409 1779 25467 1785
rect 37826 1776 37832 1828
rect 37884 1816 37890 1828
rect 37921 1819 37979 1825
rect 37921 1816 37933 1819
rect 37884 1788 37933 1816
rect 37884 1776 37890 1788
rect 37921 1785 37933 1788
rect 37967 1785 37979 1819
rect 37921 1779 37979 1785
rect 40310 1776 40316 1828
rect 40368 1776 40374 1828
rect 44542 1776 44548 1828
rect 44600 1816 44606 1828
rect 45281 1819 45339 1825
rect 45281 1816 45293 1819
rect 44600 1788 45293 1816
rect 44600 1776 44606 1788
rect 45281 1785 45293 1788
rect 45327 1785 45339 1819
rect 45281 1779 45339 1785
rect 50433 1819 50491 1825
rect 50433 1785 50445 1819
rect 50479 1816 50491 1819
rect 50522 1816 50528 1828
rect 50479 1788 50528 1816
rect 50479 1785 50491 1788
rect 50433 1779 50491 1785
rect 50522 1776 50528 1788
rect 50580 1776 50586 1828
rect 53101 1819 53159 1825
rect 53101 1785 53113 1819
rect 53147 1816 53159 1819
rect 53926 1816 53932 1828
rect 53147 1788 53932 1816
rect 53147 1785 53159 1788
rect 53101 1779 53159 1785
rect 53926 1776 53932 1788
rect 53984 1776 53990 1828
rect 74552 1816 74580 1847
rect 75730 1844 75736 1896
rect 75788 1844 75794 1896
rect 77202 1844 77208 1896
rect 77260 1844 77266 1896
rect 79873 1887 79931 1893
rect 79873 1853 79885 1887
rect 79919 1884 79931 1887
rect 80054 1884 80060 1896
rect 79919 1856 80060 1884
rect 79919 1853 79931 1856
rect 79873 1847 79931 1853
rect 80054 1844 80060 1856
rect 80112 1844 80118 1896
rect 81161 1887 81219 1893
rect 81161 1853 81173 1887
rect 81207 1884 81219 1887
rect 81342 1884 81348 1896
rect 81207 1856 81348 1884
rect 81207 1853 81219 1856
rect 81161 1847 81219 1853
rect 81342 1844 81348 1856
rect 81400 1844 81406 1896
rect 81434 1844 81440 1896
rect 81492 1844 81498 1896
rect 82630 1844 82636 1896
rect 82688 1884 82694 1896
rect 82725 1887 82783 1893
rect 82725 1884 82737 1887
rect 82688 1856 82737 1884
rect 82688 1844 82694 1856
rect 82725 1853 82737 1856
rect 82771 1853 82783 1887
rect 82725 1847 82783 1853
rect 83826 1844 83832 1896
rect 83884 1844 83890 1896
rect 84010 1844 84016 1896
rect 84068 1844 84074 1896
rect 85669 1887 85727 1893
rect 85669 1853 85681 1887
rect 85715 1884 85727 1887
rect 86034 1884 86040 1896
rect 85715 1856 86040 1884
rect 85715 1853 85727 1856
rect 85669 1847 85727 1853
rect 86034 1844 86040 1856
rect 86092 1844 86098 1896
rect 86126 1844 86132 1896
rect 86184 1844 86190 1896
rect 88260 1884 88288 1915
rect 89162 1912 89168 1924
rect 89220 1912 89226 1964
rect 89257 1955 89315 1961
rect 89257 1921 89269 1955
rect 89303 1921 89315 1955
rect 89257 1915 89315 1921
rect 89441 1955 89499 1961
rect 89441 1921 89453 1955
rect 89487 1952 89499 1955
rect 89898 1952 89904 1964
rect 89487 1924 89904 1952
rect 89487 1921 89499 1924
rect 89441 1915 89499 1921
rect 88518 1884 88524 1896
rect 88260 1856 88524 1884
rect 88518 1844 88524 1856
rect 88576 1844 88582 1896
rect 89070 1844 89076 1896
rect 89128 1844 89134 1896
rect 89272 1884 89300 1915
rect 89898 1912 89904 1924
rect 89956 1912 89962 1964
rect 89990 1912 89996 1964
rect 90048 1912 90054 1964
rect 90085 1955 90143 1961
rect 90085 1921 90097 1955
rect 90131 1921 90143 1955
rect 90085 1915 90143 1921
rect 89530 1884 89536 1896
rect 89272 1856 89536 1884
rect 89530 1844 89536 1856
rect 89588 1884 89594 1896
rect 90100 1884 90128 1915
rect 90726 1912 90732 1964
rect 90784 1912 90790 1964
rect 90913 1955 90971 1961
rect 90913 1921 90925 1955
rect 90959 1952 90971 1955
rect 91741 1955 91799 1961
rect 91741 1952 91753 1955
rect 90959 1924 91753 1952
rect 90959 1921 90971 1924
rect 90913 1915 90971 1921
rect 91741 1921 91753 1924
rect 91787 1952 91799 1955
rect 91787 1924 92244 1952
rect 91787 1921 91799 1924
rect 91741 1915 91799 1921
rect 90928 1884 90956 1915
rect 89588 1856 90956 1884
rect 91557 1887 91615 1893
rect 89588 1844 89594 1856
rect 91557 1853 91569 1887
rect 91603 1884 91615 1887
rect 92014 1884 92020 1896
rect 91603 1856 92020 1884
rect 91603 1853 91615 1856
rect 91557 1847 91615 1853
rect 92014 1844 92020 1856
rect 92072 1844 92078 1896
rect 92216 1884 92244 1924
rect 92290 1912 92296 1964
rect 92348 1952 92354 1964
rect 92385 1955 92443 1961
rect 92385 1952 92397 1955
rect 92348 1924 92397 1952
rect 92348 1912 92354 1924
rect 92385 1921 92397 1924
rect 92431 1921 92443 1955
rect 92385 1915 92443 1921
rect 92569 1955 92627 1961
rect 92569 1921 92581 1955
rect 92615 1921 92627 1955
rect 92569 1915 92627 1921
rect 92584 1884 92612 1915
rect 93302 1912 93308 1964
rect 93360 1912 93366 1964
rect 93397 1955 93455 1961
rect 93397 1921 93409 1955
rect 93443 1921 93455 1955
rect 93397 1915 93455 1921
rect 93412 1884 93440 1915
rect 94130 1912 94136 1964
rect 94188 1912 94194 1964
rect 94317 1955 94375 1961
rect 94317 1921 94329 1955
rect 94363 1921 94375 1955
rect 94317 1915 94375 1921
rect 94332 1884 94360 1915
rect 95142 1912 95148 1964
rect 95200 1912 95206 1964
rect 95237 1955 95295 1961
rect 95237 1921 95249 1955
rect 95283 1952 95295 1955
rect 96065 1955 96123 1961
rect 96065 1952 96077 1955
rect 95283 1924 96077 1952
rect 95283 1921 95295 1924
rect 95237 1915 95295 1921
rect 96065 1921 96077 1924
rect 96111 1952 96123 1955
rect 96893 1955 96951 1961
rect 96893 1952 96905 1955
rect 96111 1924 96905 1952
rect 96111 1921 96123 1924
rect 96065 1915 96123 1921
rect 96893 1921 96905 1924
rect 96939 1952 96951 1955
rect 97721 1955 97779 1961
rect 97721 1952 97733 1955
rect 96939 1924 97733 1952
rect 96939 1921 96951 1924
rect 96893 1915 96951 1921
rect 97721 1921 97733 1924
rect 97767 1952 97779 1955
rect 98546 1952 98552 1964
rect 97767 1924 98552 1952
rect 97767 1921 97779 1924
rect 97721 1915 97779 1921
rect 94958 1884 94964 1896
rect 92216 1856 94964 1884
rect 94958 1844 94964 1856
rect 95016 1884 95022 1896
rect 95252 1884 95280 1915
rect 98546 1912 98552 1924
rect 98604 1912 98610 1964
rect 100110 1952 100116 1964
rect 99760 1924 100116 1952
rect 95016 1856 95280 1884
rect 95881 1887 95939 1893
rect 95016 1844 95022 1856
rect 95881 1853 95893 1887
rect 95927 1853 95939 1887
rect 95881 1847 95939 1853
rect 96709 1887 96767 1893
rect 96709 1853 96721 1887
rect 96755 1853 96767 1887
rect 96709 1847 96767 1853
rect 95234 1816 95240 1828
rect 74552 1788 95240 1816
rect 95234 1776 95240 1788
rect 95292 1776 95298 1828
rect 95896 1816 95924 1847
rect 95970 1816 95976 1828
rect 95896 1788 95976 1816
rect 95970 1776 95976 1788
rect 96028 1776 96034 1828
rect 96724 1816 96752 1847
rect 97534 1844 97540 1896
rect 97592 1844 97598 1896
rect 98362 1844 98368 1896
rect 98420 1844 98426 1896
rect 99760 1893 99788 1924
rect 100110 1912 100116 1924
rect 100168 1952 100174 1964
rect 100481 1955 100539 1961
rect 100481 1952 100493 1955
rect 100168 1924 100493 1952
rect 100168 1912 100174 1924
rect 100481 1921 100493 1924
rect 100527 1921 100539 1955
rect 100481 1915 100539 1921
rect 100665 1955 100723 1961
rect 100665 1921 100677 1955
rect 100711 1952 100723 1955
rect 101125 1955 101183 1961
rect 101125 1952 101137 1955
rect 100711 1924 101137 1952
rect 100711 1921 100723 1924
rect 100665 1915 100723 1921
rect 101125 1921 101137 1924
rect 101171 1921 101183 1955
rect 101861 1955 101919 1961
rect 101861 1952 101873 1955
rect 101125 1915 101183 1921
rect 101232 1924 101873 1952
rect 99745 1887 99803 1893
rect 99745 1853 99757 1887
rect 99791 1853 99803 1887
rect 99745 1847 99803 1853
rect 99834 1844 99840 1896
rect 99892 1884 99898 1896
rect 100297 1887 100355 1893
rect 100297 1884 100309 1887
rect 99892 1856 100309 1884
rect 99892 1844 99898 1856
rect 100297 1853 100309 1856
rect 100343 1853 100355 1887
rect 100297 1847 100355 1853
rect 96798 1816 96804 1828
rect 96724 1788 96804 1816
rect 96798 1776 96804 1788
rect 96856 1776 96862 1828
rect 98733 1819 98791 1825
rect 98733 1785 98745 1819
rect 98779 1816 98791 1819
rect 101232 1816 101260 1924
rect 101861 1921 101873 1924
rect 101907 1921 101919 1955
rect 101861 1915 101919 1921
rect 98779 1788 101260 1816
rect 103808 1816 103836 1992
rect 120920 1992 121184 2020
rect 107102 1912 107108 1964
rect 107160 1912 107166 1964
rect 112254 1912 112260 1964
rect 112312 1912 112318 1964
rect 117314 1912 117320 1964
rect 117372 1952 117378 1964
rect 120920 1961 120948 1992
rect 121178 1980 121184 1992
rect 121236 1980 121242 2032
rect 129182 2020 129188 2032
rect 123496 1992 127756 2020
rect 117409 1955 117467 1961
rect 117409 1952 117421 1955
rect 117372 1924 117421 1952
rect 117372 1912 117378 1924
rect 117409 1921 117421 1924
rect 117455 1921 117467 1955
rect 117409 1915 117467 1921
rect 120905 1955 120963 1961
rect 120905 1921 120917 1955
rect 120951 1921 120963 1955
rect 120905 1915 120963 1921
rect 120997 1955 121055 1961
rect 120997 1921 121009 1955
rect 121043 1952 121055 1955
rect 121825 1955 121883 1961
rect 121825 1952 121837 1955
rect 121043 1924 121837 1952
rect 121043 1921 121055 1924
rect 120997 1915 121055 1921
rect 121825 1921 121837 1924
rect 121871 1952 121883 1955
rect 122653 1955 122711 1961
rect 122653 1952 122665 1955
rect 121871 1924 122665 1952
rect 121871 1921 121883 1924
rect 121825 1915 121883 1921
rect 122653 1921 122665 1924
rect 122699 1952 122711 1955
rect 122834 1952 122840 1964
rect 122699 1924 122840 1952
rect 122699 1921 122711 1924
rect 122653 1915 122711 1921
rect 122834 1912 122840 1924
rect 122892 1952 122898 1964
rect 123496 1961 123524 1992
rect 123481 1955 123539 1961
rect 123481 1952 123493 1955
rect 122892 1924 123493 1952
rect 122892 1912 122898 1924
rect 123481 1921 123493 1924
rect 123527 1921 123539 1955
rect 123481 1915 123539 1921
rect 124122 1912 124128 1964
rect 124180 1912 124186 1964
rect 124324 1961 124352 1992
rect 124309 1955 124367 1961
rect 124309 1921 124321 1955
rect 124355 1921 124367 1955
rect 124309 1915 124367 1921
rect 125042 1912 125048 1964
rect 125100 1912 125106 1964
rect 125244 1961 125272 1992
rect 125229 1955 125287 1961
rect 125229 1921 125241 1955
rect 125275 1921 125287 1955
rect 125229 1915 125287 1921
rect 125962 1912 125968 1964
rect 126020 1912 126026 1964
rect 126072 1961 126100 1992
rect 126057 1955 126115 1961
rect 126057 1921 126069 1955
rect 126103 1921 126115 1955
rect 126057 1915 126115 1921
rect 126698 1912 126704 1964
rect 126756 1912 126762 1964
rect 126900 1961 126928 1992
rect 126885 1955 126943 1961
rect 126885 1921 126897 1955
rect 126931 1921 126943 1955
rect 126885 1915 126943 1921
rect 127618 1912 127624 1964
rect 127676 1912 127682 1964
rect 127728 1961 127756 1992
rect 128556 1992 129188 2020
rect 128556 1961 128584 1992
rect 129182 1980 129188 1992
rect 129240 1980 129246 2032
rect 129550 2020 129556 2032
rect 129384 1992 129556 2020
rect 129384 1961 129412 1992
rect 129550 1980 129556 1992
rect 129608 1980 129614 2032
rect 132466 2020 132494 2060
rect 129660 1992 132494 2020
rect 127713 1955 127771 1961
rect 127713 1921 127725 1955
rect 127759 1921 127771 1955
rect 127713 1915 127771 1921
rect 128541 1955 128599 1961
rect 128541 1921 128553 1955
rect 128587 1921 128599 1955
rect 128541 1915 128599 1921
rect 128633 1955 128691 1961
rect 128633 1921 128645 1955
rect 128679 1921 128691 1955
rect 128633 1915 128691 1921
rect 129369 1955 129427 1961
rect 129369 1921 129381 1955
rect 129415 1921 129427 1955
rect 129369 1915 129427 1921
rect 129461 1955 129519 1961
rect 129461 1921 129473 1955
rect 129507 1921 129519 1955
rect 129461 1915 129519 1921
rect 121638 1844 121644 1896
rect 121696 1844 121702 1896
rect 122466 1844 122472 1896
rect 122524 1844 122530 1896
rect 123294 1844 123300 1896
rect 123352 1844 123358 1896
rect 127728 1884 127756 1915
rect 128446 1884 128452 1896
rect 127728 1856 128452 1884
rect 128446 1844 128452 1856
rect 128504 1884 128510 1896
rect 128648 1884 128676 1915
rect 129476 1884 129504 1915
rect 129550 1884 129556 1896
rect 128504 1856 129556 1884
rect 128504 1844 128510 1856
rect 129550 1844 129556 1856
rect 129608 1844 129614 1896
rect 106921 1819 106979 1825
rect 106921 1816 106933 1819
rect 103808 1788 106933 1816
rect 98779 1785 98791 1788
rect 98733 1779 98791 1785
rect 106921 1785 106933 1788
rect 106967 1785 106979 1819
rect 123312 1816 123340 1844
rect 129660 1816 129688 1992
rect 133598 1980 133604 2032
rect 133656 1980 133662 2032
rect 134978 2020 134984 2032
rect 134168 1992 134984 2020
rect 130562 1912 130568 1964
rect 130620 1912 130626 1964
rect 130657 1955 130715 1961
rect 130657 1921 130669 1955
rect 130703 1921 130715 1955
rect 130657 1915 130715 1921
rect 129734 1844 129740 1896
rect 129792 1884 129798 1896
rect 130672 1884 130700 1915
rect 131114 1912 131120 1964
rect 131172 1952 131178 1964
rect 131301 1955 131359 1961
rect 131301 1952 131313 1955
rect 131172 1924 131313 1952
rect 131172 1912 131178 1924
rect 131301 1921 131313 1924
rect 131347 1921 131359 1955
rect 131301 1915 131359 1921
rect 131485 1955 131543 1961
rect 131485 1921 131497 1955
rect 131531 1921 131543 1955
rect 131485 1915 131543 1921
rect 131500 1884 131528 1915
rect 131850 1912 131856 1964
rect 131908 1952 131914 1964
rect 132221 1955 132279 1961
rect 132221 1952 132233 1955
rect 131908 1924 132233 1952
rect 131908 1912 131914 1924
rect 132221 1921 132233 1924
rect 132267 1921 132279 1955
rect 132221 1915 132279 1921
rect 132405 1955 132463 1961
rect 132405 1921 132417 1955
rect 132451 1952 132463 1955
rect 132451 1924 132485 1952
rect 132451 1921 132463 1924
rect 132405 1915 132463 1921
rect 132420 1884 132448 1915
rect 133046 1912 133052 1964
rect 133104 1952 133110 1964
rect 134168 1961 134196 1992
rect 134978 1980 134984 1992
rect 135036 1980 135042 2032
rect 139946 1980 139952 2032
rect 140004 1980 140010 2032
rect 147646 2020 147674 2060
rect 149885 2057 149897 2091
rect 149931 2088 149943 2091
rect 150802 2088 150808 2100
rect 149931 2060 150808 2088
rect 149931 2057 149943 2060
rect 149885 2051 149943 2057
rect 150802 2048 150808 2060
rect 150860 2048 150866 2100
rect 155313 2091 155371 2097
rect 155313 2057 155325 2091
rect 155359 2088 155371 2091
rect 157886 2088 157892 2100
rect 155359 2060 157892 2088
rect 155359 2057 155371 2060
rect 155313 2051 155371 2057
rect 157886 2048 157892 2060
rect 157944 2048 157950 2100
rect 157978 2048 157984 2100
rect 158036 2088 158042 2100
rect 162118 2088 162124 2100
rect 158036 2060 162124 2088
rect 158036 2048 158042 2060
rect 162118 2048 162124 2060
rect 162176 2048 162182 2100
rect 162302 2048 162308 2100
rect 162360 2048 162366 2100
rect 163958 2048 163964 2100
rect 164016 2048 164022 2100
rect 165614 2048 165620 2100
rect 165672 2048 165678 2100
rect 165890 2048 165896 2100
rect 165948 2088 165954 2100
rect 166629 2091 166687 2097
rect 166629 2088 166641 2091
rect 165948 2060 166641 2088
rect 165948 2048 165954 2060
rect 166629 2057 166641 2060
rect 166675 2057 166687 2091
rect 166629 2051 166687 2057
rect 167454 2048 167460 2100
rect 167512 2048 167518 2100
rect 167546 2048 167552 2100
rect 167604 2088 167610 2100
rect 167604 2060 187188 2088
rect 167604 2048 167610 2060
rect 157150 2020 157156 2032
rect 147646 1992 157156 2020
rect 157150 1980 157156 1992
rect 157208 1980 157214 2032
rect 157260 1992 179460 2020
rect 133233 1955 133291 1961
rect 133233 1952 133245 1955
rect 133104 1924 133245 1952
rect 133104 1912 133110 1924
rect 133233 1921 133245 1924
rect 133279 1921 133291 1955
rect 133233 1915 133291 1921
rect 133417 1955 133475 1961
rect 133417 1921 133429 1955
rect 133463 1921 133475 1955
rect 133417 1915 133475 1921
rect 134153 1955 134211 1961
rect 134153 1921 134165 1955
rect 134199 1921 134211 1955
rect 134153 1915 134211 1921
rect 134245 1955 134303 1961
rect 134245 1921 134257 1955
rect 134291 1952 134303 1955
rect 134429 1955 134487 1961
rect 134291 1924 134380 1952
rect 134291 1921 134303 1924
rect 134245 1915 134303 1921
rect 133138 1884 133144 1896
rect 129792 1856 133144 1884
rect 129792 1844 129798 1856
rect 133138 1844 133144 1856
rect 133196 1884 133202 1896
rect 133432 1884 133460 1915
rect 134058 1884 134064 1896
rect 133196 1856 134064 1884
rect 133196 1844 133202 1856
rect 134058 1844 134064 1856
rect 134116 1884 134122 1896
rect 134352 1884 134380 1924
rect 134429 1921 134441 1955
rect 134475 1952 134487 1955
rect 135349 1955 135407 1961
rect 135349 1952 135361 1955
rect 134475 1924 135361 1952
rect 134475 1921 134487 1924
rect 134429 1915 134487 1921
rect 135349 1921 135361 1924
rect 135395 1921 135407 1955
rect 135349 1915 135407 1921
rect 138106 1912 138112 1964
rect 138164 1912 138170 1964
rect 139026 1912 139032 1964
rect 139084 1912 139090 1964
rect 139210 1961 139216 1964
rect 139167 1955 139216 1961
rect 139167 1921 139179 1955
rect 139213 1921 139216 1955
rect 139167 1915 139216 1921
rect 139210 1912 139216 1915
rect 139268 1912 139274 1964
rect 140406 1912 140412 1964
rect 140464 1952 140470 1964
rect 140501 1955 140559 1961
rect 140501 1952 140513 1955
rect 140464 1924 140513 1952
rect 140464 1912 140470 1924
rect 140501 1921 140513 1924
rect 140547 1921 140559 1955
rect 140501 1915 140559 1921
rect 141418 1912 141424 1964
rect 141476 1912 141482 1964
rect 141694 1912 141700 1964
rect 141752 1912 141758 1964
rect 142982 1912 142988 1964
rect 143040 1912 143046 1964
rect 144914 1912 144920 1964
rect 144972 1912 144978 1964
rect 150066 1912 150072 1964
rect 150124 1912 150130 1964
rect 155129 1955 155187 1961
rect 155129 1921 155141 1955
rect 155175 1921 155187 1955
rect 155129 1915 155187 1921
rect 155957 1955 156015 1961
rect 155957 1921 155969 1955
rect 156003 1952 156015 1955
rect 156690 1952 156696 1964
rect 156003 1924 156696 1952
rect 156003 1921 156015 1924
rect 155957 1915 156015 1921
rect 134116 1856 134380 1884
rect 134116 1844 134122 1856
rect 138290 1844 138296 1896
rect 138348 1844 138354 1896
rect 138382 1844 138388 1896
rect 138440 1884 138446 1896
rect 138753 1887 138811 1893
rect 138753 1884 138765 1887
rect 138440 1856 138765 1884
rect 138440 1844 138446 1856
rect 138753 1853 138765 1856
rect 138799 1853 138811 1887
rect 138753 1847 138811 1853
rect 123312 1788 129688 1816
rect 106921 1779 106979 1785
rect 23658 1748 23664 1760
rect 22066 1720 23664 1748
rect 23658 1708 23664 1720
rect 23716 1708 23722 1760
rect 23750 1708 23756 1760
rect 23808 1748 23814 1760
rect 24673 1751 24731 1757
rect 24673 1748 24685 1751
rect 23808 1720 24685 1748
rect 23808 1708 23814 1720
rect 24673 1717 24685 1720
rect 24719 1717 24731 1751
rect 24673 1711 24731 1717
rect 24854 1708 24860 1760
rect 24912 1748 24918 1760
rect 27341 1751 27399 1757
rect 27341 1748 27353 1751
rect 24912 1720 27353 1748
rect 24912 1708 24918 1720
rect 27341 1717 27353 1720
rect 27387 1717 27399 1751
rect 27341 1711 27399 1717
rect 28902 1708 28908 1760
rect 28960 1748 28966 1760
rect 28997 1751 29055 1757
rect 28997 1748 29009 1751
rect 28960 1720 29009 1748
rect 28960 1708 28966 1720
rect 28997 1717 29009 1720
rect 29043 1717 29055 1751
rect 28997 1711 29055 1717
rect 29730 1708 29736 1760
rect 29788 1748 29794 1760
rect 29825 1751 29883 1757
rect 29825 1748 29837 1751
rect 29788 1720 29837 1748
rect 29788 1708 29794 1720
rect 29825 1717 29837 1720
rect 29871 1717 29883 1751
rect 29825 1711 29883 1717
rect 30558 1708 30564 1760
rect 30616 1748 30622 1760
rect 30745 1751 30803 1757
rect 30745 1748 30757 1751
rect 30616 1720 30757 1748
rect 30616 1708 30622 1720
rect 30745 1717 30757 1720
rect 30791 1717 30803 1751
rect 30745 1711 30803 1717
rect 31754 1708 31760 1760
rect 31812 1708 31818 1760
rect 33134 1708 33140 1760
rect 33192 1748 33198 1760
rect 33321 1751 33379 1757
rect 33321 1748 33333 1751
rect 33192 1720 33333 1748
rect 33192 1708 33198 1720
rect 33321 1717 33333 1720
rect 33367 1717 33379 1751
rect 33321 1711 33379 1717
rect 36814 1708 36820 1760
rect 36872 1708 36878 1760
rect 53466 1708 53472 1760
rect 53524 1708 53530 1760
rect 55861 1751 55919 1757
rect 55861 1717 55873 1751
rect 55907 1748 55919 1751
rect 56042 1748 56048 1760
rect 55907 1720 56048 1748
rect 55907 1717 55919 1720
rect 55861 1711 55919 1717
rect 56042 1708 56048 1720
rect 56100 1708 56106 1760
rect 56689 1751 56747 1757
rect 56689 1717 56701 1751
rect 56735 1748 56747 1751
rect 56870 1748 56876 1760
rect 56735 1720 56876 1748
rect 56735 1717 56747 1720
rect 56689 1711 56747 1717
rect 56870 1708 56876 1720
rect 56928 1708 56934 1760
rect 58253 1751 58311 1757
rect 58253 1717 58265 1751
rect 58299 1748 58311 1751
rect 58434 1748 58440 1760
rect 58299 1720 58440 1748
rect 58299 1717 58311 1720
rect 58253 1711 58311 1717
rect 58434 1708 58440 1720
rect 58492 1708 58498 1760
rect 60185 1751 60243 1757
rect 60185 1717 60197 1751
rect 60231 1748 60243 1751
rect 60642 1748 60648 1760
rect 60231 1720 60648 1748
rect 60231 1717 60243 1720
rect 60185 1711 60243 1717
rect 60642 1708 60648 1720
rect 60700 1708 60706 1760
rect 61013 1751 61071 1757
rect 61013 1717 61025 1751
rect 61059 1748 61071 1751
rect 61378 1748 61384 1760
rect 61059 1720 61384 1748
rect 61059 1717 61071 1720
rect 61013 1711 61071 1717
rect 61378 1708 61384 1720
rect 61436 1708 61442 1760
rect 61838 1708 61844 1760
rect 61896 1708 61902 1760
rect 63586 1708 63592 1760
rect 63644 1708 63650 1760
rect 64322 1708 64328 1760
rect 64380 1748 64386 1760
rect 64417 1751 64475 1757
rect 64417 1748 64429 1751
rect 64380 1720 64429 1748
rect 64380 1708 64386 1720
rect 64417 1717 64429 1720
rect 64463 1717 64475 1751
rect 64417 1711 64475 1717
rect 65978 1708 65984 1760
rect 66036 1748 66042 1760
rect 66073 1751 66131 1757
rect 66073 1748 66085 1751
rect 66036 1720 66085 1748
rect 66036 1708 66042 1720
rect 66073 1717 66085 1720
rect 66119 1717 66131 1751
rect 66073 1711 66131 1717
rect 67542 1708 67548 1760
rect 67600 1708 67606 1760
rect 86034 1708 86040 1760
rect 86092 1708 86098 1760
rect 90269 1751 90327 1757
rect 90269 1717 90281 1751
rect 90315 1748 90327 1751
rect 90450 1748 90456 1760
rect 90315 1720 90456 1748
rect 90315 1717 90327 1720
rect 90269 1711 90327 1717
rect 90450 1708 90456 1720
rect 90508 1708 90514 1760
rect 91925 1751 91983 1757
rect 91925 1717 91937 1751
rect 91971 1748 91983 1751
rect 92014 1748 92020 1760
rect 91971 1720 92020 1748
rect 91971 1717 91983 1720
rect 91925 1711 91983 1717
rect 92014 1708 92020 1720
rect 92072 1708 92078 1760
rect 93302 1708 93308 1760
rect 93360 1748 93366 1760
rect 93581 1751 93639 1757
rect 93581 1748 93593 1751
rect 93360 1720 93593 1748
rect 93360 1708 93366 1720
rect 93581 1717 93593 1720
rect 93627 1717 93639 1751
rect 93581 1711 93639 1717
rect 96614 1708 96620 1760
rect 96672 1748 96678 1760
rect 97077 1751 97135 1757
rect 97077 1748 97089 1751
rect 96672 1720 97089 1748
rect 96672 1708 96678 1720
rect 97077 1717 97089 1720
rect 97123 1717 97135 1751
rect 97077 1711 97135 1717
rect 97166 1708 97172 1760
rect 97224 1748 97230 1760
rect 97905 1751 97963 1757
rect 97905 1748 97917 1751
rect 97224 1720 97917 1748
rect 97224 1708 97230 1720
rect 97905 1717 97917 1720
rect 97951 1717 97963 1751
rect 97905 1711 97963 1717
rect 98546 1708 98552 1760
rect 98604 1748 98610 1760
rect 100110 1748 100116 1760
rect 98604 1720 100116 1748
rect 98604 1708 98610 1720
rect 100110 1708 100116 1720
rect 100168 1708 100174 1760
rect 101306 1708 101312 1760
rect 101364 1708 101370 1760
rect 121178 1708 121184 1760
rect 121236 1708 121242 1760
rect 122837 1751 122895 1757
rect 122837 1717 122849 1751
rect 122883 1748 122895 1751
rect 122926 1748 122932 1760
rect 122883 1720 122932 1748
rect 122883 1717 122895 1720
rect 122837 1711 122895 1717
rect 122926 1708 122932 1720
rect 122984 1708 122990 1760
rect 123665 1751 123723 1757
rect 123665 1717 123677 1751
rect 123711 1748 123723 1751
rect 123754 1748 123760 1760
rect 123711 1720 123760 1748
rect 123711 1717 123723 1720
rect 123665 1711 123723 1717
rect 123754 1708 123760 1720
rect 123812 1708 123818 1760
rect 125410 1708 125416 1760
rect 125468 1708 125474 1760
rect 127066 1708 127072 1760
rect 127124 1708 127130 1760
rect 128817 1751 128875 1757
rect 128817 1717 128829 1751
rect 128863 1748 128875 1751
rect 129090 1748 129096 1760
rect 128863 1720 129096 1748
rect 128863 1717 128875 1720
rect 128817 1711 128875 1717
rect 129090 1708 129096 1720
rect 129148 1708 129154 1760
rect 130654 1708 130660 1760
rect 130712 1748 130718 1760
rect 130841 1751 130899 1757
rect 130841 1748 130853 1751
rect 130712 1720 130853 1748
rect 130712 1708 130718 1720
rect 130841 1717 130853 1720
rect 130887 1717 130899 1751
rect 130841 1711 130899 1717
rect 132586 1708 132592 1760
rect 132644 1708 132650 1760
rect 135254 1708 135260 1760
rect 135312 1748 135318 1760
rect 135533 1751 135591 1757
rect 135533 1748 135545 1751
rect 135312 1720 135545 1748
rect 135312 1708 135318 1720
rect 135533 1717 135545 1720
rect 135579 1717 135591 1751
rect 138768 1748 138796 1847
rect 138842 1844 138848 1896
rect 138900 1884 138906 1896
rect 139305 1887 139363 1893
rect 139305 1884 139317 1887
rect 138900 1856 139317 1884
rect 138900 1844 138906 1856
rect 139305 1853 139317 1856
rect 139351 1853 139363 1887
rect 139305 1847 139363 1853
rect 140682 1844 140688 1896
rect 140740 1844 140746 1896
rect 141510 1844 141516 1896
rect 141568 1893 141574 1896
rect 141568 1887 141596 1893
rect 141584 1853 141596 1887
rect 141568 1847 141596 1853
rect 141568 1844 141574 1847
rect 143166 1844 143172 1896
rect 143224 1884 143230 1896
rect 155034 1884 155040 1896
rect 143224 1856 155040 1884
rect 143224 1844 143230 1856
rect 155034 1844 155040 1856
rect 155092 1844 155098 1896
rect 155144 1884 155172 1915
rect 156690 1912 156696 1924
rect 156748 1912 156754 1964
rect 156782 1912 156788 1964
rect 156840 1912 156846 1964
rect 157260 1952 157288 1992
rect 156892 1924 157288 1952
rect 155144 1856 156368 1884
rect 141142 1816 141148 1828
rect 140700 1788 141148 1816
rect 140700 1748 140728 1788
rect 141142 1776 141148 1788
rect 141200 1776 141206 1828
rect 142798 1776 142804 1828
rect 142856 1776 142862 1828
rect 144733 1819 144791 1825
rect 144733 1785 144745 1819
rect 144779 1816 144791 1819
rect 148134 1816 148140 1828
rect 144779 1788 148140 1816
rect 144779 1785 144791 1788
rect 144733 1779 144791 1785
rect 148134 1776 148140 1788
rect 148192 1776 148198 1828
rect 155770 1816 155776 1828
rect 152476 1788 155776 1816
rect 138768 1720 140728 1748
rect 135533 1711 135591 1717
rect 140774 1708 140780 1760
rect 140832 1748 140838 1760
rect 142341 1751 142399 1757
rect 142341 1748 142353 1751
rect 140832 1720 142353 1748
rect 140832 1708 140838 1720
rect 142341 1717 142353 1720
rect 142387 1717 142399 1751
rect 142341 1711 142399 1717
rect 146478 1708 146484 1760
rect 146536 1748 146542 1760
rect 152476 1748 152504 1788
rect 155770 1776 155776 1788
rect 155828 1776 155834 1828
rect 146536 1720 152504 1748
rect 146536 1708 146542 1720
rect 155954 1708 155960 1760
rect 156012 1748 156018 1760
rect 156141 1751 156199 1757
rect 156141 1748 156153 1751
rect 156012 1720 156153 1748
rect 156012 1708 156018 1720
rect 156141 1717 156153 1720
rect 156187 1717 156199 1751
rect 156340 1748 156368 1856
rect 156506 1844 156512 1896
rect 156564 1884 156570 1896
rect 156892 1884 156920 1924
rect 157978 1912 157984 1964
rect 158036 1912 158042 1964
rect 159266 1912 159272 1964
rect 159324 1952 159330 1964
rect 159324 1924 159588 1952
rect 159324 1912 159330 1924
rect 156564 1856 156920 1884
rect 156564 1844 156570 1856
rect 157058 1844 157064 1896
rect 157116 1844 157122 1896
rect 158162 1844 158168 1896
rect 158220 1884 158226 1896
rect 158257 1887 158315 1893
rect 158257 1884 158269 1887
rect 158220 1856 158269 1884
rect 158220 1844 158226 1856
rect 158257 1853 158269 1856
rect 158303 1853 158315 1887
rect 158257 1847 158315 1853
rect 158530 1844 158536 1896
rect 158588 1884 158594 1896
rect 159085 1887 159143 1893
rect 159085 1884 159097 1887
rect 158588 1856 159097 1884
rect 158588 1844 158594 1856
rect 159085 1853 159097 1856
rect 159131 1853 159143 1887
rect 159560 1884 159588 1924
rect 159634 1912 159640 1964
rect 159692 1952 159698 1964
rect 159913 1955 159971 1961
rect 159913 1952 159925 1955
rect 159692 1924 159925 1952
rect 159692 1912 159698 1924
rect 159913 1921 159925 1924
rect 159959 1921 159971 1955
rect 159913 1915 159971 1921
rect 160097 1955 160155 1961
rect 160097 1921 160109 1955
rect 160143 1921 160155 1955
rect 160097 1915 160155 1921
rect 160002 1884 160008 1896
rect 159560 1856 160008 1884
rect 159085 1847 159143 1853
rect 160002 1844 160008 1856
rect 160060 1884 160066 1896
rect 160112 1884 160140 1915
rect 161198 1912 161204 1964
rect 161256 1912 161262 1964
rect 161293 1955 161351 1961
rect 161293 1921 161305 1955
rect 161339 1952 161351 1955
rect 161339 1924 161474 1952
rect 161339 1921 161351 1924
rect 161293 1915 161351 1921
rect 161308 1884 161336 1915
rect 160060 1856 161336 1884
rect 161446 1884 161474 1924
rect 161566 1912 161572 1964
rect 161624 1952 161630 1964
rect 161937 1955 161995 1961
rect 161937 1952 161949 1955
rect 161624 1924 161949 1952
rect 161624 1912 161630 1924
rect 161937 1921 161949 1924
rect 161983 1921 161995 1955
rect 161937 1915 161995 1921
rect 162121 1955 162179 1961
rect 162121 1921 162133 1955
rect 162167 1921 162179 1955
rect 162121 1915 162179 1921
rect 162136 1884 162164 1915
rect 162210 1912 162216 1964
rect 162268 1952 162274 1964
rect 162765 1955 162823 1961
rect 162765 1952 162777 1955
rect 162268 1924 162777 1952
rect 162268 1912 162274 1924
rect 162765 1921 162777 1924
rect 162811 1921 162823 1955
rect 162765 1915 162823 1921
rect 162949 1955 163007 1961
rect 162949 1921 162961 1955
rect 162995 1921 163007 1955
rect 162949 1915 163007 1921
rect 162964 1884 162992 1915
rect 163682 1912 163688 1964
rect 163740 1912 163746 1964
rect 163774 1912 163780 1964
rect 163832 1952 163838 1964
rect 163832 1924 163912 1952
rect 163832 1912 163838 1924
rect 163130 1884 163136 1896
rect 161446 1856 163136 1884
rect 160060 1844 160066 1856
rect 163130 1844 163136 1856
rect 163188 1884 163194 1896
rect 163884 1884 163912 1924
rect 164326 1912 164332 1964
rect 164384 1952 164390 1964
rect 164421 1955 164479 1961
rect 164421 1952 164433 1955
rect 164384 1924 164433 1952
rect 164384 1912 164390 1924
rect 164421 1921 164433 1924
rect 164467 1921 164479 1955
rect 164421 1915 164479 1921
rect 164605 1955 164663 1961
rect 164605 1921 164617 1955
rect 164651 1921 164663 1955
rect 164605 1915 164663 1921
rect 164620 1884 164648 1915
rect 165246 1912 165252 1964
rect 165304 1912 165310 1964
rect 165433 1955 165491 1961
rect 165433 1921 165445 1955
rect 165479 1921 165491 1955
rect 165433 1915 165491 1921
rect 165448 1884 165476 1915
rect 166258 1912 166264 1964
rect 166316 1912 166322 1964
rect 166445 1955 166503 1961
rect 166445 1921 166457 1955
rect 166491 1921 166503 1955
rect 166445 1915 166503 1921
rect 166460 1884 166488 1915
rect 167086 1912 167092 1964
rect 167144 1912 167150 1964
rect 167273 1955 167331 1961
rect 167273 1921 167285 1955
rect 167319 1921 167331 1955
rect 167273 1915 167331 1921
rect 167178 1884 167184 1896
rect 163188 1856 167184 1884
rect 163188 1844 163194 1856
rect 167178 1844 167184 1856
rect 167236 1884 167242 1896
rect 167288 1884 167316 1915
rect 167914 1912 167920 1964
rect 167972 1912 167978 1964
rect 168101 1955 168159 1961
rect 168101 1921 168113 1955
rect 168147 1921 168159 1955
rect 168101 1915 168159 1921
rect 168285 1955 168343 1961
rect 168285 1921 168297 1955
rect 168331 1952 168343 1955
rect 168745 1955 168803 1961
rect 168745 1952 168757 1955
rect 168331 1924 168757 1952
rect 168331 1921 168343 1924
rect 168285 1915 168343 1921
rect 168745 1921 168757 1924
rect 168791 1921 168803 1955
rect 168745 1915 168803 1921
rect 167822 1884 167828 1896
rect 167236 1856 167828 1884
rect 167236 1844 167242 1856
rect 167822 1844 167828 1856
rect 167880 1884 167886 1896
rect 168116 1884 168144 1915
rect 173250 1912 173256 1964
rect 173308 1912 173314 1964
rect 174722 1912 174728 1964
rect 174780 1912 174786 1964
rect 176838 1912 176844 1964
rect 176896 1912 176902 1964
rect 179432 1961 179460 1992
rect 179417 1955 179475 1961
rect 179417 1921 179429 1955
rect 179463 1921 179475 1955
rect 179417 1915 179475 1921
rect 181898 1912 181904 1964
rect 181956 1912 181962 1964
rect 183554 1912 183560 1964
rect 183612 1912 183618 1964
rect 185026 1912 185032 1964
rect 185084 1912 185090 1964
rect 187160 1961 187188 2060
rect 190362 2048 190368 2100
rect 190420 2088 190426 2100
rect 191101 2091 191159 2097
rect 191101 2088 191113 2091
rect 190420 2060 191113 2088
rect 190420 2048 190426 2060
rect 191101 2057 191113 2060
rect 191147 2057 191159 2091
rect 191101 2051 191159 2057
rect 192386 2048 192392 2100
rect 192444 2048 192450 2100
rect 195698 2048 195704 2100
rect 195756 2048 195762 2100
rect 196250 2048 196256 2100
rect 196308 2088 196314 2100
rect 197541 2091 197599 2097
rect 197541 2088 197553 2091
rect 196308 2060 197553 2088
rect 196308 2048 196314 2060
rect 197541 2057 197553 2060
rect 197587 2057 197599 2091
rect 197541 2051 197599 2057
rect 199194 2048 199200 2100
rect 199252 2048 199258 2100
rect 200850 2048 200856 2100
rect 200908 2048 200914 2100
rect 201310 2048 201316 2100
rect 201368 2048 201374 2100
rect 207014 2048 207020 2100
rect 207072 2088 207078 2100
rect 211154 2088 211160 2100
rect 207072 2060 211160 2088
rect 207072 2048 207078 2060
rect 211154 2048 211160 2060
rect 211212 2048 211218 2100
rect 211525 2091 211583 2097
rect 211525 2057 211537 2091
rect 211571 2088 211583 2091
rect 215386 2088 215392 2100
rect 211571 2060 215392 2088
rect 211571 2057 211583 2060
rect 211525 2051 211583 2057
rect 215386 2048 215392 2060
rect 215444 2048 215450 2100
rect 216125 2091 216183 2097
rect 216125 2057 216137 2091
rect 216171 2088 216183 2091
rect 216950 2088 216956 2100
rect 216171 2060 216956 2088
rect 216171 2057 216183 2060
rect 216125 2051 216183 2057
rect 216950 2048 216956 2060
rect 217008 2048 217014 2100
rect 217134 2048 217140 2100
rect 217192 2048 217198 2100
rect 221645 2091 221703 2097
rect 221645 2057 221657 2091
rect 221691 2088 221703 2091
rect 221826 2088 221832 2100
rect 221691 2060 221832 2088
rect 221691 2057 221703 2060
rect 221645 2051 221703 2057
rect 221826 2048 221832 2060
rect 221884 2048 221890 2100
rect 223022 2048 223028 2100
rect 223080 2088 223086 2100
rect 224218 2088 224224 2100
rect 223080 2060 224224 2088
rect 223080 2048 223086 2060
rect 224218 2048 224224 2060
rect 224276 2048 224282 2100
rect 225322 2048 225328 2100
rect 225380 2048 225386 2100
rect 226150 2048 226156 2100
rect 226208 2048 226214 2100
rect 226978 2048 226984 2100
rect 227036 2048 227042 2100
rect 228082 2048 228088 2100
rect 228140 2088 228146 2100
rect 228453 2091 228511 2097
rect 228453 2088 228465 2091
rect 228140 2060 228465 2088
rect 228140 2048 228146 2060
rect 228453 2057 228465 2060
rect 228499 2057 228511 2091
rect 228453 2051 228511 2057
rect 229186 2048 229192 2100
rect 229244 2088 229250 2100
rect 235994 2088 236000 2100
rect 229244 2060 236000 2088
rect 229244 2048 229250 2060
rect 235994 2048 236000 2060
rect 236052 2048 236058 2100
rect 236086 2048 236092 2100
rect 236144 2048 236150 2100
rect 245059 2091 245117 2097
rect 245059 2088 245071 2091
rect 238128 2060 245071 2088
rect 192294 2020 192300 2032
rect 192128 1992 192300 2020
rect 187145 1955 187203 1961
rect 187145 1921 187157 1955
rect 187191 1921 187203 1955
rect 187145 1915 187203 1921
rect 189718 1912 189724 1964
rect 189776 1912 189782 1964
rect 190822 1912 190828 1964
rect 190880 1912 190886 1964
rect 190914 1912 190920 1964
rect 190972 1912 190978 1964
rect 192128 1961 192156 1992
rect 192294 1980 192300 1992
rect 192352 1980 192358 2032
rect 193306 2020 193312 2032
rect 192956 1992 193312 2020
rect 192956 1961 192984 1992
rect 193306 1980 193312 1992
rect 193364 1980 193370 2032
rect 201328 2020 201356 2048
rect 200086 1992 202552 2020
rect 192113 1955 192171 1961
rect 192113 1921 192125 1955
rect 192159 1921 192171 1955
rect 192113 1915 192171 1921
rect 192205 1955 192263 1961
rect 192205 1921 192217 1955
rect 192251 1921 192263 1955
rect 192205 1915 192263 1921
rect 192941 1955 192999 1961
rect 192941 1921 192953 1955
rect 192987 1921 192999 1955
rect 192941 1915 192999 1921
rect 193033 1955 193091 1961
rect 193033 1921 193045 1955
rect 193079 1921 193091 1955
rect 193033 1915 193091 1921
rect 167880 1856 168144 1884
rect 167880 1844 167886 1856
rect 172974 1844 172980 1896
rect 173032 1844 173038 1896
rect 174446 1844 174452 1896
rect 174504 1844 174510 1896
rect 176562 1844 176568 1896
rect 176620 1844 176626 1896
rect 177850 1844 177856 1896
rect 177908 1844 177914 1896
rect 178129 1887 178187 1893
rect 178129 1853 178141 1887
rect 178175 1853 178187 1887
rect 178129 1847 178187 1853
rect 156874 1776 156880 1828
rect 156932 1816 156938 1828
rect 178144 1816 178172 1847
rect 179138 1844 179144 1896
rect 179196 1844 179202 1896
rect 183278 1844 183284 1896
rect 183336 1844 183342 1896
rect 184750 1844 184756 1896
rect 184808 1844 184814 1896
rect 186314 1844 186320 1896
rect 186372 1884 186378 1896
rect 186869 1887 186927 1893
rect 186869 1884 186881 1887
rect 186372 1856 186881 1884
rect 186372 1844 186378 1856
rect 186869 1853 186881 1856
rect 186915 1853 186927 1887
rect 186869 1847 186927 1853
rect 188154 1844 188160 1896
rect 188212 1844 188218 1896
rect 188433 1887 188491 1893
rect 188433 1853 188445 1887
rect 188479 1853 188491 1887
rect 188433 1847 188491 1853
rect 156932 1788 178172 1816
rect 156932 1776 156938 1788
rect 179506 1776 179512 1828
rect 179564 1816 179570 1828
rect 188448 1816 188476 1847
rect 189442 1844 189448 1896
rect 189500 1844 189506 1896
rect 190932 1884 190960 1912
rect 192220 1884 192248 1915
rect 193048 1884 193076 1915
rect 193214 1912 193220 1964
rect 193272 1952 193278 1964
rect 193677 1955 193735 1961
rect 193677 1952 193689 1955
rect 193272 1924 193689 1952
rect 193272 1912 193278 1924
rect 193677 1921 193689 1924
rect 193723 1921 193735 1955
rect 193677 1915 193735 1921
rect 193861 1955 193919 1961
rect 193861 1921 193873 1955
rect 193907 1921 193919 1955
rect 193861 1915 193919 1921
rect 193876 1884 193904 1915
rect 194594 1912 194600 1964
rect 194652 1912 194658 1964
rect 194689 1955 194747 1961
rect 194689 1921 194701 1955
rect 194735 1921 194747 1955
rect 194689 1915 194747 1921
rect 194704 1884 194732 1915
rect 195422 1912 195428 1964
rect 195480 1912 195486 1964
rect 195517 1955 195575 1961
rect 195517 1921 195529 1955
rect 195563 1921 195575 1955
rect 195517 1915 195575 1921
rect 195532 1884 195560 1915
rect 196158 1912 196164 1964
rect 196216 1912 196222 1964
rect 196345 1955 196403 1961
rect 196345 1921 196357 1955
rect 196391 1921 196403 1955
rect 196345 1915 196403 1921
rect 196360 1884 196388 1915
rect 196434 1912 196440 1964
rect 196492 1952 196498 1964
rect 197173 1955 197231 1961
rect 197173 1952 197185 1955
rect 196492 1924 197185 1952
rect 196492 1912 196498 1924
rect 197173 1921 197185 1924
rect 197219 1921 197231 1955
rect 197173 1915 197231 1921
rect 197262 1912 197268 1964
rect 197320 1952 197326 1964
rect 197357 1955 197415 1961
rect 197357 1952 197369 1955
rect 197320 1924 197369 1952
rect 197320 1912 197326 1924
rect 197357 1921 197369 1924
rect 197403 1921 197415 1955
rect 197357 1915 197415 1921
rect 197372 1884 197400 1915
rect 197998 1912 198004 1964
rect 198056 1912 198062 1964
rect 198185 1955 198243 1961
rect 198185 1921 198197 1955
rect 198231 1921 198243 1955
rect 198185 1915 198243 1921
rect 198200 1884 198228 1915
rect 198826 1912 198832 1964
rect 198884 1912 198890 1964
rect 199013 1955 199071 1961
rect 199013 1921 199025 1955
rect 199059 1921 199071 1955
rect 199013 1915 199071 1921
rect 199028 1884 199056 1915
rect 199654 1912 199660 1964
rect 199712 1912 199718 1964
rect 199841 1955 199899 1961
rect 199841 1921 199853 1955
rect 199887 1952 199899 1955
rect 200086 1952 200114 1992
rect 199887 1924 200114 1952
rect 199887 1921 199899 1924
rect 199841 1915 199899 1921
rect 199856 1884 199884 1915
rect 200482 1912 200488 1964
rect 200540 1912 200546 1964
rect 200684 1961 200712 1992
rect 200669 1955 200727 1961
rect 200669 1921 200681 1955
rect 200715 1921 200727 1955
rect 200669 1915 200727 1921
rect 201126 1912 201132 1964
rect 201184 1952 201190 1964
rect 201512 1961 201540 1992
rect 201313 1955 201371 1961
rect 201313 1952 201325 1955
rect 201184 1924 201325 1952
rect 201184 1912 201190 1924
rect 201313 1921 201325 1924
rect 201359 1921 201371 1955
rect 201313 1915 201371 1921
rect 201497 1955 201555 1961
rect 201497 1921 201509 1955
rect 201543 1921 201555 1955
rect 201497 1915 201555 1921
rect 202230 1912 202236 1964
rect 202288 1952 202294 1964
rect 202524 1961 202552 1992
rect 216674 1980 216680 2032
rect 216732 1980 216738 2032
rect 202325 1955 202383 1961
rect 202325 1952 202337 1955
rect 202288 1924 202337 1952
rect 202288 1912 202294 1924
rect 202325 1921 202337 1924
rect 202371 1921 202383 1955
rect 202325 1915 202383 1921
rect 202509 1955 202567 1961
rect 202509 1921 202521 1955
rect 202555 1921 202567 1955
rect 202509 1915 202567 1921
rect 202693 1955 202751 1961
rect 202693 1921 202705 1955
rect 202739 1952 202751 1955
rect 203153 1955 203211 1961
rect 203153 1952 203165 1955
rect 202739 1924 203165 1952
rect 202739 1921 202751 1924
rect 202693 1915 202751 1921
rect 203153 1921 203165 1924
rect 203199 1921 203211 1955
rect 203153 1915 203211 1921
rect 211706 1912 211712 1964
rect 211764 1912 211770 1964
rect 216309 1955 216367 1961
rect 216309 1921 216321 1955
rect 216355 1921 216367 1955
rect 216309 1915 216367 1921
rect 190932 1856 199884 1884
rect 179564 1788 188476 1816
rect 216324 1816 216352 1915
rect 216398 1912 216404 1964
rect 216456 1912 216462 1964
rect 217152 1952 217180 2048
rect 218425 2023 218483 2029
rect 218425 1989 218437 2023
rect 218471 2020 218483 2023
rect 218471 1992 219848 2020
rect 218471 1989 218483 1992
rect 218425 1983 218483 1989
rect 217781 1955 217839 1961
rect 217781 1952 217793 1955
rect 217152 1924 217793 1952
rect 217781 1921 217793 1924
rect 217827 1952 217839 1955
rect 218701 1955 218759 1961
rect 218701 1952 218713 1955
rect 217827 1924 218713 1952
rect 217827 1921 217839 1924
rect 217781 1915 217839 1921
rect 218701 1921 218713 1924
rect 218747 1921 218759 1955
rect 218701 1915 218759 1921
rect 218885 1955 218943 1961
rect 218885 1921 218897 1955
rect 218931 1952 218943 1955
rect 219434 1952 219440 1964
rect 218931 1924 219440 1952
rect 218931 1921 218943 1924
rect 218885 1915 218943 1921
rect 219434 1912 219440 1924
rect 219492 1912 219498 1964
rect 219820 1961 219848 1992
rect 222562 1980 222568 2032
rect 222620 2020 222626 2032
rect 222620 1992 223896 2020
rect 222620 1980 222626 1992
rect 219805 1955 219863 1961
rect 219805 1921 219817 1955
rect 219851 1921 219863 1955
rect 219805 1915 219863 1921
rect 220078 1912 220084 1964
rect 220136 1912 220142 1964
rect 220722 1912 220728 1964
rect 220780 1912 220786 1964
rect 220814 1912 220820 1964
rect 220872 1952 220878 1964
rect 221829 1955 221887 1961
rect 221829 1952 221841 1955
rect 220872 1924 221841 1952
rect 220872 1912 220878 1924
rect 221829 1921 221841 1924
rect 221875 1921 221887 1955
rect 221829 1915 221887 1921
rect 222470 1912 222476 1964
rect 222528 1952 222534 1964
rect 222933 1955 222991 1961
rect 222933 1952 222945 1955
rect 222528 1924 222945 1952
rect 222528 1912 222534 1924
rect 222933 1921 222945 1924
rect 222979 1921 222991 1955
rect 222933 1915 222991 1921
rect 223206 1912 223212 1964
rect 223264 1912 223270 1964
rect 223868 1961 223896 1992
rect 223942 1980 223948 2032
rect 224000 2020 224006 2032
rect 225506 2020 225512 2032
rect 224000 1992 225512 2020
rect 224000 1980 224006 1992
rect 225506 1980 225512 1992
rect 225564 1980 225570 2032
rect 230032 1992 231624 2020
rect 223853 1955 223911 1961
rect 223853 1921 223865 1955
rect 223899 1921 223911 1955
rect 223853 1915 223911 1921
rect 224402 1912 224408 1964
rect 224460 1952 224466 1964
rect 224770 1952 224776 1964
rect 224460 1924 224776 1952
rect 224460 1912 224466 1924
rect 224770 1912 224776 1924
rect 224828 1952 224834 1964
rect 224957 1955 225015 1961
rect 224957 1952 224969 1955
rect 224828 1924 224969 1952
rect 224828 1912 224834 1924
rect 224957 1921 224969 1924
rect 225003 1921 225015 1955
rect 224957 1915 225015 1921
rect 225141 1955 225199 1961
rect 225141 1921 225153 1955
rect 225187 1952 225199 1955
rect 225187 1924 225276 1952
rect 225187 1921 225199 1924
rect 225141 1915 225199 1921
rect 217965 1887 218023 1893
rect 217965 1853 217977 1887
rect 218011 1884 218023 1887
rect 218054 1884 218060 1896
rect 218011 1856 218060 1884
rect 218011 1853 218023 1856
rect 217965 1847 218023 1853
rect 218054 1844 218060 1856
rect 218112 1844 218118 1896
rect 219161 1887 219219 1893
rect 219161 1853 219173 1887
rect 219207 1853 219219 1887
rect 219161 1847 219219 1853
rect 216674 1816 216680 1828
rect 216324 1788 216680 1816
rect 179564 1776 179570 1788
rect 216674 1776 216680 1788
rect 216732 1776 216738 1828
rect 219176 1816 219204 1847
rect 220998 1844 221004 1896
rect 221056 1844 221062 1896
rect 222102 1844 222108 1896
rect 222160 1884 222166 1896
rect 224129 1887 224187 1893
rect 222160 1856 223988 1884
rect 222160 1844 222166 1856
rect 223850 1816 223856 1828
rect 219176 1788 223856 1816
rect 223850 1776 223856 1788
rect 223908 1776 223914 1828
rect 223960 1816 223988 1856
rect 224129 1853 224141 1887
rect 224175 1884 224187 1887
rect 224862 1884 224868 1896
rect 224175 1856 224868 1884
rect 224175 1853 224187 1856
rect 224129 1847 224187 1853
rect 224862 1844 224868 1856
rect 224920 1844 224926 1896
rect 225248 1884 225276 1924
rect 225874 1912 225880 1964
rect 225932 1912 225938 1964
rect 225969 1955 226027 1961
rect 225969 1921 225981 1955
rect 226015 1921 226027 1955
rect 225969 1915 226027 1921
rect 225984 1884 226012 1915
rect 226702 1912 226708 1964
rect 226760 1912 226766 1964
rect 226800 1955 226858 1961
rect 226800 1921 226812 1955
rect 226846 1952 226858 1955
rect 226846 1924 226932 1952
rect 226846 1921 226858 1924
rect 226800 1915 226858 1921
rect 226610 1884 226616 1896
rect 224972 1856 225184 1884
rect 225248 1856 226616 1884
rect 224972 1816 225000 1856
rect 223960 1788 225000 1816
rect 225156 1816 225184 1856
rect 226610 1844 226616 1856
rect 226668 1884 226674 1896
rect 226904 1884 226932 1924
rect 227714 1912 227720 1964
rect 227772 1952 227778 1964
rect 228085 1955 228143 1961
rect 228085 1952 228097 1955
rect 227772 1924 228097 1952
rect 227772 1912 227778 1924
rect 228085 1921 228097 1924
rect 228131 1921 228143 1955
rect 228085 1915 228143 1921
rect 228269 1955 228327 1961
rect 228269 1921 228281 1955
rect 228315 1921 228327 1955
rect 228269 1915 228327 1921
rect 228284 1884 228312 1915
rect 228910 1912 228916 1964
rect 228968 1912 228974 1964
rect 229097 1955 229155 1961
rect 229097 1921 229109 1955
rect 229143 1952 229155 1955
rect 229462 1952 229468 1964
rect 229143 1924 229468 1952
rect 229143 1921 229155 1924
rect 229097 1915 229155 1921
rect 228358 1884 228364 1896
rect 226668 1856 228364 1884
rect 226668 1844 226674 1856
rect 228358 1844 228364 1856
rect 228416 1884 228422 1896
rect 229112 1884 229140 1915
rect 229462 1912 229468 1924
rect 229520 1912 229526 1964
rect 229738 1912 229744 1964
rect 229796 1912 229802 1964
rect 229922 1912 229928 1964
rect 229980 1961 229986 1964
rect 229980 1955 230003 1961
rect 229991 1952 230003 1955
rect 230032 1952 230060 1992
rect 230768 1964 230796 1992
rect 231596 1964 231624 1992
rect 231762 1980 231768 2032
rect 231820 1980 231826 2032
rect 231854 1980 231860 2032
rect 231912 2020 231918 2032
rect 232593 2023 232651 2029
rect 232593 2020 232605 2023
rect 231912 1992 232605 2020
rect 231912 1980 231918 1992
rect 232593 1989 232605 1992
rect 232639 1989 232651 2023
rect 233694 2020 233700 2032
rect 232593 1983 232651 1989
rect 233344 1992 233700 2020
rect 229991 1924 230060 1952
rect 229991 1921 230003 1924
rect 229980 1915 230003 1921
rect 229980 1912 229986 1915
rect 230106 1912 230112 1964
rect 230164 1952 230170 1964
rect 230569 1955 230627 1961
rect 230569 1952 230581 1955
rect 230164 1924 230581 1952
rect 230164 1912 230170 1924
rect 230569 1921 230581 1924
rect 230615 1921 230627 1955
rect 230569 1915 230627 1921
rect 230750 1912 230756 1964
rect 230808 1912 230814 1964
rect 231486 1912 231492 1964
rect 231544 1912 231550 1964
rect 231578 1912 231584 1964
rect 231636 1912 231642 1964
rect 232130 1912 232136 1964
rect 232188 1952 232194 1964
rect 232225 1955 232283 1961
rect 232225 1952 232237 1955
rect 232188 1924 232237 1952
rect 232188 1912 232194 1924
rect 232225 1921 232237 1924
rect 232271 1921 232283 1955
rect 232225 1915 232283 1921
rect 232314 1912 232320 1964
rect 232372 1952 232378 1964
rect 232409 1955 232467 1961
rect 232409 1952 232421 1955
rect 232372 1924 232421 1952
rect 232372 1912 232378 1924
rect 232409 1921 232421 1924
rect 232455 1952 232467 1955
rect 233234 1952 233240 1964
rect 232455 1924 233240 1952
rect 232455 1921 232467 1924
rect 232409 1915 232467 1921
rect 233234 1912 233240 1924
rect 233292 1912 233298 1964
rect 233344 1961 233372 1992
rect 233694 1980 233700 1992
rect 233752 1980 233758 2032
rect 233878 1980 233884 2032
rect 233936 2020 233942 2032
rect 238128 2020 238156 2060
rect 245059 2057 245071 2060
rect 245105 2057 245117 2091
rect 245059 2051 245117 2057
rect 251450 2048 251456 2100
rect 251508 2048 251514 2100
rect 257614 2048 257620 2100
rect 257672 2088 257678 2100
rect 257985 2091 258043 2097
rect 257985 2088 257997 2091
rect 257672 2060 257997 2088
rect 257672 2048 257678 2060
rect 257985 2057 257997 2060
rect 258031 2088 258043 2091
rect 258902 2088 258908 2100
rect 258031 2060 258908 2088
rect 258031 2057 258043 2060
rect 257985 2051 258043 2057
rect 258902 2048 258908 2060
rect 258960 2048 258966 2100
rect 258994 2048 259000 2100
rect 259052 2088 259058 2100
rect 259365 2091 259423 2097
rect 259365 2088 259377 2091
rect 259052 2060 259377 2088
rect 259052 2048 259058 2060
rect 259365 2057 259377 2060
rect 259411 2057 259423 2091
rect 259365 2051 259423 2057
rect 259564 2060 260052 2088
rect 233936 1992 238156 2020
rect 238220 1992 241652 2020
rect 233936 1980 233942 1992
rect 233329 1955 233387 1961
rect 233329 1921 233341 1955
rect 233375 1921 233387 1955
rect 233329 1915 233387 1921
rect 233418 1912 233424 1964
rect 233476 1952 233482 1964
rect 234249 1955 234307 1961
rect 234249 1952 234261 1955
rect 233476 1924 234261 1952
rect 233476 1912 233482 1924
rect 234249 1921 234261 1924
rect 234295 1921 234307 1955
rect 234249 1915 234307 1921
rect 228416 1856 229140 1884
rect 228416 1844 228422 1856
rect 229830 1844 229836 1896
rect 229888 1884 229894 1896
rect 229888 1856 234016 1884
rect 229888 1844 229894 1856
rect 233988 1816 234016 1856
rect 234062 1844 234068 1896
rect 234120 1844 234126 1896
rect 234264 1884 234292 1915
rect 234890 1912 234896 1964
rect 234948 1912 234954 1964
rect 235077 1955 235135 1961
rect 235077 1921 235089 1955
rect 235123 1952 235135 1955
rect 235905 1955 235963 1961
rect 235905 1952 235917 1955
rect 235123 1924 235917 1952
rect 235123 1921 235135 1924
rect 235077 1915 235135 1921
rect 235905 1921 235917 1924
rect 235951 1952 235963 1955
rect 235994 1952 236000 1964
rect 235951 1924 236000 1952
rect 235951 1921 235963 1924
rect 235905 1915 235963 1921
rect 235092 1884 235120 1915
rect 235994 1912 236000 1924
rect 236052 1952 236058 1964
rect 236733 1955 236791 1961
rect 236733 1952 236745 1955
rect 236052 1924 236745 1952
rect 236052 1912 236058 1924
rect 236733 1921 236745 1924
rect 236779 1921 236791 1955
rect 236733 1915 236791 1921
rect 236917 1955 236975 1961
rect 236917 1921 236929 1955
rect 236963 1952 236975 1955
rect 237377 1955 237435 1961
rect 237377 1952 237389 1955
rect 236963 1924 237389 1952
rect 236963 1921 236975 1924
rect 236917 1915 236975 1921
rect 237377 1921 237389 1924
rect 237423 1921 237435 1955
rect 237377 1915 237435 1921
rect 237926 1912 237932 1964
rect 237984 1952 237990 1964
rect 238220 1952 238248 1992
rect 237984 1924 238248 1952
rect 237984 1912 237990 1924
rect 240042 1912 240048 1964
rect 240100 1952 240106 1964
rect 241517 1955 241575 1961
rect 241517 1952 241529 1955
rect 240100 1924 241529 1952
rect 240100 1912 240106 1924
rect 241517 1921 241529 1924
rect 241563 1921 241575 1955
rect 241624 1952 241652 1992
rect 243170 1980 243176 2032
rect 243228 2020 243234 2032
rect 257798 2020 257804 2032
rect 243228 1992 257804 2020
rect 243228 1980 243234 1992
rect 257798 1980 257804 1992
rect 257856 2020 257862 2032
rect 259086 2020 259092 2032
rect 257856 1992 258028 2020
rect 257856 1980 257862 1992
rect 250257 1955 250315 1961
rect 250257 1952 250269 1955
rect 241624 1924 250269 1952
rect 241517 1915 241575 1921
rect 250257 1921 250269 1924
rect 250303 1921 250315 1955
rect 250257 1915 250315 1921
rect 251174 1912 251180 1964
rect 251232 1952 251238 1964
rect 251361 1955 251419 1961
rect 251361 1952 251373 1955
rect 251232 1924 251373 1952
rect 251232 1912 251238 1924
rect 251361 1921 251373 1924
rect 251407 1921 251419 1955
rect 251361 1915 251419 1921
rect 252554 1912 252560 1964
rect 252612 1912 252618 1964
rect 255406 1912 255412 1964
rect 255464 1912 255470 1964
rect 256697 1955 256755 1961
rect 256697 1921 256709 1955
rect 256743 1952 256755 1955
rect 256878 1952 256884 1964
rect 256743 1924 256884 1952
rect 256743 1921 256755 1924
rect 256697 1915 256755 1921
rect 256878 1912 256884 1924
rect 256936 1912 256942 1964
rect 257890 1912 257896 1964
rect 257948 1912 257954 1964
rect 258000 1952 258028 1992
rect 258828 1992 259092 2020
rect 258828 1952 258856 1992
rect 259086 1980 259092 1992
rect 259144 2020 259150 2032
rect 259564 2020 259592 2060
rect 259144 1992 259592 2020
rect 259144 1980 259150 1992
rect 258000 1924 258856 1952
rect 258902 1912 258908 1964
rect 258960 1952 258966 1964
rect 259196 1961 259224 1992
rect 258997 1955 259055 1961
rect 258997 1952 259009 1955
rect 258960 1924 259009 1952
rect 258960 1912 258966 1924
rect 258997 1921 259009 1924
rect 259043 1921 259055 1955
rect 258997 1915 259055 1921
rect 259181 1955 259239 1961
rect 259181 1921 259193 1955
rect 259227 1921 259239 1955
rect 259181 1915 259239 1921
rect 259822 1912 259828 1964
rect 259880 1952 259886 1964
rect 260024 1961 260052 2060
rect 261570 2048 261576 2100
rect 261628 2088 261634 2100
rect 261849 2091 261907 2097
rect 261849 2088 261861 2091
rect 261628 2060 261861 2088
rect 261628 2048 261634 2060
rect 261849 2057 261861 2060
rect 261895 2057 261907 2091
rect 261849 2051 261907 2057
rect 269666 2048 269672 2100
rect 269724 2048 269730 2100
rect 269758 2048 269764 2100
rect 269816 2088 269822 2100
rect 269816 2060 270356 2088
rect 269816 2048 269822 2060
rect 260098 1980 260104 2032
rect 260156 2020 260162 2032
rect 264146 2020 264152 2032
rect 260156 1992 264152 2020
rect 260156 1980 260162 1992
rect 264146 1980 264152 1992
rect 264204 1980 264210 2032
rect 267550 1980 267556 2032
rect 267608 2020 267614 2032
rect 267608 1992 270264 2020
rect 267608 1980 267614 1992
rect 259917 1955 259975 1961
rect 259917 1952 259929 1955
rect 259880 1924 259929 1952
rect 259880 1912 259886 1924
rect 259917 1921 259929 1924
rect 259963 1921 259975 1955
rect 259917 1915 259975 1921
rect 260009 1955 260067 1961
rect 260009 1921 260021 1955
rect 260055 1952 260067 1955
rect 260055 1924 260236 1952
rect 260055 1921 260067 1924
rect 260009 1915 260067 1921
rect 234264 1856 235120 1884
rect 235718 1844 235724 1896
rect 235776 1844 235782 1896
rect 235810 1844 235816 1896
rect 235868 1884 235874 1896
rect 236549 1887 236607 1893
rect 236549 1884 236561 1887
rect 235868 1856 236561 1884
rect 235868 1844 235874 1856
rect 236549 1853 236561 1856
rect 236595 1853 236607 1887
rect 236549 1847 236607 1853
rect 241238 1844 241244 1896
rect 241296 1844 241302 1896
rect 242894 1844 242900 1896
rect 242952 1884 242958 1896
rect 243541 1887 243599 1893
rect 243541 1884 243553 1887
rect 242952 1856 243553 1884
rect 242952 1844 242958 1856
rect 243541 1853 243553 1856
rect 243587 1853 243599 1887
rect 243541 1847 243599 1853
rect 243814 1844 243820 1896
rect 243872 1844 243878 1896
rect 244274 1844 244280 1896
rect 244332 1884 244338 1896
rect 244829 1887 244887 1893
rect 244829 1884 244841 1887
rect 244332 1856 244841 1884
rect 244332 1844 244338 1856
rect 244829 1853 244841 1856
rect 244875 1853 244887 1887
rect 244829 1847 244887 1853
rect 246114 1844 246120 1896
rect 246172 1844 246178 1896
rect 246393 1887 246451 1893
rect 246393 1853 246405 1887
rect 246439 1853 246451 1887
rect 246393 1847 246451 1853
rect 239490 1816 239496 1828
rect 225156 1788 233740 1816
rect 233988 1788 239496 1816
rect 159453 1751 159511 1757
rect 159453 1748 159465 1751
rect 156340 1720 159465 1748
rect 156141 1711 156199 1717
rect 159453 1717 159465 1720
rect 159499 1717 159511 1751
rect 159453 1711 159511 1717
rect 160186 1708 160192 1760
rect 160244 1748 160250 1760
rect 160281 1751 160339 1757
rect 160281 1748 160293 1751
rect 160244 1720 160293 1748
rect 160244 1708 160250 1720
rect 160281 1717 160293 1720
rect 160327 1717 160339 1751
rect 160281 1711 160339 1717
rect 161474 1708 161480 1760
rect 161532 1708 161538 1760
rect 163130 1708 163136 1760
rect 163188 1708 163194 1760
rect 164510 1708 164516 1760
rect 164568 1748 164574 1760
rect 164789 1751 164847 1757
rect 164789 1748 164801 1751
rect 164568 1720 164801 1748
rect 164568 1708 164574 1720
rect 164789 1717 164801 1720
rect 164835 1717 164847 1751
rect 164789 1711 164847 1717
rect 168374 1708 168380 1760
rect 168432 1748 168438 1760
rect 168929 1751 168987 1757
rect 168929 1748 168941 1751
rect 168432 1720 168941 1748
rect 168432 1708 168438 1720
rect 168929 1717 168941 1720
rect 168975 1717 168987 1751
rect 168929 1711 168987 1717
rect 181990 1708 181996 1760
rect 182048 1708 182054 1760
rect 193214 1708 193220 1760
rect 193272 1708 193278 1760
rect 193306 1708 193312 1760
rect 193364 1748 193370 1760
rect 194045 1751 194103 1757
rect 194045 1748 194057 1751
rect 193364 1720 194057 1748
rect 193364 1708 193370 1720
rect 194045 1717 194057 1720
rect 194091 1717 194103 1751
rect 194045 1711 194103 1717
rect 194594 1708 194600 1760
rect 194652 1748 194658 1760
rect 194873 1751 194931 1757
rect 194873 1748 194885 1751
rect 194652 1720 194885 1748
rect 194652 1708 194658 1720
rect 194873 1717 194885 1720
rect 194919 1717 194931 1751
rect 194873 1711 194931 1717
rect 196526 1708 196532 1760
rect 196584 1708 196590 1760
rect 197906 1708 197912 1760
rect 197964 1748 197970 1760
rect 198369 1751 198427 1757
rect 198369 1748 198381 1751
rect 197964 1720 198381 1748
rect 197964 1708 197970 1720
rect 198369 1717 198381 1720
rect 198415 1717 198427 1751
rect 198369 1711 198427 1717
rect 199746 1708 199752 1760
rect 199804 1748 199810 1760
rect 200025 1751 200083 1757
rect 200025 1748 200037 1751
rect 199804 1720 200037 1748
rect 199804 1708 199810 1720
rect 200025 1717 200037 1720
rect 200071 1717 200083 1751
rect 200025 1711 200083 1717
rect 201678 1708 201684 1760
rect 201736 1708 201742 1760
rect 202874 1708 202880 1760
rect 202932 1748 202938 1760
rect 203337 1751 203395 1757
rect 203337 1748 203349 1751
rect 202932 1720 203349 1748
rect 202932 1708 202938 1720
rect 203337 1717 203349 1720
rect 203383 1717 203395 1751
rect 203337 1711 203395 1717
rect 216122 1708 216128 1760
rect 216180 1748 216186 1760
rect 224310 1748 224316 1760
rect 216180 1720 224316 1748
rect 216180 1708 216186 1720
rect 224310 1708 224316 1720
rect 224368 1708 224374 1760
rect 225506 1708 225512 1760
rect 225564 1748 225570 1760
rect 229186 1748 229192 1760
rect 225564 1720 229192 1748
rect 225564 1708 225570 1720
rect 229186 1708 229192 1720
rect 229244 1708 229250 1760
rect 229278 1708 229284 1760
rect 229336 1708 229342 1760
rect 229646 1708 229652 1760
rect 229704 1748 229710 1760
rect 230109 1751 230167 1757
rect 230109 1748 230121 1751
rect 229704 1720 230121 1748
rect 229704 1708 229710 1720
rect 230109 1717 230121 1720
rect 230155 1717 230167 1751
rect 230109 1711 230167 1717
rect 230658 1708 230664 1760
rect 230716 1748 230722 1760
rect 230937 1751 230995 1757
rect 230937 1748 230949 1751
rect 230716 1720 230949 1748
rect 230716 1708 230722 1720
rect 230937 1717 230949 1720
rect 230983 1717 230995 1751
rect 230937 1711 230995 1717
rect 231578 1708 231584 1760
rect 231636 1748 231642 1760
rect 232314 1748 232320 1760
rect 231636 1720 232320 1748
rect 231636 1708 231642 1720
rect 232314 1708 232320 1720
rect 232372 1708 232378 1760
rect 233234 1708 233240 1760
rect 233292 1748 233298 1760
rect 233605 1751 233663 1757
rect 233605 1748 233617 1751
rect 233292 1720 233617 1748
rect 233292 1708 233298 1720
rect 233605 1717 233617 1720
rect 233651 1717 233663 1751
rect 233712 1748 233740 1788
rect 239490 1776 239496 1788
rect 239548 1776 239554 1828
rect 242526 1776 242532 1828
rect 242584 1816 242590 1828
rect 246408 1816 246436 1847
rect 248414 1844 248420 1896
rect 248472 1884 248478 1896
rect 248693 1887 248751 1893
rect 248693 1884 248705 1887
rect 248472 1856 248705 1884
rect 248472 1844 248478 1856
rect 248693 1853 248705 1856
rect 248739 1853 248751 1887
rect 248693 1847 248751 1853
rect 248966 1844 248972 1896
rect 249024 1844 249030 1896
rect 249794 1844 249800 1896
rect 249852 1884 249858 1896
rect 249981 1887 250039 1893
rect 249981 1884 249993 1887
rect 249852 1856 249993 1884
rect 249852 1844 249858 1856
rect 249981 1853 249993 1856
rect 250027 1853 250039 1887
rect 249981 1847 250039 1853
rect 252278 1844 252284 1896
rect 252336 1844 252342 1896
rect 253842 1844 253848 1896
rect 253900 1844 253906 1896
rect 254026 1844 254032 1896
rect 254084 1884 254090 1896
rect 254121 1887 254179 1893
rect 254121 1884 254133 1887
rect 254084 1856 254133 1884
rect 254084 1844 254090 1856
rect 254121 1853 254133 1856
rect 254167 1853 254179 1887
rect 254121 1847 254179 1853
rect 255130 1844 255136 1896
rect 255188 1844 255194 1896
rect 256418 1844 256424 1896
rect 256476 1844 256482 1896
rect 260208 1884 260236 1924
rect 260282 1912 260288 1964
rect 260340 1952 260346 1964
rect 260653 1955 260711 1961
rect 260653 1952 260665 1955
rect 260340 1924 260665 1952
rect 260340 1912 260346 1924
rect 260653 1921 260665 1924
rect 260699 1921 260711 1955
rect 260653 1915 260711 1921
rect 260837 1955 260895 1961
rect 260837 1921 260849 1955
rect 260883 1921 260895 1955
rect 260837 1915 260895 1921
rect 260852 1884 260880 1915
rect 261478 1912 261484 1964
rect 261536 1912 261542 1964
rect 261665 1955 261723 1961
rect 261665 1921 261677 1955
rect 261711 1921 261723 1955
rect 261665 1915 261723 1921
rect 261680 1884 261708 1915
rect 262306 1912 262312 1964
rect 262364 1912 262370 1964
rect 262493 1955 262551 1961
rect 262493 1921 262505 1955
rect 262539 1921 262551 1955
rect 262493 1915 262551 1921
rect 262508 1884 262536 1915
rect 262582 1912 262588 1964
rect 262640 1952 262646 1964
rect 263137 1955 263195 1961
rect 263137 1952 263149 1955
rect 262640 1924 263149 1952
rect 262640 1912 262646 1924
rect 263137 1921 263149 1924
rect 263183 1921 263195 1955
rect 263137 1915 263195 1921
rect 263321 1955 263379 1961
rect 263321 1921 263333 1955
rect 263367 1952 263379 1955
rect 264238 1952 264244 1964
rect 263367 1924 264244 1952
rect 263367 1921 263379 1924
rect 263321 1915 263379 1921
rect 263336 1884 263364 1915
rect 264238 1912 264244 1924
rect 264296 1952 264302 1964
rect 264333 1955 264391 1961
rect 264333 1952 264345 1955
rect 264296 1924 264345 1952
rect 264296 1912 264302 1924
rect 264333 1921 264345 1924
rect 264379 1952 264391 1955
rect 265161 1955 265219 1961
rect 265161 1952 265173 1955
rect 264379 1924 265173 1952
rect 264379 1921 264391 1924
rect 264333 1915 264391 1921
rect 265161 1921 265173 1924
rect 265207 1952 265219 1955
rect 265989 1955 266047 1961
rect 265989 1952 266001 1955
rect 265207 1924 266001 1952
rect 265207 1921 265219 1924
rect 265161 1915 265219 1921
rect 265989 1921 266001 1924
rect 266035 1952 266047 1955
rect 266817 1955 266875 1961
rect 266817 1952 266829 1955
rect 266035 1924 266829 1952
rect 266035 1921 266047 1924
rect 265989 1915 266047 1921
rect 266817 1921 266829 1924
rect 266863 1952 266875 1955
rect 267645 1955 267703 1961
rect 267645 1952 267657 1955
rect 266863 1924 267657 1952
rect 266863 1921 266875 1924
rect 266817 1915 266875 1921
rect 267645 1921 267657 1924
rect 267691 1952 267703 1955
rect 268473 1955 268531 1961
rect 268473 1952 268485 1955
rect 267691 1924 268485 1952
rect 267691 1921 267703 1924
rect 267645 1915 267703 1921
rect 268473 1921 268485 1924
rect 268519 1952 268531 1955
rect 269206 1952 269212 1964
rect 268519 1924 269212 1952
rect 268519 1921 268531 1924
rect 268473 1915 268531 1921
rect 269206 1912 269212 1924
rect 269264 1952 269270 1964
rect 269485 1955 269543 1961
rect 269485 1952 269497 1955
rect 269264 1924 269497 1952
rect 269264 1912 269270 1924
rect 269485 1921 269497 1924
rect 269531 1952 269543 1955
rect 269758 1952 269764 1964
rect 269531 1924 269764 1952
rect 269531 1921 269543 1924
rect 269485 1915 269543 1921
rect 269758 1912 269764 1924
rect 269816 1912 269822 1964
rect 270236 1961 270264 1992
rect 270328 1961 270356 2060
rect 270494 2048 270500 2100
rect 270552 2048 270558 2100
rect 271138 1980 271144 2032
rect 271196 2020 271202 2032
rect 272150 2020 272156 2032
rect 271196 1992 272156 2020
rect 271196 1980 271202 1992
rect 272150 1980 272156 1992
rect 272208 1980 272214 2032
rect 270221 1955 270279 1961
rect 270221 1921 270233 1955
rect 270267 1921 270279 1955
rect 270221 1915 270279 1921
rect 270313 1955 270371 1961
rect 270313 1921 270325 1955
rect 270359 1921 270371 1955
rect 270313 1915 270371 1921
rect 260208 1856 263364 1884
rect 263410 1844 263416 1896
rect 263468 1884 263474 1896
rect 264149 1887 264207 1893
rect 264149 1884 264161 1887
rect 263468 1856 264161 1884
rect 263468 1844 263474 1856
rect 264149 1853 264161 1856
rect 264195 1853 264207 1887
rect 264149 1847 264207 1853
rect 264977 1887 265035 1893
rect 264977 1853 264989 1887
rect 265023 1884 265035 1887
rect 265066 1884 265072 1896
rect 265023 1856 265072 1884
rect 265023 1853 265035 1856
rect 264977 1847 265035 1853
rect 265066 1844 265072 1856
rect 265124 1844 265130 1896
rect 265802 1844 265808 1896
rect 265860 1844 265866 1896
rect 266630 1844 266636 1896
rect 266688 1844 266694 1896
rect 266722 1844 266728 1896
rect 266780 1884 266786 1896
rect 267461 1887 267519 1893
rect 267461 1884 267473 1887
rect 266780 1856 267473 1884
rect 266780 1844 266786 1856
rect 267461 1853 267473 1856
rect 267507 1853 267519 1887
rect 267461 1847 267519 1853
rect 268286 1844 268292 1896
rect 268344 1844 268350 1896
rect 269301 1887 269359 1893
rect 269301 1853 269313 1887
rect 269347 1884 269359 1887
rect 270862 1884 270868 1896
rect 269347 1856 270868 1884
rect 269347 1853 269359 1856
rect 269301 1847 269359 1853
rect 270862 1844 270868 1856
rect 270920 1844 270926 1896
rect 242584 1788 246436 1816
rect 242584 1776 242590 1788
rect 259270 1776 259276 1828
rect 259328 1816 259334 1828
rect 269022 1816 269028 1828
rect 259328 1788 269028 1816
rect 259328 1776 259334 1788
rect 269022 1776 269028 1788
rect 269080 1776 269086 1828
rect 233878 1748 233884 1760
rect 233712 1720 233884 1748
rect 233605 1711 233663 1717
rect 233878 1708 233884 1720
rect 233936 1708 233942 1760
rect 233970 1708 233976 1760
rect 234028 1748 234034 1760
rect 234433 1751 234491 1757
rect 234433 1748 234445 1751
rect 234028 1720 234445 1748
rect 234028 1708 234034 1720
rect 234433 1717 234445 1720
rect 234479 1717 234491 1751
rect 234433 1711 234491 1717
rect 234706 1708 234712 1760
rect 234764 1748 234770 1760
rect 235261 1751 235319 1757
rect 235261 1748 235273 1751
rect 234764 1720 235273 1748
rect 234764 1708 234770 1720
rect 235261 1717 235273 1720
rect 235307 1717 235319 1751
rect 235261 1711 235319 1717
rect 237282 1708 237288 1760
rect 237340 1748 237346 1760
rect 237561 1751 237619 1757
rect 237561 1748 237573 1751
rect 237340 1720 237573 1748
rect 237340 1708 237346 1720
rect 237561 1717 237573 1720
rect 237607 1717 237619 1751
rect 237561 1711 237619 1717
rect 257890 1708 257896 1760
rect 257948 1748 257954 1760
rect 260098 1748 260104 1760
rect 257948 1720 260104 1748
rect 257948 1708 257954 1720
rect 260098 1708 260104 1720
rect 260156 1708 260162 1760
rect 260193 1751 260251 1757
rect 260193 1717 260205 1751
rect 260239 1748 260251 1751
rect 260282 1748 260288 1760
rect 260239 1720 260288 1748
rect 260239 1717 260251 1720
rect 260193 1711 260251 1717
rect 260282 1708 260288 1720
rect 260340 1708 260346 1760
rect 261021 1751 261079 1757
rect 261021 1717 261033 1751
rect 261067 1748 261079 1751
rect 261570 1748 261576 1760
rect 261067 1720 261576 1748
rect 261067 1717 261079 1720
rect 261021 1711 261079 1717
rect 261570 1708 261576 1720
rect 261628 1708 261634 1760
rect 262306 1708 262312 1760
rect 262364 1748 262370 1760
rect 262677 1751 262735 1757
rect 262677 1748 262689 1751
rect 262364 1720 262689 1748
rect 262364 1708 262370 1720
rect 262677 1717 262689 1720
rect 262723 1717 262735 1751
rect 262677 1711 262735 1717
rect 263042 1708 263048 1760
rect 263100 1748 263106 1760
rect 263505 1751 263563 1757
rect 263505 1748 263517 1751
rect 263100 1720 263517 1748
rect 263100 1708 263106 1720
rect 263505 1717 263517 1720
rect 263551 1717 263563 1751
rect 263505 1711 263563 1717
rect 264146 1708 264152 1760
rect 264204 1748 264210 1760
rect 264517 1751 264575 1757
rect 264517 1748 264529 1751
rect 264204 1720 264529 1748
rect 264204 1708 264210 1720
rect 264517 1717 264529 1720
rect 264563 1717 264575 1751
rect 264517 1711 264575 1717
rect 265158 1708 265164 1760
rect 265216 1748 265222 1760
rect 265345 1751 265403 1757
rect 265345 1748 265357 1751
rect 265216 1720 265357 1748
rect 265216 1708 265222 1720
rect 265345 1717 265357 1720
rect 265391 1717 265403 1751
rect 265345 1711 265403 1717
rect 265894 1708 265900 1760
rect 265952 1748 265958 1760
rect 266173 1751 266231 1757
rect 266173 1748 266185 1751
rect 265952 1720 266185 1748
rect 265952 1708 265958 1720
rect 266173 1717 266185 1720
rect 266219 1717 266231 1751
rect 266173 1711 266231 1717
rect 266722 1708 266728 1760
rect 266780 1748 266786 1760
rect 267001 1751 267059 1757
rect 267001 1748 267013 1751
rect 266780 1720 267013 1748
rect 266780 1708 266786 1720
rect 267001 1717 267013 1720
rect 267047 1717 267059 1751
rect 267001 1711 267059 1717
rect 267826 1708 267832 1760
rect 267884 1708 267890 1760
rect 268194 1708 268200 1760
rect 268252 1748 268258 1760
rect 268657 1751 268715 1757
rect 268657 1748 268669 1751
rect 268252 1720 268669 1748
rect 268252 1708 268258 1720
rect 268657 1717 268669 1720
rect 268703 1717 268715 1751
rect 268657 1711 268715 1717
rect 1104 1658 271492 1680
rect 1104 1606 34748 1658
rect 34800 1606 34812 1658
rect 34864 1606 34876 1658
rect 34928 1606 34940 1658
rect 34992 1606 35004 1658
rect 35056 1606 102345 1658
rect 102397 1606 102409 1658
rect 102461 1606 102473 1658
rect 102525 1606 102537 1658
rect 102589 1606 102601 1658
rect 102653 1606 169942 1658
rect 169994 1606 170006 1658
rect 170058 1606 170070 1658
rect 170122 1606 170134 1658
rect 170186 1606 170198 1658
rect 170250 1606 237539 1658
rect 237591 1606 237603 1658
rect 237655 1606 237667 1658
rect 237719 1606 237731 1658
rect 237783 1606 237795 1658
rect 237847 1606 271492 1658
rect 1104 1584 271492 1606
rect 22094 1504 22100 1556
rect 22152 1544 22158 1556
rect 25961 1547 26019 1553
rect 25961 1544 25973 1547
rect 22152 1516 25973 1544
rect 22152 1504 22158 1516
rect 25961 1513 25973 1516
rect 26007 1513 26019 1547
rect 25961 1507 26019 1513
rect 28353 1547 28411 1553
rect 28353 1513 28365 1547
rect 28399 1544 28411 1547
rect 28534 1544 28540 1556
rect 28399 1516 28540 1544
rect 28399 1513 28411 1516
rect 28353 1507 28411 1513
rect 28534 1504 28540 1516
rect 28592 1504 28598 1556
rect 35437 1547 35495 1553
rect 35437 1513 35449 1547
rect 35483 1544 35495 1547
rect 35526 1544 35532 1556
rect 35483 1516 35532 1544
rect 35483 1513 35495 1516
rect 35437 1507 35495 1513
rect 35526 1504 35532 1516
rect 35584 1504 35590 1556
rect 35618 1504 35624 1556
rect 35676 1544 35682 1556
rect 58894 1544 58900 1556
rect 35676 1516 58900 1544
rect 35676 1504 35682 1516
rect 58894 1504 58900 1516
rect 58952 1504 58958 1556
rect 59998 1504 60004 1556
rect 60056 1504 60062 1556
rect 94406 1504 94412 1556
rect 94464 1544 94470 1556
rect 95145 1547 95203 1553
rect 95145 1544 95157 1547
rect 94464 1516 95157 1544
rect 94464 1504 94470 1516
rect 95145 1513 95157 1516
rect 95191 1513 95203 1547
rect 95145 1507 95203 1513
rect 95234 1504 95240 1556
rect 95292 1544 95298 1556
rect 99190 1544 99196 1556
rect 95292 1516 99196 1544
rect 95292 1504 95298 1516
rect 99190 1504 99196 1516
rect 99248 1504 99254 1556
rect 99374 1504 99380 1556
rect 99432 1544 99438 1556
rect 107378 1544 107384 1556
rect 99432 1516 107384 1544
rect 99432 1504 99438 1516
rect 107378 1504 107384 1516
rect 107436 1504 107442 1556
rect 113266 1504 113272 1556
rect 113324 1544 113330 1556
rect 113361 1547 113419 1553
rect 113361 1544 113373 1547
rect 113324 1516 113373 1544
rect 113324 1504 113330 1516
rect 113361 1513 113373 1516
rect 113407 1513 113419 1547
rect 113361 1507 113419 1513
rect 121638 1504 121644 1556
rect 121696 1544 121702 1556
rect 156506 1544 156512 1556
rect 121696 1516 156512 1544
rect 121696 1504 121702 1516
rect 156506 1504 156512 1516
rect 156564 1504 156570 1556
rect 156690 1504 156696 1556
rect 156748 1544 156754 1556
rect 156785 1547 156843 1553
rect 156785 1544 156797 1547
rect 156748 1516 156797 1544
rect 156748 1504 156754 1516
rect 156785 1513 156797 1516
rect 156831 1513 156843 1547
rect 156785 1507 156843 1513
rect 157334 1504 157340 1556
rect 157392 1544 157398 1556
rect 157613 1547 157671 1553
rect 157613 1544 157625 1547
rect 157392 1516 157625 1544
rect 157392 1504 157398 1516
rect 157613 1513 157625 1516
rect 157659 1513 157671 1547
rect 157613 1507 157671 1513
rect 175826 1504 175832 1556
rect 175884 1544 175890 1556
rect 175884 1516 177068 1544
rect 175884 1504 175890 1516
rect 23658 1436 23664 1488
rect 23716 1476 23722 1488
rect 30926 1476 30932 1488
rect 23716 1448 30932 1476
rect 23716 1436 23722 1448
rect 30926 1436 30932 1448
rect 30984 1436 30990 1488
rect 31018 1436 31024 1488
rect 31076 1476 31082 1488
rect 31076 1448 35894 1476
rect 31076 1436 31082 1448
rect 842 1368 848 1420
rect 900 1408 906 1420
rect 1765 1411 1823 1417
rect 1765 1408 1777 1411
rect 900 1380 1777 1408
rect 900 1368 906 1380
rect 1765 1377 1777 1380
rect 1811 1377 1823 1411
rect 1765 1371 1823 1377
rect 24026 1368 24032 1420
rect 24084 1408 24090 1420
rect 24946 1408 24952 1420
rect 24084 1380 24952 1408
rect 24084 1368 24090 1380
rect 2593 1343 2651 1349
rect 2593 1309 2605 1343
rect 2639 1309 2651 1343
rect 2593 1303 2651 1309
rect 2608 1272 2636 1303
rect 2866 1300 2872 1352
rect 2924 1300 2930 1352
rect 5166 1300 5172 1352
rect 5224 1300 5230 1352
rect 5442 1300 5448 1352
rect 5500 1300 5506 1352
rect 6546 1300 6552 1352
rect 6604 1300 6610 1352
rect 6825 1343 6883 1349
rect 6825 1309 6837 1343
rect 6871 1340 6883 1343
rect 9398 1340 9404 1352
rect 6871 1312 9404 1340
rect 6871 1309 6883 1312
rect 6825 1303 6883 1309
rect 9398 1300 9404 1312
rect 9456 1300 9462 1352
rect 9493 1343 9551 1349
rect 9493 1309 9505 1343
rect 9539 1340 9551 1343
rect 9582 1340 9588 1352
rect 9539 1312 9588 1340
rect 9539 1309 9551 1312
rect 9493 1303 9551 1309
rect 9582 1300 9588 1312
rect 9640 1300 9646 1352
rect 11146 1300 11152 1352
rect 11204 1300 11210 1352
rect 12158 1300 12164 1352
rect 12216 1300 12222 1352
rect 14826 1300 14832 1352
rect 14884 1300 14890 1352
rect 15102 1300 15108 1352
rect 15160 1300 15166 1352
rect 23750 1300 23756 1352
rect 23808 1300 23814 1352
rect 24688 1349 24716 1380
rect 24946 1368 24952 1380
rect 25004 1368 25010 1420
rect 25038 1368 25044 1420
rect 25096 1408 25102 1420
rect 25096 1380 25176 1408
rect 25096 1368 25102 1380
rect 25148 1349 25176 1380
rect 25866 1368 25872 1420
rect 25924 1408 25930 1420
rect 27157 1411 27215 1417
rect 27157 1408 27169 1411
rect 25924 1380 27169 1408
rect 25924 1368 25930 1380
rect 27157 1377 27169 1380
rect 27203 1377 27215 1411
rect 27157 1371 27215 1377
rect 27798 1368 27804 1420
rect 27856 1408 27862 1420
rect 27985 1411 28043 1417
rect 27985 1408 27997 1411
rect 27856 1380 27997 1408
rect 27856 1368 27862 1380
rect 27985 1377 27997 1380
rect 28031 1377 28043 1411
rect 27985 1371 28043 1377
rect 34333 1411 34391 1417
rect 34333 1377 34345 1411
rect 34379 1408 34391 1411
rect 34422 1408 34428 1420
rect 34379 1380 34428 1408
rect 34379 1377 34391 1380
rect 34333 1371 34391 1377
rect 34422 1368 34428 1380
rect 34480 1368 34486 1420
rect 35866 1408 35894 1448
rect 36722 1436 36728 1488
rect 36780 1436 36786 1488
rect 38654 1436 38660 1488
rect 38712 1436 38718 1488
rect 43346 1436 43352 1488
rect 43404 1476 43410 1488
rect 44453 1479 44511 1485
rect 44453 1476 44465 1479
rect 43404 1448 44465 1476
rect 43404 1436 43410 1448
rect 44453 1445 44465 1448
rect 44499 1445 44511 1479
rect 54110 1476 54116 1488
rect 44453 1439 44511 1445
rect 53944 1448 54116 1476
rect 53466 1408 53472 1420
rect 35866 1380 53472 1408
rect 53466 1368 53472 1380
rect 53524 1368 53530 1420
rect 53944 1417 53972 1448
rect 54110 1436 54116 1448
rect 54168 1436 54174 1488
rect 86034 1436 86040 1488
rect 86092 1476 86098 1488
rect 99006 1476 99012 1488
rect 86092 1448 99012 1476
rect 86092 1436 86098 1448
rect 99006 1436 99012 1448
rect 99064 1436 99070 1488
rect 101582 1436 101588 1488
rect 101640 1476 101646 1488
rect 133230 1476 133236 1488
rect 101640 1448 133236 1476
rect 101640 1436 101646 1448
rect 133230 1436 133236 1448
rect 133288 1436 133294 1488
rect 133322 1436 133328 1488
rect 133380 1436 133386 1488
rect 134334 1436 134340 1488
rect 134392 1436 134398 1488
rect 138014 1436 138020 1488
rect 138072 1476 138078 1488
rect 138109 1479 138167 1485
rect 138109 1476 138121 1479
rect 138072 1448 138121 1476
rect 138072 1436 138078 1448
rect 138109 1445 138121 1448
rect 138155 1445 138167 1479
rect 138109 1439 138167 1445
rect 138290 1436 138296 1488
rect 138348 1476 138354 1488
rect 139213 1479 139271 1485
rect 139213 1476 139225 1479
rect 138348 1448 139225 1476
rect 138348 1436 138354 1448
rect 139213 1445 139225 1448
rect 139259 1445 139271 1479
rect 139213 1439 139271 1445
rect 140501 1479 140559 1485
rect 140501 1445 140513 1479
rect 140547 1476 140559 1479
rect 140682 1476 140688 1488
rect 140547 1448 140688 1476
rect 140547 1445 140559 1448
rect 140501 1439 140559 1445
rect 140682 1436 140688 1448
rect 140740 1436 140746 1488
rect 144178 1436 144184 1488
rect 144236 1476 144242 1488
rect 176930 1476 176936 1488
rect 144236 1448 176936 1476
rect 144236 1436 144242 1448
rect 176930 1436 176936 1448
rect 176988 1436 176994 1488
rect 177040 1476 177068 1516
rect 180610 1504 180616 1556
rect 180668 1504 180674 1556
rect 216582 1544 216588 1556
rect 180766 1516 216588 1544
rect 180766 1476 180794 1516
rect 216582 1504 216588 1516
rect 216640 1504 216646 1556
rect 220630 1504 220636 1556
rect 220688 1544 220694 1556
rect 221645 1547 221703 1553
rect 221645 1544 221657 1547
rect 220688 1516 221657 1544
rect 220688 1504 220694 1516
rect 221645 1513 221657 1516
rect 221691 1513 221703 1547
rect 221645 1507 221703 1513
rect 225877 1547 225935 1553
rect 225877 1513 225889 1547
rect 225923 1544 225935 1547
rect 226242 1544 226248 1556
rect 225923 1516 226248 1544
rect 225923 1513 225935 1516
rect 225877 1507 225935 1513
rect 226242 1504 226248 1516
rect 226300 1504 226306 1556
rect 226426 1504 226432 1556
rect 226484 1544 226490 1556
rect 228453 1547 228511 1553
rect 226484 1516 228404 1544
rect 226484 1504 226490 1516
rect 177040 1448 180794 1476
rect 191374 1436 191380 1488
rect 191432 1436 191438 1488
rect 213273 1479 213331 1485
rect 213273 1445 213285 1479
rect 213319 1445 213331 1479
rect 213273 1439 213331 1445
rect 53929 1411 53987 1417
rect 53929 1377 53941 1411
rect 53975 1377 53987 1411
rect 53929 1371 53987 1377
rect 69106 1368 69112 1420
rect 69164 1368 69170 1420
rect 87782 1368 87788 1420
rect 87840 1408 87846 1420
rect 88061 1411 88119 1417
rect 88061 1408 88073 1411
rect 87840 1380 88073 1408
rect 87840 1368 87846 1380
rect 88061 1377 88073 1380
rect 88107 1377 88119 1411
rect 88518 1408 88524 1420
rect 88061 1371 88119 1377
rect 88260 1380 88524 1408
rect 24673 1343 24731 1349
rect 24673 1309 24685 1343
rect 24719 1309 24731 1343
rect 24673 1303 24731 1309
rect 25133 1343 25191 1349
rect 25133 1309 25145 1343
rect 25179 1340 25191 1343
rect 27341 1343 27399 1349
rect 27341 1340 27353 1343
rect 25179 1312 27353 1340
rect 25179 1309 25191 1312
rect 25133 1303 25191 1309
rect 27341 1309 27353 1312
rect 27387 1309 27399 1343
rect 27341 1303 27399 1309
rect 2958 1272 2964 1284
rect 2608 1244 2964 1272
rect 2958 1232 2964 1244
rect 3016 1232 3022 1284
rect 4062 1232 4068 1284
rect 4120 1232 4126 1284
rect 8202 1232 8208 1284
rect 8260 1272 8266 1284
rect 8297 1275 8355 1281
rect 8297 1272 8309 1275
rect 8260 1244 8309 1272
rect 8260 1232 8266 1244
rect 8297 1241 8309 1244
rect 8343 1241 8355 1275
rect 8297 1235 8355 1241
rect 9674 1232 9680 1284
rect 9732 1232 9738 1284
rect 10226 1232 10232 1284
rect 10284 1232 10290 1284
rect 10410 1232 10416 1284
rect 10468 1232 10474 1284
rect 10962 1232 10968 1284
rect 11020 1232 11026 1284
rect 11974 1232 11980 1284
rect 12032 1232 12038 1284
rect 12710 1232 12716 1284
rect 12768 1232 12774 1284
rect 13446 1232 13452 1284
rect 13504 1232 13510 1284
rect 17126 1232 17132 1284
rect 17184 1232 17190 1284
rect 17862 1232 17868 1284
rect 17920 1232 17926 1284
rect 18598 1232 18604 1284
rect 18656 1232 18662 1284
rect 25317 1275 25375 1281
rect 25317 1241 25329 1275
rect 25363 1272 25375 1275
rect 25869 1275 25927 1281
rect 25869 1272 25881 1275
rect 25363 1244 25881 1272
rect 25363 1241 25375 1244
rect 25317 1235 25375 1241
rect 25869 1241 25881 1244
rect 25915 1241 25927 1275
rect 27356 1272 27384 1303
rect 27522 1300 27528 1352
rect 27580 1300 27586 1352
rect 28169 1343 28227 1349
rect 28169 1309 28181 1343
rect 28215 1309 28227 1343
rect 28169 1303 28227 1309
rect 28184 1272 28212 1303
rect 28902 1300 28908 1352
rect 28960 1300 28966 1352
rect 29730 1300 29736 1352
rect 29788 1300 29794 1352
rect 30558 1300 30564 1352
rect 30616 1300 30622 1352
rect 31389 1343 31447 1349
rect 31389 1309 31401 1343
rect 31435 1340 31447 1343
rect 31754 1340 31760 1352
rect 31435 1312 31760 1340
rect 31435 1309 31447 1312
rect 31389 1303 31447 1309
rect 31754 1300 31760 1312
rect 31812 1300 31818 1352
rect 32306 1300 32312 1352
rect 32364 1300 32370 1352
rect 35618 1300 35624 1352
rect 35676 1300 35682 1352
rect 36262 1300 36268 1352
rect 36320 1300 36326 1352
rect 36906 1300 36912 1352
rect 36964 1300 36970 1352
rect 38197 1343 38255 1349
rect 38197 1309 38209 1343
rect 38243 1340 38255 1343
rect 38562 1340 38568 1352
rect 38243 1312 38568 1340
rect 38243 1309 38255 1312
rect 38197 1303 38255 1309
rect 38562 1300 38568 1312
rect 38620 1300 38626 1352
rect 38838 1300 38844 1352
rect 38896 1300 38902 1352
rect 39485 1343 39543 1349
rect 39485 1309 39497 1343
rect 39531 1340 39543 1343
rect 39942 1340 39948 1352
rect 39531 1312 39948 1340
rect 39531 1309 39543 1312
rect 39485 1303 39543 1309
rect 39942 1300 39948 1312
rect 40000 1300 40006 1352
rect 40770 1300 40776 1352
rect 40828 1300 40834 1352
rect 41414 1300 41420 1352
rect 41472 1300 41478 1352
rect 42058 1300 42064 1352
rect 42116 1300 42122 1352
rect 43254 1300 43260 1352
rect 43312 1300 43318 1352
rect 43990 1300 43996 1352
rect 44048 1300 44054 1352
rect 44634 1300 44640 1352
rect 44692 1300 44698 1352
rect 45922 1300 45928 1352
rect 45980 1300 45986 1352
rect 46566 1300 46572 1352
rect 46624 1300 46630 1352
rect 47210 1300 47216 1352
rect 47268 1300 47274 1352
rect 48314 1300 48320 1352
rect 48372 1340 48378 1352
rect 48409 1343 48467 1349
rect 48409 1340 48421 1343
rect 48372 1312 48421 1340
rect 48372 1300 48378 1312
rect 48409 1309 48421 1312
rect 48455 1309 48467 1343
rect 48409 1303 48467 1309
rect 49142 1300 49148 1352
rect 49200 1300 49206 1352
rect 49786 1300 49792 1352
rect 49844 1300 49850 1352
rect 51074 1300 51080 1352
rect 51132 1300 51138 1352
rect 51718 1300 51724 1352
rect 51776 1300 51782 1352
rect 52362 1300 52368 1352
rect 52420 1300 52426 1352
rect 53193 1343 53251 1349
rect 53193 1309 53205 1343
rect 53239 1340 53251 1343
rect 53834 1340 53840 1352
rect 53239 1312 53840 1340
rect 53239 1309 53251 1312
rect 53193 1303 53251 1309
rect 53834 1300 53840 1312
rect 53892 1300 53898 1352
rect 54018 1300 54024 1352
rect 54076 1340 54082 1352
rect 54113 1343 54171 1349
rect 54113 1340 54125 1343
rect 54076 1312 54125 1340
rect 54076 1300 54082 1312
rect 54113 1309 54125 1312
rect 54159 1309 54171 1343
rect 54113 1303 54171 1309
rect 56042 1300 56048 1352
rect 56100 1300 56106 1352
rect 56870 1300 56876 1352
rect 56928 1300 56934 1352
rect 58434 1300 58440 1352
rect 58492 1300 58498 1352
rect 59357 1343 59415 1349
rect 59357 1309 59369 1343
rect 59403 1340 59415 1343
rect 59722 1340 59728 1352
rect 59403 1312 59728 1340
rect 59403 1309 59415 1312
rect 59357 1303 59415 1309
rect 59722 1300 59728 1312
rect 59780 1300 59786 1352
rect 59817 1343 59875 1349
rect 59817 1309 59829 1343
rect 59863 1340 59875 1343
rect 59906 1340 59912 1352
rect 59863 1312 59912 1340
rect 59863 1309 59875 1312
rect 59817 1303 59875 1309
rect 59906 1300 59912 1312
rect 59964 1300 59970 1352
rect 60642 1300 60648 1352
rect 60700 1300 60706 1352
rect 61378 1300 61384 1352
rect 61436 1300 61442 1352
rect 61838 1300 61844 1352
rect 61896 1340 61902 1352
rect 62117 1343 62175 1349
rect 62117 1340 62129 1343
rect 61896 1312 62129 1340
rect 61896 1300 61902 1312
rect 62117 1309 62129 1312
rect 62163 1309 62175 1343
rect 62117 1303 62175 1309
rect 63586 1300 63592 1352
rect 63644 1300 63650 1352
rect 64322 1300 64328 1352
rect 64380 1300 64386 1352
rect 65978 1300 65984 1352
rect 66036 1300 66042 1352
rect 69566 1300 69572 1352
rect 69624 1300 69630 1352
rect 69842 1300 69848 1352
rect 69900 1300 69906 1352
rect 72142 1300 72148 1352
rect 72200 1300 72206 1352
rect 72418 1300 72424 1352
rect 72476 1300 72482 1352
rect 74718 1300 74724 1352
rect 74776 1300 74782 1352
rect 74994 1300 75000 1352
rect 75052 1300 75058 1352
rect 77297 1343 77355 1349
rect 77297 1309 77309 1343
rect 77343 1309 77355 1343
rect 77297 1303 77355 1309
rect 27356 1244 28212 1272
rect 25869 1235 25927 1241
rect 42978 1232 42984 1284
rect 43036 1272 43042 1284
rect 43036 1244 43852 1272
rect 43036 1232 43042 1244
rect 4154 1164 4160 1216
rect 4212 1164 4218 1216
rect 8386 1164 8392 1216
rect 8444 1164 8450 1216
rect 12802 1164 12808 1216
rect 12860 1164 12866 1216
rect 13538 1164 13544 1216
rect 13596 1164 13602 1216
rect 17218 1164 17224 1216
rect 17276 1164 17282 1216
rect 17954 1164 17960 1216
rect 18012 1164 18018 1216
rect 18690 1164 18696 1216
rect 18748 1164 18754 1216
rect 23934 1164 23940 1216
rect 23992 1164 23998 1216
rect 28994 1164 29000 1216
rect 29052 1204 29058 1216
rect 29089 1207 29147 1213
rect 29089 1204 29101 1207
rect 29052 1176 29101 1204
rect 29052 1164 29058 1176
rect 29089 1173 29101 1176
rect 29135 1173 29147 1207
rect 29089 1167 29147 1173
rect 29914 1164 29920 1216
rect 29972 1164 29978 1216
rect 30374 1164 30380 1216
rect 30432 1204 30438 1216
rect 30745 1207 30803 1213
rect 30745 1204 30757 1207
rect 30432 1176 30757 1204
rect 30432 1164 30438 1176
rect 30745 1173 30757 1176
rect 30791 1173 30803 1207
rect 30745 1167 30803 1173
rect 31570 1164 31576 1216
rect 31628 1164 31634 1216
rect 32490 1164 32496 1216
rect 32548 1164 32554 1216
rect 36078 1164 36084 1216
rect 36136 1164 36142 1216
rect 38010 1164 38016 1216
rect 38068 1164 38074 1216
rect 39301 1207 39359 1213
rect 39301 1173 39313 1207
rect 39347 1204 39359 1207
rect 39850 1204 39856 1216
rect 39347 1176 39856 1204
rect 39347 1173 39359 1176
rect 39301 1167 39359 1173
rect 39850 1164 39856 1176
rect 39908 1164 39914 1216
rect 40586 1164 40592 1216
rect 40644 1164 40650 1216
rect 41230 1164 41236 1216
rect 41288 1164 41294 1216
rect 41506 1164 41512 1216
rect 41564 1204 41570 1216
rect 41877 1207 41935 1213
rect 41877 1204 41889 1207
rect 41564 1176 41889 1204
rect 41564 1164 41570 1176
rect 41877 1173 41889 1176
rect 41923 1173 41935 1207
rect 41877 1167 41935 1173
rect 43070 1164 43076 1216
rect 43128 1164 43134 1216
rect 43824 1213 43852 1244
rect 46658 1232 46664 1284
rect 46716 1272 46722 1284
rect 46716 1244 48268 1272
rect 46716 1232 46722 1244
rect 43809 1207 43867 1213
rect 43809 1173 43821 1207
rect 43855 1173 43867 1207
rect 43809 1167 43867 1173
rect 45002 1164 45008 1216
rect 45060 1204 45066 1216
rect 45741 1207 45799 1213
rect 45741 1204 45753 1207
rect 45060 1176 45753 1204
rect 45060 1164 45066 1176
rect 45741 1173 45753 1176
rect 45787 1173 45799 1207
rect 45741 1167 45799 1173
rect 45830 1164 45836 1216
rect 45888 1204 45894 1216
rect 46385 1207 46443 1213
rect 46385 1204 46397 1207
rect 45888 1176 46397 1204
rect 45888 1164 45894 1176
rect 46385 1173 46397 1176
rect 46431 1173 46443 1207
rect 46385 1167 46443 1173
rect 46842 1164 46848 1216
rect 46900 1204 46906 1216
rect 48240 1213 48268 1244
rect 52914 1232 52920 1284
rect 52972 1272 52978 1284
rect 54297 1275 54355 1281
rect 54297 1272 54309 1275
rect 52972 1244 54309 1272
rect 52972 1232 52978 1244
rect 54297 1241 54309 1244
rect 54343 1241 54355 1275
rect 77312 1272 77340 1303
rect 77570 1300 77576 1352
rect 77628 1300 77634 1352
rect 79873 1343 79931 1349
rect 79873 1309 79885 1343
rect 79919 1340 79931 1343
rect 79962 1340 79968 1352
rect 79919 1312 79968 1340
rect 79919 1309 79931 1312
rect 79873 1303 79931 1309
rect 79962 1300 79968 1312
rect 80020 1300 80026 1352
rect 80149 1343 80207 1349
rect 80149 1309 80161 1343
rect 80195 1309 80207 1343
rect 80149 1303 80207 1309
rect 82449 1343 82507 1349
rect 82449 1309 82461 1343
rect 82495 1309 82507 1343
rect 82449 1303 82507 1309
rect 78582 1272 78588 1284
rect 77312 1244 78588 1272
rect 54297 1235 54355 1241
rect 78582 1232 78588 1244
rect 78640 1232 78646 1284
rect 47029 1207 47087 1213
rect 47029 1204 47041 1207
rect 46900 1176 47041 1204
rect 46900 1164 46906 1176
rect 47029 1173 47041 1176
rect 47075 1173 47087 1207
rect 47029 1167 47087 1173
rect 48225 1207 48283 1213
rect 48225 1173 48237 1207
rect 48271 1173 48283 1207
rect 48225 1167 48283 1173
rect 48866 1164 48872 1216
rect 48924 1204 48930 1216
rect 48961 1207 49019 1213
rect 48961 1204 48973 1207
rect 48924 1176 48973 1204
rect 48924 1164 48930 1176
rect 48961 1173 48973 1176
rect 49007 1173 49019 1207
rect 48961 1167 49019 1173
rect 49602 1164 49608 1216
rect 49660 1164 49666 1216
rect 50706 1164 50712 1216
rect 50764 1204 50770 1216
rect 50893 1207 50951 1213
rect 50893 1204 50905 1207
rect 50764 1176 50905 1204
rect 50764 1164 50770 1176
rect 50893 1173 50905 1176
rect 50939 1173 50951 1207
rect 50893 1167 50951 1173
rect 51534 1164 51540 1216
rect 51592 1164 51598 1216
rect 51994 1164 52000 1216
rect 52052 1204 52058 1216
rect 52181 1207 52239 1213
rect 52181 1204 52193 1207
rect 52052 1176 52193 1204
rect 52052 1164 52058 1176
rect 52181 1173 52193 1176
rect 52227 1173 52239 1207
rect 52181 1167 52239 1173
rect 53374 1164 53380 1216
rect 53432 1164 53438 1216
rect 56226 1164 56232 1216
rect 56284 1164 56290 1216
rect 57054 1164 57060 1216
rect 57112 1164 57118 1216
rect 58618 1164 58624 1216
rect 58676 1164 58682 1216
rect 60826 1164 60832 1216
rect 60884 1164 60890 1216
rect 61562 1164 61568 1216
rect 61620 1164 61626 1216
rect 62298 1164 62304 1216
rect 62356 1164 62362 1216
rect 63770 1164 63776 1216
rect 63828 1164 63834 1216
rect 64506 1164 64512 1216
rect 64564 1164 64570 1216
rect 66162 1164 66168 1216
rect 66220 1164 66226 1216
rect 80164 1204 80192 1303
rect 82464 1272 82492 1303
rect 82722 1300 82728 1352
rect 82780 1300 82786 1352
rect 85022 1300 85028 1352
rect 85080 1300 85086 1352
rect 85298 1300 85304 1352
rect 85356 1300 85362 1352
rect 86770 1300 86776 1352
rect 86828 1300 86834 1352
rect 87046 1300 87052 1352
rect 87104 1300 87110 1352
rect 88260 1349 88288 1380
rect 88518 1368 88524 1380
rect 88576 1408 88582 1420
rect 89530 1408 89536 1420
rect 88576 1380 89536 1408
rect 88576 1368 88582 1380
rect 88245 1343 88303 1349
rect 88245 1309 88257 1343
rect 88291 1309 88303 1343
rect 88245 1303 88303 1309
rect 88334 1300 88340 1352
rect 88392 1340 88398 1352
rect 88429 1343 88487 1349
rect 88429 1340 88441 1343
rect 88392 1312 88441 1340
rect 88392 1300 88398 1312
rect 88429 1309 88441 1312
rect 88475 1309 88487 1343
rect 88429 1303 88487 1309
rect 89070 1300 89076 1352
rect 89128 1300 89134 1352
rect 89180 1349 89208 1380
rect 89530 1368 89536 1380
rect 89588 1368 89594 1420
rect 98270 1368 98276 1420
rect 98328 1408 98334 1420
rect 98365 1411 98423 1417
rect 98365 1408 98377 1411
rect 98328 1380 98377 1408
rect 98328 1368 98334 1380
rect 98365 1377 98377 1380
rect 98411 1377 98423 1411
rect 98365 1371 98423 1377
rect 98472 1380 98684 1408
rect 89165 1343 89223 1349
rect 89165 1309 89177 1343
rect 89211 1309 89223 1343
rect 89165 1303 89223 1309
rect 89254 1300 89260 1352
rect 89312 1340 89318 1352
rect 89349 1343 89407 1349
rect 89349 1340 89361 1343
rect 89312 1312 89361 1340
rect 89312 1300 89318 1312
rect 89349 1309 89361 1312
rect 89395 1309 89407 1343
rect 89349 1303 89407 1309
rect 90450 1300 90456 1352
rect 90508 1300 90514 1352
rect 92014 1300 92020 1352
rect 92072 1300 92078 1352
rect 93302 1300 93308 1352
rect 93360 1300 93366 1352
rect 94866 1300 94872 1352
rect 94924 1300 94930 1352
rect 94958 1300 94964 1352
rect 95016 1300 95022 1352
rect 95881 1343 95939 1349
rect 95881 1309 95893 1343
rect 95927 1340 95939 1343
rect 96614 1340 96620 1352
rect 95927 1312 96620 1340
rect 95927 1309 95939 1312
rect 95881 1303 95939 1309
rect 96614 1300 96620 1312
rect 96672 1300 96678 1352
rect 96893 1343 96951 1349
rect 96893 1309 96905 1343
rect 96939 1340 96951 1343
rect 97166 1340 97172 1352
rect 96939 1312 97172 1340
rect 96939 1309 96951 1312
rect 96893 1303 96951 1309
rect 97166 1300 97172 1312
rect 97224 1300 97230 1352
rect 97629 1343 97687 1349
rect 97629 1309 97641 1343
rect 97675 1340 97687 1343
rect 98472 1340 98500 1380
rect 97675 1312 98500 1340
rect 97675 1309 97687 1312
rect 97629 1303 97687 1309
rect 98546 1300 98552 1352
rect 98604 1300 98610 1352
rect 98656 1340 98684 1380
rect 99558 1368 99564 1420
rect 99616 1408 99622 1420
rect 99929 1411 99987 1417
rect 99929 1408 99941 1411
rect 99616 1380 99941 1408
rect 99616 1368 99622 1380
rect 99929 1377 99941 1380
rect 99975 1377 99987 1411
rect 99929 1371 99987 1377
rect 100220 1380 100892 1408
rect 98733 1343 98791 1349
rect 98733 1340 98745 1343
rect 98656 1312 98745 1340
rect 98733 1309 98745 1312
rect 98779 1309 98791 1343
rect 98733 1303 98791 1309
rect 99285 1343 99343 1349
rect 99285 1309 99297 1343
rect 99331 1340 99343 1343
rect 99834 1340 99840 1352
rect 99331 1312 99840 1340
rect 99331 1309 99343 1312
rect 99285 1303 99343 1309
rect 99834 1300 99840 1312
rect 99892 1300 99898 1352
rect 100110 1300 100116 1352
rect 100168 1300 100174 1352
rect 84470 1272 84476 1284
rect 82464 1244 84476 1272
rect 84470 1232 84476 1244
rect 84528 1232 84534 1284
rect 100220 1272 100248 1380
rect 100297 1343 100355 1349
rect 100297 1309 100309 1343
rect 100343 1340 100355 1343
rect 100757 1343 100815 1349
rect 100757 1340 100769 1343
rect 100343 1312 100769 1340
rect 100343 1309 100355 1312
rect 100297 1303 100355 1309
rect 100757 1309 100769 1312
rect 100803 1309 100815 1343
rect 100864 1340 100892 1380
rect 103238 1368 103244 1420
rect 103296 1368 103302 1420
rect 109972 1380 110184 1408
rect 100864 1312 103836 1340
rect 100757 1303 100815 1309
rect 88352 1244 100248 1272
rect 88352 1204 88380 1244
rect 100570 1232 100576 1284
rect 100628 1272 100634 1284
rect 103808 1272 103836 1312
rect 103882 1300 103888 1352
rect 103940 1300 103946 1352
rect 104710 1300 104716 1352
rect 104768 1340 104774 1352
rect 104897 1343 104955 1349
rect 104897 1340 104909 1343
rect 104768 1312 104909 1340
rect 104768 1300 104774 1312
rect 104897 1309 104909 1312
rect 104943 1309 104955 1343
rect 104897 1303 104955 1309
rect 105630 1300 105636 1352
rect 105688 1300 105694 1352
rect 106182 1300 106188 1352
rect 106240 1340 106246 1352
rect 106369 1343 106427 1349
rect 106369 1340 106381 1343
rect 106240 1312 106381 1340
rect 106240 1300 106246 1312
rect 106369 1309 106381 1312
rect 106415 1309 106427 1343
rect 106369 1303 106427 1309
rect 107746 1300 107752 1352
rect 107804 1300 107810 1352
rect 108390 1300 108396 1352
rect 108448 1300 108454 1352
rect 109034 1300 109040 1352
rect 109092 1300 109098 1352
rect 109218 1300 109224 1352
rect 109276 1340 109282 1352
rect 109972 1340 110000 1380
rect 109276 1312 110000 1340
rect 109276 1300 109282 1312
rect 110046 1300 110052 1352
rect 110104 1300 110110 1352
rect 110156 1340 110184 1380
rect 110966 1368 110972 1420
rect 111024 1408 111030 1420
rect 149238 1408 149244 1420
rect 111024 1380 149244 1408
rect 111024 1368 111030 1380
rect 149238 1368 149244 1380
rect 149296 1368 149302 1420
rect 154132 1380 154988 1408
rect 110156 1312 110736 1340
rect 104250 1272 104256 1284
rect 100628 1244 103744 1272
rect 103808 1244 104256 1272
rect 100628 1232 100634 1244
rect 80164 1176 88380 1204
rect 90634 1164 90640 1216
rect 90692 1164 90698 1216
rect 92198 1164 92204 1216
rect 92256 1164 92262 1216
rect 93486 1164 93492 1216
rect 93544 1164 93550 1216
rect 96065 1207 96123 1213
rect 96065 1173 96077 1207
rect 96111 1204 96123 1207
rect 96522 1204 96528 1216
rect 96111 1176 96528 1204
rect 96111 1173 96123 1176
rect 96065 1167 96123 1173
rect 96522 1164 96528 1176
rect 96580 1164 96586 1216
rect 97074 1164 97080 1216
rect 97132 1164 97138 1216
rect 97813 1207 97871 1213
rect 97813 1173 97825 1207
rect 97859 1204 97871 1207
rect 98454 1204 98460 1216
rect 97859 1176 98460 1204
rect 97859 1173 97871 1176
rect 97813 1167 97871 1173
rect 98454 1164 98460 1176
rect 98512 1164 98518 1216
rect 100018 1164 100024 1216
rect 100076 1204 100082 1216
rect 103716 1213 103744 1244
rect 104250 1232 104256 1244
rect 104308 1232 104314 1284
rect 104802 1232 104808 1284
rect 104860 1272 104866 1284
rect 104860 1244 106228 1272
rect 104860 1232 104866 1244
rect 100941 1207 100999 1213
rect 100941 1204 100953 1207
rect 100076 1176 100953 1204
rect 100076 1164 100082 1176
rect 100941 1173 100953 1176
rect 100987 1173 100999 1207
rect 100941 1167 100999 1173
rect 103701 1207 103759 1213
rect 103701 1173 103713 1207
rect 103747 1173 103759 1207
rect 103701 1167 103759 1173
rect 104618 1164 104624 1216
rect 104676 1204 104682 1216
rect 104713 1207 104771 1213
rect 104713 1204 104725 1207
rect 104676 1176 104725 1204
rect 104676 1164 104682 1176
rect 104713 1173 104725 1176
rect 104759 1173 104771 1207
rect 104713 1167 104771 1173
rect 105446 1164 105452 1216
rect 105504 1164 105510 1216
rect 106200 1213 106228 1244
rect 107470 1232 107476 1284
rect 107528 1272 107534 1284
rect 107528 1244 107700 1272
rect 107528 1232 107534 1244
rect 106185 1207 106243 1213
rect 106185 1173 106197 1207
rect 106231 1173 106243 1207
rect 106185 1167 106243 1173
rect 106274 1164 106280 1216
rect 106332 1204 106338 1216
rect 107565 1207 107623 1213
rect 107565 1204 107577 1207
rect 106332 1176 107577 1204
rect 106332 1164 106338 1176
rect 107565 1173 107577 1176
rect 107611 1173 107623 1207
rect 107672 1204 107700 1244
rect 108114 1232 108120 1284
rect 108172 1272 108178 1284
rect 110708 1272 110736 1312
rect 110782 1300 110788 1352
rect 110840 1300 110846 1352
rect 111518 1300 111524 1352
rect 111576 1300 111582 1352
rect 112898 1300 112904 1352
rect 112956 1300 112962 1352
rect 113082 1300 113088 1352
rect 113140 1340 113146 1352
rect 113140 1312 113496 1340
rect 113140 1300 113146 1312
rect 108172 1244 110644 1272
rect 110708 1244 112852 1272
rect 108172 1232 108178 1244
rect 108209 1207 108267 1213
rect 108209 1204 108221 1207
rect 107672 1176 108221 1204
rect 107565 1167 107623 1173
rect 108209 1173 108221 1176
rect 108255 1173 108267 1207
rect 108209 1167 108267 1173
rect 108850 1164 108856 1216
rect 108908 1164 108914 1216
rect 109862 1164 109868 1216
rect 109920 1164 109926 1216
rect 110616 1213 110644 1244
rect 110601 1207 110659 1213
rect 110601 1173 110613 1207
rect 110647 1173 110659 1207
rect 110601 1167 110659 1173
rect 111334 1164 111340 1216
rect 111392 1164 111398 1216
rect 112714 1164 112720 1216
rect 112772 1164 112778 1216
rect 112824 1204 112852 1244
rect 112990 1232 112996 1284
rect 113048 1272 113054 1284
rect 113358 1272 113364 1284
rect 113048 1244 113364 1272
rect 113048 1232 113054 1244
rect 113358 1232 113364 1244
rect 113416 1232 113422 1284
rect 113468 1272 113496 1312
rect 113542 1300 113548 1352
rect 113600 1300 113606 1352
rect 113634 1300 113640 1352
rect 113692 1340 113698 1352
rect 113692 1312 113772 1340
rect 113692 1300 113698 1312
rect 113744 1272 113772 1312
rect 114186 1300 114192 1352
rect 114244 1300 114250 1352
rect 115198 1300 115204 1352
rect 115256 1300 115262 1352
rect 115750 1300 115756 1352
rect 115808 1340 115814 1352
rect 115937 1343 115995 1349
rect 115937 1340 115949 1343
rect 115808 1312 115949 1340
rect 115808 1300 115814 1312
rect 115937 1309 115949 1312
rect 115983 1309 115995 1343
rect 115937 1303 115995 1309
rect 116670 1300 116676 1352
rect 116728 1300 116734 1352
rect 118050 1300 118056 1352
rect 118108 1300 118114 1352
rect 118694 1300 118700 1352
rect 118752 1300 118758 1352
rect 119338 1300 119344 1352
rect 119396 1300 119402 1352
rect 120350 1300 120356 1352
rect 120408 1300 120414 1352
rect 121086 1300 121092 1352
rect 121144 1300 121150 1352
rect 121178 1300 121184 1352
rect 121236 1340 121242 1352
rect 121641 1343 121699 1349
rect 121641 1340 121653 1343
rect 121236 1312 121653 1340
rect 121236 1300 121242 1312
rect 121641 1309 121653 1312
rect 121687 1309 121699 1343
rect 121641 1303 121699 1309
rect 122926 1300 122932 1352
rect 122984 1300 122990 1352
rect 123754 1300 123760 1352
rect 123812 1300 123818 1352
rect 125410 1300 125416 1352
rect 125468 1300 125474 1352
rect 126793 1343 126851 1349
rect 126793 1309 126805 1343
rect 126839 1340 126851 1343
rect 127066 1340 127072 1352
rect 126839 1312 127072 1340
rect 126839 1309 126851 1312
rect 126793 1303 126851 1309
rect 127066 1300 127072 1312
rect 127124 1300 127130 1352
rect 128262 1300 128268 1352
rect 128320 1300 128326 1352
rect 128446 1300 128452 1352
rect 128504 1300 128510 1352
rect 128630 1300 128636 1352
rect 128688 1300 128694 1352
rect 129090 1300 129096 1352
rect 129148 1300 129154 1352
rect 130654 1300 130660 1352
rect 130712 1300 130718 1352
rect 131945 1343 132003 1349
rect 131945 1309 131957 1343
rect 131991 1340 132003 1343
rect 132586 1340 132592 1352
rect 131991 1312 132592 1340
rect 131991 1309 132003 1312
rect 131945 1303 132003 1309
rect 132586 1300 132592 1312
rect 132644 1300 132650 1352
rect 132770 1300 132776 1352
rect 132828 1340 132834 1352
rect 132957 1343 133015 1349
rect 132957 1340 132969 1343
rect 132828 1312 132969 1340
rect 132828 1300 132834 1312
rect 132957 1309 132969 1312
rect 133003 1309 133015 1343
rect 132957 1303 133015 1309
rect 133138 1300 133144 1352
rect 133196 1300 133202 1352
rect 133874 1300 133880 1352
rect 133932 1340 133938 1352
rect 133969 1343 134027 1349
rect 133969 1340 133981 1343
rect 133932 1312 133981 1340
rect 133932 1300 133938 1312
rect 133969 1309 133981 1312
rect 134015 1309 134027 1343
rect 133969 1303 134027 1309
rect 134058 1300 134064 1352
rect 134116 1340 134122 1352
rect 134153 1343 134211 1349
rect 134153 1340 134165 1343
rect 134116 1312 134165 1340
rect 134116 1300 134122 1312
rect 134153 1309 134165 1312
rect 134199 1309 134211 1343
rect 134153 1303 134211 1309
rect 138750 1300 138756 1352
rect 138808 1300 138814 1352
rect 138842 1300 138848 1352
rect 138900 1340 138906 1352
rect 139397 1343 139455 1349
rect 139397 1340 139409 1343
rect 138900 1312 139409 1340
rect 138900 1300 138906 1312
rect 139397 1309 139409 1312
rect 139443 1309 139455 1343
rect 139397 1303 139455 1309
rect 140682 1300 140688 1352
rect 140740 1300 140746 1352
rect 140774 1300 140780 1352
rect 140832 1340 140838 1352
rect 141329 1343 141387 1349
rect 141329 1340 141341 1343
rect 140832 1312 141341 1340
rect 140832 1300 140838 1312
rect 141329 1309 141341 1312
rect 141375 1309 141387 1343
rect 141329 1303 141387 1309
rect 141970 1300 141976 1352
rect 142028 1300 142034 1352
rect 142062 1300 142068 1352
rect 142120 1340 142126 1352
rect 143261 1343 143319 1349
rect 143261 1340 143273 1343
rect 142120 1312 143273 1340
rect 142120 1300 142126 1312
rect 143261 1309 143273 1312
rect 143307 1309 143319 1343
rect 143261 1303 143319 1309
rect 143534 1300 143540 1352
rect 143592 1340 143598 1352
rect 143905 1343 143963 1349
rect 143905 1340 143917 1343
rect 143592 1312 143917 1340
rect 143592 1300 143598 1312
rect 143905 1309 143917 1312
rect 143951 1309 143963 1343
rect 143905 1303 143963 1309
rect 144546 1300 144552 1352
rect 144604 1300 144610 1352
rect 145834 1300 145840 1352
rect 145892 1300 145898 1352
rect 146202 1300 146208 1352
rect 146260 1340 146266 1352
rect 146481 1343 146539 1349
rect 146481 1340 146493 1343
rect 146260 1312 146493 1340
rect 146260 1300 146266 1312
rect 146481 1309 146493 1312
rect 146527 1309 146539 1343
rect 146481 1303 146539 1309
rect 147122 1300 147128 1352
rect 147180 1300 147186 1352
rect 148410 1300 148416 1352
rect 148468 1300 148474 1352
rect 148502 1300 148508 1352
rect 148560 1340 148566 1352
rect 149057 1343 149115 1349
rect 149057 1340 149069 1343
rect 148560 1312 149069 1340
rect 148560 1300 148566 1312
rect 149057 1309 149069 1312
rect 149103 1309 149115 1343
rect 149057 1303 149115 1309
rect 149698 1300 149704 1352
rect 149756 1300 149762 1352
rect 150986 1300 150992 1352
rect 151044 1300 151050 1352
rect 151630 1300 151636 1352
rect 151688 1300 151694 1352
rect 152274 1300 152280 1352
rect 152332 1300 152338 1352
rect 153194 1300 153200 1352
rect 153252 1340 153258 1352
rect 153565 1343 153623 1349
rect 153565 1340 153577 1343
rect 153252 1312 153577 1340
rect 153252 1300 153258 1312
rect 153565 1309 153577 1312
rect 153611 1309 153623 1343
rect 154132 1340 154160 1380
rect 153565 1303 153623 1309
rect 153948 1312 154160 1340
rect 113468 1244 113588 1272
rect 113744 1244 115796 1272
rect 113266 1204 113272 1216
rect 112824 1176 113272 1204
rect 113266 1164 113272 1176
rect 113324 1164 113330 1216
rect 113560 1204 113588 1244
rect 114005 1207 114063 1213
rect 114005 1204 114017 1207
rect 113560 1176 114017 1204
rect 114005 1173 114017 1176
rect 114051 1173 114063 1207
rect 114005 1167 114063 1173
rect 115014 1164 115020 1216
rect 115072 1164 115078 1216
rect 115768 1213 115796 1244
rect 123570 1232 123576 1284
rect 123628 1272 123634 1284
rect 148778 1272 148784 1284
rect 123628 1244 148784 1272
rect 123628 1232 123634 1244
rect 148778 1232 148784 1244
rect 148836 1232 148842 1284
rect 150618 1272 150624 1284
rect 148888 1244 150624 1272
rect 115753 1207 115811 1213
rect 115753 1173 115765 1207
rect 115799 1173 115811 1207
rect 115753 1167 115811 1173
rect 115842 1164 115848 1216
rect 115900 1204 115906 1216
rect 116489 1207 116547 1213
rect 116489 1204 116501 1207
rect 115900 1176 116501 1204
rect 115900 1164 115906 1176
rect 116489 1173 116501 1176
rect 116535 1173 116547 1207
rect 116489 1167 116547 1173
rect 117222 1164 117228 1216
rect 117280 1204 117286 1216
rect 117869 1207 117927 1213
rect 117869 1204 117881 1207
rect 117280 1176 117881 1204
rect 117280 1164 117286 1176
rect 117869 1173 117881 1176
rect 117915 1173 117927 1207
rect 117869 1167 117927 1173
rect 118510 1164 118516 1216
rect 118568 1164 118574 1216
rect 119157 1207 119215 1213
rect 119157 1173 119169 1207
rect 119203 1204 119215 1207
rect 119246 1204 119252 1216
rect 119203 1176 119252 1204
rect 119203 1173 119215 1176
rect 119157 1167 119215 1173
rect 119246 1164 119252 1176
rect 119304 1164 119310 1216
rect 120166 1164 120172 1216
rect 120224 1164 120230 1216
rect 120810 1164 120816 1216
rect 120868 1204 120874 1216
rect 120905 1207 120963 1213
rect 120905 1204 120917 1207
rect 120868 1176 120917 1204
rect 120868 1164 120874 1176
rect 120905 1173 120917 1176
rect 120951 1173 120963 1207
rect 120905 1167 120963 1173
rect 121822 1164 121828 1216
rect 121880 1164 121886 1216
rect 123110 1164 123116 1216
rect 123168 1164 123174 1216
rect 123938 1164 123944 1216
rect 123996 1164 124002 1216
rect 125318 1164 125324 1216
rect 125376 1204 125382 1216
rect 125597 1207 125655 1213
rect 125597 1204 125609 1207
rect 125376 1176 125609 1204
rect 125376 1164 125382 1176
rect 125597 1173 125609 1176
rect 125643 1173 125655 1207
rect 125597 1167 125655 1173
rect 126790 1164 126796 1216
rect 126848 1204 126854 1216
rect 126977 1207 127035 1213
rect 126977 1204 126989 1207
rect 126848 1176 126989 1204
rect 126848 1164 126854 1176
rect 126977 1173 126989 1176
rect 127023 1173 127035 1207
rect 126977 1167 127035 1173
rect 129274 1164 129280 1216
rect 129332 1164 129338 1216
rect 130838 1164 130844 1216
rect 130896 1164 130902 1216
rect 132126 1164 132132 1216
rect 132184 1164 132190 1216
rect 137922 1164 137928 1216
rect 137980 1204 137986 1216
rect 138569 1207 138627 1213
rect 138569 1204 138581 1207
rect 137980 1176 138581 1204
rect 137980 1164 137986 1176
rect 138569 1173 138581 1176
rect 138615 1173 138627 1207
rect 138569 1167 138627 1173
rect 140866 1164 140872 1216
rect 140924 1204 140930 1216
rect 141145 1207 141203 1213
rect 141145 1204 141157 1207
rect 140924 1176 141157 1204
rect 140924 1164 140930 1176
rect 141145 1173 141157 1176
rect 141191 1173 141203 1207
rect 141145 1167 141203 1173
rect 141789 1207 141847 1213
rect 141789 1173 141801 1207
rect 141835 1204 141847 1207
rect 141878 1204 141884 1216
rect 141835 1176 141884 1204
rect 141835 1173 141847 1176
rect 141789 1167 141847 1173
rect 141878 1164 141884 1176
rect 141936 1164 141942 1216
rect 143074 1164 143080 1216
rect 143132 1164 143138 1216
rect 143721 1207 143779 1213
rect 143721 1173 143733 1207
rect 143767 1204 143779 1207
rect 143810 1204 143816 1216
rect 143767 1176 143816 1204
rect 143767 1173 143779 1176
rect 143721 1167 143779 1173
rect 143810 1164 143816 1176
rect 143868 1164 143874 1216
rect 144362 1164 144368 1216
rect 144420 1164 144426 1216
rect 145650 1164 145656 1216
rect 145708 1164 145714 1216
rect 146110 1164 146116 1216
rect 146168 1204 146174 1216
rect 146297 1207 146355 1213
rect 146297 1204 146309 1207
rect 146168 1176 146309 1204
rect 146168 1164 146174 1176
rect 146297 1173 146309 1176
rect 146343 1173 146355 1207
rect 146297 1167 146355 1173
rect 146386 1164 146392 1216
rect 146444 1204 146450 1216
rect 146941 1207 146999 1213
rect 146941 1204 146953 1207
rect 146444 1176 146953 1204
rect 146444 1164 146450 1176
rect 146941 1173 146953 1176
rect 146987 1173 146999 1207
rect 146941 1167 146999 1173
rect 148226 1164 148232 1216
rect 148284 1164 148290 1216
rect 148888 1213 148916 1244
rect 150618 1232 150624 1244
rect 150676 1232 150682 1284
rect 153286 1272 153292 1284
rect 151464 1244 153292 1272
rect 148873 1207 148931 1213
rect 148873 1173 148885 1207
rect 148919 1173 148931 1207
rect 148873 1167 148931 1173
rect 149517 1207 149575 1213
rect 149517 1173 149529 1207
rect 149563 1204 149575 1207
rect 150710 1204 150716 1216
rect 149563 1176 150716 1204
rect 149563 1173 149575 1176
rect 149517 1167 149575 1173
rect 150710 1164 150716 1176
rect 150768 1164 150774 1216
rect 150805 1207 150863 1213
rect 150805 1173 150817 1207
rect 150851 1204 150863 1207
rect 150894 1204 150900 1216
rect 150851 1176 150900 1204
rect 150851 1173 150863 1176
rect 150805 1167 150863 1173
rect 150894 1164 150900 1176
rect 150952 1164 150958 1216
rect 151464 1213 151492 1244
rect 153286 1232 153292 1244
rect 153344 1232 153350 1284
rect 151449 1207 151507 1213
rect 151449 1173 151461 1207
rect 151495 1173 151507 1207
rect 151449 1167 151507 1173
rect 152090 1164 152096 1216
rect 152148 1164 152154 1216
rect 153381 1207 153439 1213
rect 153381 1173 153393 1207
rect 153427 1204 153439 1207
rect 153948 1204 153976 1312
rect 154206 1300 154212 1352
rect 154264 1300 154270 1352
rect 154574 1300 154580 1352
rect 154632 1340 154638 1352
rect 154853 1343 154911 1349
rect 154853 1340 154865 1343
rect 154632 1312 154865 1340
rect 154632 1300 154638 1312
rect 154853 1309 154865 1312
rect 154899 1309 154911 1343
rect 154960 1340 154988 1380
rect 156506 1368 156512 1420
rect 156564 1408 156570 1420
rect 157058 1408 157064 1420
rect 156564 1380 157064 1408
rect 156564 1368 156570 1380
rect 157058 1368 157064 1380
rect 157116 1408 157122 1420
rect 157245 1411 157303 1417
rect 157245 1408 157257 1411
rect 157116 1380 157257 1408
rect 157116 1368 157122 1380
rect 157245 1377 157257 1380
rect 157291 1377 157303 1411
rect 157245 1371 157303 1377
rect 158162 1368 158168 1420
rect 158220 1408 158226 1420
rect 158533 1411 158591 1417
rect 158533 1408 158545 1411
rect 158220 1380 158545 1408
rect 158220 1368 158226 1380
rect 158533 1377 158545 1380
rect 158579 1377 158591 1411
rect 158533 1371 158591 1377
rect 159082 1368 159088 1420
rect 159140 1408 159146 1420
rect 159361 1411 159419 1417
rect 159361 1408 159373 1411
rect 159140 1380 159373 1408
rect 159140 1368 159146 1380
rect 159361 1377 159373 1380
rect 159407 1377 159419 1411
rect 160370 1408 160376 1420
rect 159361 1371 159419 1377
rect 160112 1380 160376 1408
rect 156138 1340 156144 1352
rect 154960 1312 156144 1340
rect 154853 1303 154911 1309
rect 156138 1300 156144 1312
rect 156196 1300 156202 1352
rect 156417 1343 156475 1349
rect 156417 1309 156429 1343
rect 156463 1309 156475 1343
rect 156417 1303 156475 1309
rect 156601 1343 156659 1349
rect 156601 1309 156613 1343
rect 156647 1309 156659 1343
rect 156601 1303 156659 1309
rect 157429 1343 157487 1349
rect 157429 1309 157441 1343
rect 157475 1309 157487 1343
rect 157429 1303 157487 1309
rect 158717 1343 158775 1349
rect 158717 1309 158729 1343
rect 158763 1340 158775 1343
rect 159266 1340 159272 1352
rect 158763 1312 159272 1340
rect 158763 1309 158775 1312
rect 158717 1303 158775 1309
rect 156230 1272 156236 1284
rect 154040 1244 156236 1272
rect 154040 1213 154068 1244
rect 156230 1232 156236 1244
rect 156288 1232 156294 1284
rect 153427 1176 153976 1204
rect 154025 1207 154083 1213
rect 153427 1173 153439 1176
rect 153381 1167 153439 1173
rect 154025 1173 154037 1207
rect 154071 1173 154083 1207
rect 154025 1167 154083 1173
rect 154669 1207 154727 1213
rect 154669 1173 154681 1207
rect 154715 1204 154727 1207
rect 156046 1204 156052 1216
rect 154715 1176 156052 1204
rect 154715 1173 154727 1176
rect 154669 1167 154727 1173
rect 156046 1164 156052 1176
rect 156104 1164 156110 1216
rect 156432 1204 156460 1303
rect 156616 1272 156644 1303
rect 157444 1272 157472 1303
rect 158732 1272 158760 1303
rect 159266 1300 159272 1312
rect 159324 1340 159330 1352
rect 159545 1343 159603 1349
rect 159545 1340 159557 1343
rect 159324 1312 159557 1340
rect 159324 1300 159330 1312
rect 159545 1309 159557 1312
rect 159591 1309 159603 1343
rect 159545 1303 159603 1309
rect 159729 1343 159787 1349
rect 159729 1309 159741 1343
rect 159775 1340 159787 1343
rect 160112 1340 160140 1380
rect 160370 1368 160376 1380
rect 160428 1368 160434 1420
rect 163685 1411 163743 1417
rect 163685 1377 163697 1411
rect 163731 1408 163743 1411
rect 164142 1408 164148 1420
rect 163731 1380 164148 1408
rect 163731 1377 163743 1380
rect 163685 1371 163743 1377
rect 164142 1368 164148 1380
rect 164200 1368 164206 1420
rect 166997 1411 167055 1417
rect 166997 1377 167009 1411
rect 167043 1408 167055 1411
rect 168098 1408 168104 1420
rect 167043 1380 168104 1408
rect 167043 1377 167055 1380
rect 166997 1371 167055 1377
rect 168098 1368 168104 1380
rect 168156 1368 168162 1420
rect 171686 1368 171692 1420
rect 171744 1368 171750 1420
rect 190914 1368 190920 1420
rect 190972 1408 190978 1420
rect 201221 1411 201279 1417
rect 190972 1380 191236 1408
rect 190972 1368 190978 1380
rect 159775 1312 160140 1340
rect 159775 1309 159787 1312
rect 159729 1303 159787 1309
rect 160186 1300 160192 1352
rect 160244 1300 160250 1352
rect 161109 1343 161167 1349
rect 161109 1309 161121 1343
rect 161155 1340 161167 1343
rect 161474 1340 161480 1352
rect 161155 1312 161480 1340
rect 161155 1309 161167 1312
rect 161109 1303 161167 1309
rect 161474 1300 161480 1312
rect 161532 1300 161538 1352
rect 162305 1343 162363 1349
rect 162305 1309 162317 1343
rect 162351 1340 162363 1343
rect 163130 1340 163136 1352
rect 162351 1312 163136 1340
rect 162351 1309 162363 1312
rect 162305 1303 162363 1309
rect 163130 1300 163136 1312
rect 163188 1300 163194 1352
rect 163774 1300 163780 1352
rect 163832 1340 163838 1352
rect 163869 1343 163927 1349
rect 163869 1340 163881 1343
rect 163832 1312 163881 1340
rect 163832 1300 163838 1312
rect 163869 1309 163881 1312
rect 163915 1309 163927 1343
rect 163869 1303 163927 1309
rect 164053 1343 164111 1349
rect 164053 1309 164065 1343
rect 164099 1340 164111 1343
rect 164418 1340 164424 1352
rect 164099 1312 164424 1340
rect 164099 1309 164111 1312
rect 164053 1303 164111 1309
rect 164418 1300 164424 1312
rect 164476 1300 164482 1352
rect 164510 1300 164516 1352
rect 164568 1300 164574 1352
rect 167178 1300 167184 1352
rect 167236 1300 167242 1352
rect 167365 1343 167423 1349
rect 167365 1309 167377 1343
rect 167411 1340 167423 1343
rect 167825 1343 167883 1349
rect 167825 1340 167837 1343
rect 167411 1312 167837 1340
rect 167411 1309 167423 1312
rect 167365 1303 167423 1309
rect 167825 1309 167837 1312
rect 167871 1309 167883 1343
rect 167825 1303 167883 1309
rect 168006 1300 168012 1352
rect 168064 1340 168070 1352
rect 168837 1343 168895 1349
rect 168837 1340 168849 1343
rect 168064 1312 168849 1340
rect 168064 1300 168070 1312
rect 168837 1309 168849 1312
rect 168883 1309 168895 1343
rect 168837 1303 168895 1309
rect 172238 1300 172244 1352
rect 172296 1300 172302 1352
rect 172514 1300 172520 1352
rect 172572 1300 172578 1352
rect 173802 1300 173808 1352
rect 173860 1340 173866 1352
rect 173989 1343 174047 1349
rect 173989 1340 174001 1343
rect 173860 1312 174001 1340
rect 173860 1300 173866 1312
rect 173989 1309 174001 1312
rect 174035 1309 174047 1343
rect 173989 1303 174047 1309
rect 174262 1300 174268 1352
rect 174320 1300 174326 1352
rect 175182 1300 175188 1352
rect 175240 1340 175246 1352
rect 176565 1343 176623 1349
rect 176565 1340 176577 1343
rect 175240 1312 176577 1340
rect 175240 1300 175246 1312
rect 176565 1309 176577 1312
rect 176611 1309 176623 1343
rect 176565 1303 176623 1309
rect 176838 1300 176844 1352
rect 176896 1300 176902 1352
rect 178402 1300 178408 1352
rect 178460 1340 178466 1352
rect 179141 1343 179199 1349
rect 179141 1340 179153 1343
rect 178460 1312 179153 1340
rect 178460 1300 178466 1312
rect 179141 1309 179153 1312
rect 179187 1309 179199 1343
rect 179141 1303 179199 1309
rect 179414 1300 179420 1352
rect 179472 1300 179478 1352
rect 182542 1300 182548 1352
rect 182600 1300 182606 1352
rect 182818 1300 182824 1352
rect 182876 1300 182882 1352
rect 184290 1300 184296 1352
rect 184348 1300 184354 1352
rect 184566 1300 184572 1352
rect 184624 1300 184630 1352
rect 185578 1300 185584 1352
rect 185636 1340 185642 1352
rect 186869 1343 186927 1349
rect 186869 1340 186881 1343
rect 185636 1312 186881 1340
rect 185636 1300 185642 1312
rect 186869 1309 186881 1312
rect 186915 1309 186927 1343
rect 186869 1303 186927 1309
rect 187142 1300 187148 1352
rect 187200 1300 187206 1352
rect 188522 1300 188528 1352
rect 188580 1340 188586 1352
rect 189445 1343 189503 1349
rect 189445 1340 189457 1343
rect 188580 1312 189457 1340
rect 188580 1300 188586 1312
rect 189445 1309 189457 1312
rect 189491 1309 189503 1343
rect 189445 1303 189503 1309
rect 189718 1300 189724 1352
rect 189776 1300 189782 1352
rect 191098 1300 191104 1352
rect 191156 1300 191162 1352
rect 191208 1349 191236 1380
rect 201221 1377 201233 1411
rect 201267 1408 201279 1411
rect 202046 1408 202052 1420
rect 201267 1380 202052 1408
rect 201267 1377 201279 1380
rect 201221 1371 201279 1377
rect 202046 1368 202052 1380
rect 202104 1368 202110 1420
rect 202322 1368 202328 1420
rect 202380 1368 202386 1420
rect 205818 1368 205824 1420
rect 205876 1368 205882 1420
rect 191193 1343 191251 1349
rect 191193 1309 191205 1343
rect 191239 1309 191251 1343
rect 191193 1303 191251 1309
rect 192481 1343 192539 1349
rect 192481 1309 192493 1343
rect 192527 1340 192539 1343
rect 193214 1340 193220 1352
rect 192527 1312 193220 1340
rect 192527 1309 192539 1312
rect 192481 1303 192539 1309
rect 193214 1300 193220 1312
rect 193272 1300 193278 1352
rect 193306 1300 193312 1352
rect 193364 1300 193370 1352
rect 194594 1300 194600 1352
rect 194652 1300 194658 1352
rect 195609 1343 195667 1349
rect 195609 1309 195621 1343
rect 195655 1340 195667 1343
rect 196526 1340 196532 1352
rect 195655 1312 196532 1340
rect 195655 1309 195667 1312
rect 195609 1303 195667 1309
rect 196526 1300 196532 1312
rect 196584 1300 196590 1352
rect 197173 1343 197231 1349
rect 197173 1309 197185 1343
rect 197219 1340 197231 1343
rect 197446 1340 197452 1352
rect 197219 1312 197452 1340
rect 197219 1309 197231 1312
rect 197173 1303 197231 1309
rect 197446 1300 197452 1312
rect 197504 1300 197510 1352
rect 197906 1300 197912 1352
rect 197964 1300 197970 1352
rect 199746 1300 199752 1352
rect 199804 1300 199810 1352
rect 200485 1343 200543 1349
rect 200485 1309 200497 1343
rect 200531 1309 200543 1343
rect 200485 1303 200543 1309
rect 156616 1244 158760 1272
rect 158806 1232 158812 1284
rect 158864 1272 158870 1284
rect 158864 1244 160416 1272
rect 158864 1232 158870 1244
rect 156966 1204 156972 1216
rect 156432 1176 156972 1204
rect 156966 1164 156972 1176
rect 157024 1164 157030 1216
rect 157702 1164 157708 1216
rect 157760 1204 157766 1216
rect 160388 1213 160416 1244
rect 161382 1232 161388 1284
rect 161440 1272 161446 1284
rect 179506 1272 179512 1284
rect 161440 1244 179512 1272
rect 161440 1232 161446 1244
rect 179506 1232 179512 1244
rect 179564 1232 179570 1284
rect 180518 1232 180524 1284
rect 180576 1232 180582 1284
rect 181806 1232 181812 1284
rect 181864 1232 181870 1284
rect 197262 1232 197268 1284
rect 197320 1272 197326 1284
rect 200500 1272 200528 1303
rect 201310 1300 201316 1352
rect 201368 1340 201374 1352
rect 201405 1343 201463 1349
rect 201405 1340 201417 1343
rect 201368 1312 201417 1340
rect 201368 1300 201374 1312
rect 201405 1309 201417 1312
rect 201451 1340 201463 1343
rect 202509 1343 202567 1349
rect 202509 1340 202521 1343
rect 201451 1312 202521 1340
rect 201451 1309 201463 1312
rect 201405 1303 201463 1309
rect 202509 1309 202521 1312
rect 202555 1309 202567 1343
rect 202509 1303 202567 1309
rect 202693 1343 202751 1349
rect 202693 1309 202705 1343
rect 202739 1340 202751 1343
rect 203153 1343 203211 1349
rect 203153 1340 203165 1343
rect 202739 1312 203165 1340
rect 202739 1309 202751 1312
rect 202693 1303 202751 1309
rect 203153 1309 203165 1312
rect 203199 1309 203211 1343
rect 203153 1303 203211 1309
rect 206554 1300 206560 1352
rect 206612 1300 206618 1352
rect 207658 1300 207664 1352
rect 207716 1300 207722 1352
rect 208302 1300 208308 1352
rect 208360 1300 208366 1352
rect 208946 1300 208952 1352
rect 209004 1300 209010 1352
rect 209774 1300 209780 1352
rect 209832 1340 209838 1352
rect 210237 1343 210295 1349
rect 210237 1340 210249 1343
rect 209832 1312 210249 1340
rect 209832 1300 209838 1312
rect 210237 1309 210249 1312
rect 210283 1309 210295 1343
rect 210237 1303 210295 1309
rect 210878 1300 210884 1352
rect 210936 1300 210942 1352
rect 211522 1300 211528 1352
rect 211580 1300 211586 1352
rect 212258 1300 212264 1352
rect 212316 1340 212322 1352
rect 212813 1343 212871 1349
rect 212813 1340 212825 1343
rect 212316 1312 212825 1340
rect 212316 1300 212322 1312
rect 212813 1309 212825 1312
rect 212859 1309 212871 1343
rect 212813 1303 212871 1309
rect 201678 1272 201684 1284
rect 197320 1244 198136 1272
rect 200500 1244 201684 1272
rect 197320 1232 197326 1244
rect 158901 1207 158959 1213
rect 158901 1204 158913 1207
rect 157760 1176 158913 1204
rect 157760 1164 157766 1176
rect 158901 1173 158913 1176
rect 158947 1173 158959 1207
rect 158901 1167 158959 1173
rect 160373 1207 160431 1213
rect 160373 1173 160385 1207
rect 160419 1173 160431 1207
rect 160373 1167 160431 1173
rect 161290 1164 161296 1216
rect 161348 1164 161354 1216
rect 162486 1164 162492 1216
rect 162544 1164 162550 1216
rect 164694 1164 164700 1216
rect 164752 1164 164758 1216
rect 168006 1164 168012 1216
rect 168064 1164 168070 1216
rect 169018 1164 169024 1216
rect 169076 1164 169082 1216
rect 181898 1164 181904 1216
rect 181956 1164 181962 1216
rect 192662 1164 192668 1216
rect 192720 1164 192726 1216
rect 192938 1164 192944 1216
rect 192996 1204 193002 1216
rect 193493 1207 193551 1213
rect 193493 1204 193505 1207
rect 192996 1176 193505 1204
rect 192996 1164 193002 1176
rect 193493 1173 193505 1176
rect 193539 1173 193551 1207
rect 193493 1167 193551 1173
rect 193674 1164 193680 1216
rect 193732 1204 193738 1216
rect 194781 1207 194839 1213
rect 194781 1204 194793 1207
rect 193732 1176 194793 1204
rect 193732 1164 193738 1176
rect 194781 1173 194793 1176
rect 194827 1173 194839 1207
rect 194781 1167 194839 1173
rect 195790 1164 195796 1216
rect 195848 1164 195854 1216
rect 196618 1164 196624 1216
rect 196676 1204 196682 1216
rect 198108 1213 198136 1244
rect 201678 1232 201684 1244
rect 201736 1232 201742 1284
rect 209958 1272 209964 1284
rect 208136 1244 209964 1272
rect 197357 1207 197415 1213
rect 197357 1204 197369 1207
rect 196676 1176 197369 1204
rect 196676 1164 196682 1176
rect 197357 1173 197369 1176
rect 197403 1173 197415 1207
rect 197357 1167 197415 1173
rect 198093 1207 198151 1213
rect 198093 1173 198105 1207
rect 198139 1173 198151 1207
rect 198093 1167 198151 1173
rect 199930 1164 199936 1216
rect 199988 1164 199994 1216
rect 200666 1164 200672 1216
rect 200724 1164 200730 1216
rect 201218 1164 201224 1216
rect 201276 1204 201282 1216
rect 201589 1207 201647 1213
rect 201589 1204 201601 1207
rect 201276 1176 201601 1204
rect 201276 1164 201282 1176
rect 201589 1173 201601 1176
rect 201635 1173 201647 1207
rect 201589 1167 201647 1173
rect 203334 1164 203340 1216
rect 203392 1164 203398 1216
rect 206370 1164 206376 1216
rect 206428 1164 206434 1216
rect 207474 1164 207480 1216
rect 207532 1164 207538 1216
rect 208136 1213 208164 1244
rect 209958 1232 209964 1244
rect 210016 1232 210022 1284
rect 212534 1272 212540 1284
rect 211264 1244 212540 1272
rect 208121 1207 208179 1213
rect 208121 1173 208133 1207
rect 208167 1173 208179 1207
rect 208121 1167 208179 1173
rect 208765 1207 208823 1213
rect 208765 1173 208777 1207
rect 208811 1204 208823 1207
rect 209866 1204 209872 1216
rect 208811 1176 209872 1204
rect 208811 1173 208823 1176
rect 208765 1167 208823 1173
rect 209866 1164 209872 1176
rect 209924 1164 209930 1216
rect 210053 1207 210111 1213
rect 210053 1173 210065 1207
rect 210099 1204 210111 1207
rect 210326 1204 210332 1216
rect 210099 1176 210332 1204
rect 210099 1173 210111 1176
rect 210053 1167 210111 1173
rect 210326 1164 210332 1176
rect 210384 1164 210390 1216
rect 210697 1207 210755 1213
rect 210697 1173 210709 1207
rect 210743 1204 210755 1207
rect 211264 1204 211292 1244
rect 212534 1232 212540 1244
rect 212592 1232 212598 1284
rect 213288 1272 213316 1439
rect 224770 1436 224776 1488
rect 224828 1476 224834 1488
rect 227806 1476 227812 1488
rect 224828 1448 227812 1476
rect 224828 1436 224834 1448
rect 227806 1436 227812 1448
rect 227864 1436 227870 1488
rect 228376 1476 228404 1516
rect 228453 1513 228465 1547
rect 228499 1544 228511 1547
rect 228818 1544 228824 1556
rect 228499 1516 228824 1544
rect 228499 1513 228511 1516
rect 228453 1507 228511 1513
rect 228818 1504 228824 1516
rect 228876 1504 228882 1556
rect 232501 1547 232559 1553
rect 232501 1513 232513 1547
rect 232547 1544 232559 1547
rect 232590 1544 232596 1556
rect 232547 1516 232596 1544
rect 232547 1513 232559 1516
rect 232501 1507 232559 1513
rect 232590 1504 232596 1516
rect 232648 1504 232654 1556
rect 236181 1547 236239 1553
rect 236181 1513 236193 1547
rect 236227 1544 236239 1547
rect 236546 1544 236552 1556
rect 236227 1516 236552 1544
rect 236227 1513 236239 1516
rect 236181 1507 236239 1513
rect 236546 1504 236552 1516
rect 236604 1504 236610 1556
rect 257062 1544 257068 1556
rect 239416 1516 257068 1544
rect 239416 1476 239444 1516
rect 257062 1504 257068 1516
rect 257120 1504 257126 1556
rect 228376 1448 239444 1476
rect 239490 1436 239496 1488
rect 239548 1476 239554 1488
rect 256970 1476 256976 1488
rect 239548 1448 256976 1476
rect 239548 1436 239554 1448
rect 256970 1436 256976 1448
rect 257028 1436 257034 1488
rect 225414 1368 225420 1420
rect 225472 1408 225478 1420
rect 225509 1411 225567 1417
rect 225509 1408 225521 1411
rect 225472 1380 225521 1408
rect 225472 1368 225478 1380
rect 225509 1377 225521 1380
rect 225555 1377 225567 1411
rect 225509 1371 225567 1377
rect 226521 1411 226579 1417
rect 226521 1377 226533 1411
rect 226567 1408 226579 1411
rect 227070 1408 227076 1420
rect 226567 1380 227076 1408
rect 226567 1377 226579 1380
rect 226521 1371 226579 1377
rect 227070 1368 227076 1380
rect 227128 1368 227134 1420
rect 228085 1411 228143 1417
rect 228085 1377 228097 1411
rect 228131 1408 228143 1411
rect 228174 1408 228180 1420
rect 228131 1380 228180 1408
rect 228131 1377 228143 1380
rect 228085 1371 228143 1377
rect 228174 1368 228180 1380
rect 228232 1368 228238 1420
rect 232133 1411 232191 1417
rect 232133 1377 232145 1411
rect 232179 1408 232191 1411
rect 232498 1408 232504 1420
rect 232179 1380 232504 1408
rect 232179 1377 232191 1380
rect 232133 1371 232191 1377
rect 232498 1368 232504 1380
rect 232556 1368 232562 1420
rect 235442 1368 235448 1420
rect 235500 1408 235506 1420
rect 235813 1411 235871 1417
rect 235813 1408 235825 1411
rect 235500 1380 235825 1408
rect 235500 1368 235506 1380
rect 235813 1377 235825 1380
rect 235859 1377 235871 1411
rect 235813 1371 235871 1377
rect 237190 1368 237196 1420
rect 237248 1408 237254 1420
rect 237248 1380 239904 1408
rect 237248 1368 237254 1380
rect 213454 1300 213460 1352
rect 213512 1300 213518 1352
rect 213730 1300 213736 1352
rect 213788 1340 213794 1352
rect 214101 1343 214159 1349
rect 214101 1340 214113 1343
rect 213788 1312 214113 1340
rect 213788 1300 213794 1312
rect 214101 1309 214113 1312
rect 214147 1309 214159 1343
rect 214101 1303 214159 1309
rect 214466 1300 214472 1352
rect 214524 1340 214530 1352
rect 215389 1343 215447 1349
rect 215389 1340 215401 1343
rect 214524 1312 215401 1340
rect 214524 1300 214530 1312
rect 215389 1309 215401 1312
rect 215435 1309 215447 1343
rect 215389 1303 215447 1309
rect 216033 1343 216091 1349
rect 216033 1309 216045 1343
rect 216079 1309 216091 1343
rect 216033 1303 216091 1309
rect 214558 1272 214564 1284
rect 213288 1244 214564 1272
rect 214558 1232 214564 1244
rect 214616 1232 214622 1284
rect 215110 1232 215116 1284
rect 215168 1272 215174 1284
rect 216048 1272 216076 1303
rect 216674 1300 216680 1352
rect 216732 1300 216738 1352
rect 217778 1300 217784 1352
rect 217836 1300 217842 1352
rect 218146 1300 218152 1352
rect 218204 1340 218210 1352
rect 218701 1343 218759 1349
rect 218701 1340 218713 1343
rect 218204 1312 218713 1340
rect 218204 1300 218210 1312
rect 218701 1309 218713 1312
rect 218747 1309 218759 1343
rect 219805 1343 219863 1349
rect 219805 1340 219817 1343
rect 218701 1303 218759 1309
rect 218808 1312 219817 1340
rect 217594 1272 217600 1284
rect 215168 1244 216076 1272
rect 216508 1244 217600 1272
rect 215168 1232 215174 1244
rect 210743 1176 211292 1204
rect 211341 1207 211399 1213
rect 210743 1173 210755 1176
rect 210697 1167 210755 1173
rect 211341 1173 211353 1207
rect 211387 1204 211399 1207
rect 211798 1204 211804 1216
rect 211387 1176 211804 1204
rect 211387 1173 211399 1176
rect 211341 1167 211399 1173
rect 211798 1164 211804 1176
rect 211856 1164 211862 1216
rect 212629 1207 212687 1213
rect 212629 1173 212641 1207
rect 212675 1204 212687 1207
rect 213822 1204 213828 1216
rect 212675 1176 213828 1204
rect 212675 1173 212687 1176
rect 212629 1167 212687 1173
rect 213822 1164 213828 1176
rect 213880 1164 213886 1216
rect 213917 1207 213975 1213
rect 213917 1173 213929 1207
rect 213963 1204 213975 1207
rect 214374 1204 214380 1216
rect 213963 1176 214380 1204
rect 213963 1173 213975 1176
rect 213917 1167 213975 1173
rect 214374 1164 214380 1176
rect 214432 1164 214438 1216
rect 215202 1164 215208 1216
rect 215260 1164 215266 1216
rect 215570 1164 215576 1216
rect 215628 1204 215634 1216
rect 216508 1213 216536 1244
rect 217594 1232 217600 1244
rect 217652 1232 217658 1284
rect 218054 1232 218060 1284
rect 218112 1232 218118 1284
rect 215849 1207 215907 1213
rect 215849 1204 215861 1207
rect 215628 1176 215861 1204
rect 215628 1164 215634 1176
rect 215849 1173 215861 1176
rect 215895 1173 215907 1207
rect 215849 1167 215907 1173
rect 216493 1207 216551 1213
rect 216493 1173 216505 1207
rect 216539 1173 216551 1207
rect 216493 1167 216551 1173
rect 217410 1164 217416 1216
rect 217468 1204 217474 1216
rect 218808 1204 218836 1312
rect 219805 1309 219817 1312
rect 219851 1309 219863 1343
rect 219805 1303 219863 1309
rect 220541 1343 220599 1349
rect 220541 1309 220553 1343
rect 220587 1309 220599 1343
rect 220541 1303 220599 1309
rect 218974 1232 218980 1284
rect 219032 1232 219038 1284
rect 219434 1232 219440 1284
rect 219492 1272 219498 1284
rect 220556 1272 220584 1303
rect 221182 1300 221188 1352
rect 221240 1300 221246 1352
rect 221829 1343 221887 1349
rect 221829 1309 221841 1343
rect 221875 1309 221887 1343
rect 221829 1303 221887 1309
rect 219492 1244 220584 1272
rect 219492 1232 219498 1244
rect 220722 1232 220728 1284
rect 220780 1272 220786 1284
rect 221844 1272 221872 1303
rect 222194 1300 222200 1352
rect 222252 1340 222258 1352
rect 223117 1343 223175 1349
rect 223117 1340 223129 1343
rect 222252 1312 223129 1340
rect 222252 1300 222258 1312
rect 223117 1309 223129 1312
rect 223163 1309 223175 1343
rect 223117 1303 223175 1309
rect 223758 1300 223764 1352
rect 223816 1300 223822 1352
rect 224865 1343 224923 1349
rect 224865 1340 224877 1343
rect 223868 1312 224877 1340
rect 220780 1244 221872 1272
rect 220780 1232 220786 1244
rect 222286 1232 222292 1284
rect 222344 1272 222350 1284
rect 223868 1272 223896 1312
rect 224865 1309 224877 1312
rect 224911 1309 224923 1343
rect 224865 1303 224923 1309
rect 225693 1343 225751 1349
rect 225693 1309 225705 1343
rect 225739 1340 225751 1343
rect 226610 1340 226616 1352
rect 225739 1312 226616 1340
rect 225739 1309 225751 1312
rect 225693 1303 225751 1309
rect 226610 1300 226616 1312
rect 226668 1340 226674 1352
rect 226705 1343 226763 1349
rect 226705 1340 226717 1343
rect 226668 1312 226717 1340
rect 226668 1300 226674 1312
rect 226705 1309 226717 1312
rect 226751 1309 226763 1343
rect 226705 1303 226763 1309
rect 226886 1300 226892 1352
rect 226944 1300 226950 1352
rect 228269 1343 228327 1349
rect 228269 1309 228281 1343
rect 228315 1340 228327 1343
rect 228358 1340 228364 1352
rect 228315 1312 228364 1340
rect 228315 1309 228327 1312
rect 228269 1303 228327 1309
rect 228358 1300 228364 1312
rect 228416 1300 228422 1352
rect 228913 1343 228971 1349
rect 228913 1309 228925 1343
rect 228959 1340 228971 1343
rect 229278 1340 229284 1352
rect 228959 1312 229284 1340
rect 228959 1309 228971 1312
rect 228913 1303 228971 1309
rect 229278 1300 229284 1312
rect 229336 1300 229342 1352
rect 229646 1300 229652 1352
rect 229704 1300 229710 1352
rect 230658 1300 230664 1352
rect 230716 1300 230722 1352
rect 232314 1300 232320 1352
rect 232372 1300 232378 1352
rect 233234 1300 233240 1352
rect 233292 1300 233298 1352
rect 233970 1300 233976 1352
rect 234028 1300 234034 1352
rect 234706 1300 234712 1352
rect 234764 1300 234770 1352
rect 235994 1300 236000 1352
rect 236052 1300 236058 1352
rect 239876 1340 239904 1380
rect 239950 1368 239956 1420
rect 240008 1368 240014 1420
rect 257706 1408 257712 1420
rect 240060 1380 257712 1408
rect 240060 1340 240088 1380
rect 257706 1368 257712 1380
rect 257764 1368 257770 1420
rect 267734 1368 267740 1420
rect 267792 1408 267798 1420
rect 269301 1411 269359 1417
rect 269301 1408 269313 1411
rect 267792 1380 269313 1408
rect 267792 1368 267798 1380
rect 269301 1377 269313 1380
rect 269347 1377 269359 1411
rect 269301 1371 269359 1377
rect 239876 1312 240088 1340
rect 240962 1300 240968 1352
rect 241020 1300 241026 1352
rect 241054 1300 241060 1352
rect 241112 1340 241118 1352
rect 241241 1343 241299 1349
rect 241241 1340 241253 1343
rect 241112 1312 241253 1340
rect 241112 1300 241118 1312
rect 241241 1309 241253 1312
rect 241287 1309 241299 1343
rect 241241 1303 241299 1309
rect 241974 1300 241980 1352
rect 242032 1340 242038 1352
rect 243541 1343 243599 1349
rect 243541 1340 243553 1343
rect 242032 1312 243553 1340
rect 242032 1300 242038 1312
rect 243541 1309 243553 1312
rect 243587 1309 243599 1343
rect 243541 1303 243599 1309
rect 243814 1300 243820 1352
rect 243872 1300 243878 1352
rect 244918 1300 244924 1352
rect 244976 1340 244982 1352
rect 246117 1343 246175 1349
rect 246117 1340 246129 1343
rect 244976 1312 246129 1340
rect 244976 1300 244982 1312
rect 246117 1309 246129 1312
rect 246163 1309 246175 1343
rect 246117 1303 246175 1309
rect 246206 1300 246212 1352
rect 246264 1340 246270 1352
rect 246393 1343 246451 1349
rect 246393 1340 246405 1343
rect 246264 1312 246405 1340
rect 246264 1300 246270 1312
rect 246393 1309 246405 1312
rect 246439 1309 246451 1343
rect 246393 1303 246451 1309
rect 246482 1300 246488 1352
rect 246540 1340 246546 1352
rect 246540 1312 248460 1340
rect 246540 1300 246546 1312
rect 222344 1244 223896 1272
rect 222344 1232 222350 1244
rect 224034 1232 224040 1284
rect 224092 1232 224098 1284
rect 226242 1232 226248 1284
rect 226300 1272 226306 1284
rect 230198 1272 230204 1284
rect 226300 1244 230204 1272
rect 226300 1232 226306 1244
rect 230198 1232 230204 1244
rect 230256 1232 230262 1284
rect 230382 1232 230388 1284
rect 230440 1272 230446 1284
rect 237374 1272 237380 1284
rect 230440 1244 237380 1272
rect 230440 1232 230446 1244
rect 237374 1232 237380 1244
rect 237432 1232 237438 1284
rect 247957 1275 248015 1281
rect 247957 1241 247969 1275
rect 248003 1272 248015 1275
rect 248322 1272 248328 1284
rect 248003 1244 248328 1272
rect 248003 1241 248015 1244
rect 247957 1235 248015 1241
rect 248322 1232 248328 1244
rect 248380 1232 248386 1284
rect 248432 1272 248460 1312
rect 248506 1300 248512 1352
rect 248564 1340 248570 1352
rect 248693 1343 248751 1349
rect 248693 1340 248705 1343
rect 248564 1312 248705 1340
rect 248564 1300 248570 1312
rect 248693 1309 248705 1312
rect 248739 1309 248751 1343
rect 248693 1303 248751 1309
rect 248966 1300 248972 1352
rect 249024 1300 249030 1352
rect 249076 1312 251404 1340
rect 249076 1272 249104 1312
rect 248432 1244 249104 1272
rect 250162 1232 250168 1284
rect 250220 1232 250226 1284
rect 217468 1176 218836 1204
rect 217468 1164 217474 1176
rect 219618 1164 219624 1216
rect 219676 1164 219682 1216
rect 220354 1164 220360 1216
rect 220412 1164 220418 1216
rect 220906 1164 220912 1216
rect 220964 1204 220970 1216
rect 221001 1207 221059 1213
rect 221001 1204 221013 1207
rect 220964 1176 221013 1204
rect 220964 1164 220970 1176
rect 221001 1173 221013 1176
rect 221047 1173 221059 1207
rect 221001 1167 221059 1173
rect 222933 1207 222991 1213
rect 222933 1173 222945 1207
rect 222979 1204 222991 1207
rect 223114 1204 223120 1216
rect 222979 1176 223120 1204
rect 222979 1173 222991 1176
rect 222933 1167 222991 1173
rect 223114 1164 223120 1176
rect 223172 1164 223178 1216
rect 224681 1207 224739 1213
rect 224681 1173 224693 1207
rect 224727 1204 224739 1207
rect 225046 1204 225052 1216
rect 224727 1176 225052 1204
rect 224727 1173 224739 1176
rect 224681 1167 224739 1173
rect 225046 1164 225052 1176
rect 225104 1164 225110 1216
rect 229094 1164 229100 1216
rect 229152 1164 229158 1216
rect 229830 1164 229836 1216
rect 229888 1164 229894 1216
rect 230842 1164 230848 1216
rect 230900 1164 230906 1216
rect 233418 1164 233424 1216
rect 233476 1164 233482 1216
rect 234154 1164 234160 1216
rect 234212 1164 234218 1216
rect 234890 1164 234896 1216
rect 234948 1164 234954 1216
rect 248046 1164 248052 1216
rect 248104 1164 248110 1216
rect 250254 1164 250260 1216
rect 250312 1164 250318 1216
rect 251376 1204 251404 1312
rect 251542 1300 251548 1352
rect 251600 1300 251606 1352
rect 251818 1300 251824 1352
rect 251876 1300 251882 1352
rect 253474 1300 253480 1352
rect 253532 1340 253538 1352
rect 253845 1343 253903 1349
rect 253845 1340 253857 1343
rect 253532 1312 253857 1340
rect 253532 1300 253538 1312
rect 253845 1309 253857 1312
rect 253891 1309 253903 1343
rect 253845 1303 253903 1309
rect 254118 1300 254124 1352
rect 254176 1300 254182 1352
rect 255222 1300 255228 1352
rect 255280 1340 255286 1352
rect 256421 1343 256479 1349
rect 256421 1340 256433 1343
rect 255280 1312 256433 1340
rect 255280 1300 255286 1312
rect 256421 1309 256433 1312
rect 256467 1309 256479 1343
rect 256421 1303 256479 1309
rect 256510 1300 256516 1352
rect 256568 1340 256574 1352
rect 256697 1343 256755 1349
rect 256697 1340 256709 1343
rect 256568 1312 256709 1340
rect 256568 1300 256574 1312
rect 256697 1309 256709 1312
rect 256743 1309 256755 1343
rect 256697 1303 256755 1309
rect 257798 1300 257804 1352
rect 257856 1340 257862 1352
rect 257893 1343 257951 1349
rect 257893 1340 257905 1343
rect 257856 1312 257905 1340
rect 257856 1300 257862 1312
rect 257893 1309 257905 1312
rect 257939 1309 257951 1343
rect 257893 1303 257951 1309
rect 257982 1300 257988 1352
rect 258040 1340 258046 1352
rect 258077 1343 258135 1349
rect 258077 1340 258089 1343
rect 258040 1312 258089 1340
rect 258040 1300 258046 1312
rect 258077 1309 258089 1312
rect 258123 1309 258135 1343
rect 258077 1303 258135 1309
rect 258997 1343 259055 1349
rect 258997 1309 259009 1343
rect 259043 1309 259055 1343
rect 258997 1303 259055 1309
rect 259273 1343 259331 1349
rect 259273 1309 259285 1343
rect 259319 1309 259331 1343
rect 259273 1303 259331 1309
rect 257430 1232 257436 1284
rect 257488 1272 257494 1284
rect 259012 1272 259040 1303
rect 257488 1244 259040 1272
rect 257488 1232 257494 1244
rect 259288 1204 259316 1303
rect 260282 1300 260288 1352
rect 260340 1300 260346 1352
rect 261570 1300 261576 1352
rect 261628 1300 261634 1352
rect 262306 1300 262312 1352
rect 262364 1300 262370 1352
rect 263042 1300 263048 1352
rect 263100 1300 263106 1352
rect 264146 1300 264152 1352
rect 264204 1300 264210 1352
rect 265158 1300 265164 1352
rect 265216 1300 265222 1352
rect 265894 1300 265900 1352
rect 265952 1300 265958 1352
rect 266722 1300 266728 1352
rect 266780 1300 266786 1352
rect 267461 1343 267519 1349
rect 267461 1309 267473 1343
rect 267507 1340 267519 1343
rect 267826 1340 267832 1352
rect 267507 1312 267832 1340
rect 267507 1309 267519 1312
rect 267461 1303 267519 1309
rect 267826 1300 267832 1312
rect 267884 1300 267890 1352
rect 268194 1300 268200 1352
rect 268252 1300 268258 1352
rect 269206 1300 269212 1352
rect 269264 1340 269270 1352
rect 269485 1343 269543 1349
rect 269485 1340 269497 1343
rect 269264 1312 269497 1340
rect 269264 1300 269270 1312
rect 269485 1309 269497 1312
rect 269531 1309 269543 1343
rect 269485 1303 269543 1309
rect 269669 1343 269727 1349
rect 269669 1309 269681 1343
rect 269715 1340 269727 1343
rect 269850 1340 269856 1352
rect 269715 1312 269856 1340
rect 269715 1309 269727 1312
rect 269669 1303 269727 1309
rect 269850 1300 269856 1312
rect 269908 1300 269914 1352
rect 269942 1300 269948 1352
rect 270000 1340 270006 1352
rect 270129 1343 270187 1349
rect 270129 1340 270141 1343
rect 270000 1312 270141 1340
rect 270000 1300 270006 1312
rect 270129 1309 270141 1312
rect 270175 1309 270187 1343
rect 270129 1303 270187 1309
rect 268930 1232 268936 1284
rect 268988 1272 268994 1284
rect 271782 1272 271788 1284
rect 268988 1244 271788 1272
rect 268988 1232 268994 1244
rect 271782 1232 271788 1244
rect 271840 1232 271846 1284
rect 251376 1176 259316 1204
rect 260466 1164 260472 1216
rect 260524 1164 260530 1216
rect 261754 1164 261760 1216
rect 261812 1164 261818 1216
rect 262490 1164 262496 1216
rect 262548 1164 262554 1216
rect 263226 1164 263232 1216
rect 263284 1164 263290 1216
rect 264330 1164 264336 1216
rect 264388 1164 264394 1216
rect 265342 1164 265348 1216
rect 265400 1164 265406 1216
rect 266078 1164 266084 1216
rect 266136 1164 266142 1216
rect 266906 1164 266912 1216
rect 266964 1164 266970 1216
rect 267642 1164 267648 1216
rect 267700 1164 267706 1216
rect 268378 1164 268384 1216
rect 268436 1164 268442 1216
rect 270310 1164 270316 1216
rect 270368 1164 270374 1216
rect 1104 1114 271651 1136
rect 1104 1062 68546 1114
rect 68598 1062 68610 1114
rect 68662 1062 68674 1114
rect 68726 1062 68738 1114
rect 68790 1062 68802 1114
rect 68854 1062 136143 1114
rect 136195 1062 136207 1114
rect 136259 1062 136271 1114
rect 136323 1062 136335 1114
rect 136387 1062 136399 1114
rect 136451 1062 203740 1114
rect 203792 1062 203804 1114
rect 203856 1062 203868 1114
rect 203920 1062 203932 1114
rect 203984 1062 203996 1114
rect 204048 1062 271337 1114
rect 271389 1062 271401 1114
rect 271453 1062 271465 1114
rect 271517 1062 271529 1114
rect 271581 1062 271593 1114
rect 271645 1062 271651 1114
rect 1104 1040 271651 1062
rect 13538 960 13544 1012
rect 13596 1000 13602 1012
rect 47670 1000 47676 1012
rect 13596 972 47676 1000
rect 13596 960 13602 972
rect 47670 960 47676 972
rect 47728 960 47734 1012
rect 69842 960 69848 1012
rect 69900 1000 69906 1012
rect 96706 1000 96712 1012
rect 69900 972 96712 1000
rect 69900 960 69906 972
rect 96706 960 96712 972
rect 96764 960 96770 1012
rect 105998 960 106004 1012
rect 106056 1000 106062 1012
rect 108850 1000 108856 1012
rect 106056 972 108856 1000
rect 106056 960 106062 972
rect 108850 960 108856 972
rect 108908 960 108914 1012
rect 108942 960 108948 1012
rect 109000 1000 109006 1012
rect 109862 1000 109868 1012
rect 109000 972 109868 1000
rect 109000 960 109006 972
rect 109862 960 109868 972
rect 109920 960 109926 1012
rect 141510 960 141516 1012
rect 141568 1000 141574 1012
rect 174262 1000 174268 1012
rect 141568 972 174268 1000
rect 141568 960 141574 972
rect 174262 960 174268 972
rect 174320 960 174326 1012
rect 207474 960 207480 1012
rect 207532 1000 207538 1012
rect 210234 1000 210240 1012
rect 207532 972 210240 1000
rect 207532 960 207538 972
rect 210234 960 210240 972
rect 210292 960 210298 1012
rect 210326 960 210332 1012
rect 210384 1000 210390 1012
rect 212810 1000 212816 1012
rect 210384 972 212816 1000
rect 210384 960 210390 972
rect 212810 960 212816 972
rect 212868 960 212874 1012
rect 217962 960 217968 1012
rect 218020 1000 218026 1012
rect 219618 1000 219624 1012
rect 218020 972 219624 1000
rect 218020 960 218026 972
rect 219618 960 219624 972
rect 219676 960 219682 1012
rect 246206 1000 246212 1012
rect 220188 972 246212 1000
rect 18690 892 18696 944
rect 18748 932 18754 944
rect 53190 932 53196 944
rect 18748 904 53196 932
rect 18748 892 18754 904
rect 53190 892 53196 904
rect 53248 892 53254 944
rect 82354 892 82360 944
rect 82412 932 82418 944
rect 114830 932 114836 944
rect 82412 904 114836 932
rect 82412 892 82418 904
rect 114830 892 114836 904
rect 114888 892 114894 944
rect 145650 892 145656 944
rect 145708 932 145714 944
rect 147766 932 147772 944
rect 145708 904 147772 932
rect 145708 892 145714 904
rect 147766 892 147772 904
rect 147824 892 147830 944
rect 152090 892 152096 944
rect 152148 932 152154 944
rect 155862 932 155868 944
rect 152148 904 155868 932
rect 152148 892 152154 904
rect 155862 892 155868 904
rect 155920 892 155926 944
rect 182818 932 182824 944
rect 157306 904 182824 932
rect 17218 824 17224 876
rect 17276 864 17282 876
rect 51442 864 51448 876
rect 17276 836 51448 864
rect 17276 824 17282 836
rect 51442 824 51448 836
rect 51500 824 51506 876
rect 82630 824 82636 876
rect 82688 864 82694 876
rect 115106 864 115112 876
rect 82688 836 115112 864
rect 82688 824 82694 836
rect 115106 824 115112 836
rect 115164 824 115170 876
rect 141326 824 141332 876
rect 141384 864 141390 876
rect 152458 864 152464 876
rect 141384 836 152464 864
rect 141384 824 141390 836
rect 152458 824 152464 836
rect 152516 824 152522 876
rect 152550 824 152556 876
rect 152608 864 152614 876
rect 157306 864 157334 904
rect 182818 892 182824 904
rect 182876 892 182882 944
rect 210970 892 210976 944
rect 211028 932 211034 944
rect 216858 932 216864 944
rect 211028 904 216864 932
rect 211028 892 211034 904
rect 216858 892 216864 904
rect 216916 892 216922 944
rect 218054 892 218060 944
rect 218112 932 218118 944
rect 220078 932 220084 944
rect 218112 904 220084 932
rect 218112 892 218118 904
rect 220078 892 220084 904
rect 220136 892 220142 944
rect 152608 836 157334 864
rect 152608 824 152614 836
rect 158898 824 158904 876
rect 158956 864 158962 876
rect 189718 864 189724 876
rect 158956 836 189724 864
rect 158956 824 158962 836
rect 189718 824 189724 836
rect 189776 824 189782 876
rect 211154 824 211160 876
rect 211212 864 211218 876
rect 219802 864 219808 876
rect 211212 836 219808 864
rect 211212 824 211218 836
rect 219802 824 219808 836
rect 219860 824 219866 876
rect 4154 756 4160 808
rect 4212 796 4218 808
rect 38746 796 38752 808
rect 4212 768 38752 796
rect 4212 756 4218 768
rect 38746 756 38752 768
rect 38804 756 38810 808
rect 81434 756 81440 808
rect 81492 796 81498 808
rect 81492 768 104112 796
rect 81492 756 81498 768
rect 12802 688 12808 740
rect 12860 728 12866 740
rect 46290 728 46296 740
rect 12860 700 46296 728
rect 12860 688 12866 700
rect 46290 688 46296 700
rect 46348 688 46354 740
rect 76742 688 76748 740
rect 76800 728 76806 740
rect 100386 728 100392 740
rect 76800 700 100392 728
rect 76800 688 76806 700
rect 100386 688 100392 700
rect 100444 688 100450 740
rect 9674 620 9680 672
rect 9732 660 9738 672
rect 43898 660 43904 672
rect 9732 632 43904 660
rect 9732 620 9738 632
rect 43898 620 43904 632
rect 43956 620 43962 672
rect 73798 620 73804 672
rect 73856 660 73862 672
rect 104084 660 104112 768
rect 104250 756 104256 808
rect 104308 796 104314 808
rect 109954 796 109960 808
rect 104308 768 109960 796
rect 104308 756 104314 768
rect 109954 756 109960 768
rect 110012 756 110018 808
rect 142706 756 142712 808
rect 142764 796 142770 808
rect 204254 796 204260 808
rect 142764 768 204260 796
rect 142764 756 142770 768
rect 204254 756 204260 768
rect 204312 756 204318 808
rect 213638 756 213644 808
rect 213696 796 213702 808
rect 220188 796 220216 972
rect 246206 960 246212 972
rect 246264 960 246270 1012
rect 265526 960 265532 1012
rect 265584 1000 265590 1012
rect 269022 1000 269028 1012
rect 265584 972 269028 1000
rect 265584 960 265590 972
rect 269022 960 269028 972
rect 269080 960 269086 1012
rect 220262 892 220268 944
rect 220320 932 220326 944
rect 223574 932 223580 944
rect 220320 904 223580 932
rect 220320 892 220326 904
rect 223574 892 223580 904
rect 223632 892 223638 944
rect 224862 892 224868 944
rect 224920 932 224926 944
rect 226242 932 226248 944
rect 224920 904 226248 932
rect 224920 892 224926 904
rect 226242 892 226248 904
rect 226300 892 226306 944
rect 229738 892 229744 944
rect 229796 932 229802 944
rect 254118 932 254124 944
rect 229796 904 254124 932
rect 229796 892 229802 904
rect 254118 892 254124 904
rect 254176 892 254182 944
rect 222010 824 222016 876
rect 222068 864 222074 876
rect 250254 864 250260 876
rect 222068 836 250260 864
rect 222068 824 222074 836
rect 250254 824 250260 836
rect 250312 824 250318 876
rect 213696 768 220216 796
rect 213696 756 213702 768
rect 221550 756 221556 808
rect 221608 796 221614 808
rect 254026 796 254032 808
rect 221608 768 254032 796
rect 221608 756 221614 768
rect 254026 756 254032 768
rect 254084 756 254090 808
rect 107194 688 107200 740
rect 107252 728 107258 740
rect 108850 728 108856 740
rect 107252 700 108856 728
rect 107252 688 107258 700
rect 108850 688 108856 700
rect 108908 688 108914 740
rect 112714 728 112720 740
rect 109006 700 112720 728
rect 73856 632 89714 660
rect 104084 632 105584 660
rect 73856 620 73862 632
rect 8386 552 8392 604
rect 8444 592 8450 604
rect 40218 592 40224 604
rect 8444 564 40224 592
rect 8444 552 8450 564
rect 40218 552 40224 564
rect 40276 552 40282 604
rect 74994 552 75000 604
rect 75052 592 75058 604
rect 89686 592 89714 632
rect 101858 592 101864 604
rect 75052 564 84194 592
rect 89686 564 101864 592
rect 75052 552 75058 564
rect 17954 484 17960 536
rect 18012 524 18018 536
rect 51810 524 51816 536
rect 18012 496 51816 524
rect 18012 484 18018 496
rect 51810 484 51816 496
rect 51868 484 51874 536
rect 84166 524 84194 564
rect 101858 552 101864 564
rect 101916 552 101922 604
rect 105078 524 105084 536
rect 84166 496 105084 524
rect 105078 484 105084 496
rect 105136 484 105142 536
rect 105556 524 105584 632
rect 107562 620 107568 672
rect 107620 660 107626 672
rect 109006 660 109034 700
rect 112714 688 112720 700
rect 112772 688 112778 740
rect 146754 688 146760 740
rect 146812 728 146818 740
rect 179414 728 179420 740
rect 146812 700 179420 728
rect 146812 688 146818 700
rect 179414 688 179420 700
rect 179472 688 179478 740
rect 207198 688 207204 740
rect 207256 728 207262 740
rect 217318 728 217324 740
rect 207256 700 217324 728
rect 207256 688 207262 700
rect 217318 688 217324 700
rect 217376 688 217382 740
rect 218882 688 218888 740
rect 218940 728 218946 740
rect 221182 728 221188 740
rect 218940 700 221188 728
rect 218940 688 218946 700
rect 221182 688 221188 700
rect 221240 688 221246 740
rect 224770 688 224776 740
rect 224828 728 224834 740
rect 258350 728 258356 740
rect 224828 700 258356 728
rect 224828 688 224834 700
rect 258350 688 258356 700
rect 258408 688 258414 740
rect 107620 632 109034 660
rect 107620 620 107626 632
rect 143902 620 143908 672
rect 143960 660 143966 672
rect 176838 660 176844 672
rect 143960 632 176844 660
rect 143960 620 143966 632
rect 176838 620 176844 632
rect 176896 620 176902 672
rect 208854 620 208860 672
rect 208912 660 208918 672
rect 241054 660 241060 672
rect 208912 632 241060 660
rect 208912 620 208918 632
rect 241054 620 241060 632
rect 241112 620 241118 672
rect 111978 592 111984 604
rect 108960 564 111984 592
rect 108960 524 108988 564
rect 111978 552 111984 564
rect 112036 552 112042 604
rect 138658 552 138664 604
rect 138716 592 138722 604
rect 172514 592 172520 604
rect 138716 564 172520 592
rect 138716 552 138722 564
rect 172514 552 172520 564
rect 172572 552 172578 604
rect 217318 552 217324 604
rect 217376 592 217382 604
rect 223022 592 223028 604
rect 217376 564 223028 592
rect 217376 552 217382 564
rect 223022 552 223028 564
rect 223080 552 223086 604
rect 223114 552 223120 604
rect 223172 592 223178 604
rect 248966 592 248972 604
rect 223172 564 248972 592
rect 223172 552 223178 564
rect 248966 552 248972 564
rect 249024 552 249030 604
rect 105556 496 108988 524
rect 152458 484 152464 536
rect 152516 524 152522 536
rect 158346 524 158352 536
rect 152516 496 158352 524
rect 152516 484 152522 496
rect 158346 484 158352 496
rect 158404 484 158410 536
rect 187142 524 187148 536
rect 161446 496 187148 524
rect 5442 416 5448 468
rect 5500 456 5506 468
rect 40126 456 40132 468
rect 5500 428 40132 456
rect 5500 416 5506 428
rect 40126 416 40132 428
rect 40184 416 40190 468
rect 72418 416 72424 468
rect 72476 456 72482 468
rect 99742 456 99748 468
rect 72476 428 99748 456
rect 72476 416 72482 428
rect 99742 416 99748 428
rect 99800 416 99806 468
rect 100386 416 100392 468
rect 100444 456 100450 468
rect 106366 456 106372 468
rect 100444 428 106372 456
rect 100444 416 100450 428
rect 106366 416 106372 428
rect 106424 416 106430 468
rect 148778 416 148784 468
rect 148836 456 148842 468
rect 160462 456 160468 468
rect 148836 428 160468 456
rect 148836 416 148842 428
rect 160462 416 160468 428
rect 160520 416 160526 468
rect 2866 348 2872 400
rect 2924 388 2930 400
rect 37734 388 37740 400
rect 2924 360 37740 388
rect 2924 348 2930 360
rect 37734 348 37740 360
rect 37792 348 37798 400
rect 151538 348 151544 400
rect 151596 388 151602 400
rect 152550 388 152556 400
rect 151596 360 152556 388
rect 151596 348 151602 360
rect 152550 348 152556 360
rect 152608 348 152614 400
rect 154298 348 154304 400
rect 154356 388 154362 400
rect 161446 388 161474 496
rect 187142 484 187148 496
rect 187200 484 187206 536
rect 211062 484 211068 536
rect 211120 524 211126 536
rect 243814 524 243820 536
rect 211120 496 243820 524
rect 211120 484 211126 496
rect 243814 484 243820 496
rect 243872 484 243878 536
rect 211338 416 211344 468
rect 211396 456 211402 468
rect 211396 428 215294 456
rect 211396 416 211402 428
rect 154356 360 161474 388
rect 215266 388 215294 428
rect 216582 416 216588 468
rect 216640 456 216646 468
rect 227990 456 227996 468
rect 216640 428 227996 456
rect 216640 416 216646 428
rect 227990 416 227996 428
rect 228048 416 228054 468
rect 256510 456 256516 468
rect 234586 428 256516 456
rect 217870 388 217876 400
rect 215266 360 217876 388
rect 154356 348 154362 360
rect 217870 348 217876 360
rect 217928 348 217934 400
rect 219618 348 219624 400
rect 219676 388 219682 400
rect 220722 388 220728 400
rect 219676 360 220728 388
rect 219676 348 219682 360
rect 220722 348 220728 360
rect 220780 348 220786 400
rect 224126 348 224132 400
rect 224184 388 224190 400
rect 234586 388 234614 428
rect 256510 416 256516 428
rect 256568 416 256574 468
rect 224184 360 234614 388
rect 224184 348 224190 360
rect 235718 348 235724 400
rect 235776 388 235782 400
rect 268930 388 268936 400
rect 235776 360 268936 388
rect 235776 348 235782 360
rect 268930 348 268936 360
rect 268988 348 268994 400
rect 9398 280 9404 332
rect 9456 320 9462 332
rect 41046 320 41052 332
rect 9456 292 41052 320
rect 9456 280 9462 292
rect 41046 280 41052 292
rect 41104 280 41110 332
rect 216214 280 216220 332
rect 216272 320 216278 332
rect 223114 320 223120 332
rect 216272 292 223120 320
rect 216272 280 216278 292
rect 223114 280 223120 292
rect 223172 280 223178 332
rect 227898 280 227904 332
rect 227956 320 227962 332
rect 251818 320 251824 332
rect 227956 292 251824 320
rect 227956 280 227962 292
rect 251818 280 251824 292
rect 251876 280 251882 332
rect 222838 212 222844 264
rect 222896 252 222902 264
rect 229738 252 229744 264
rect 222896 224 229744 252
rect 222896 212 222902 224
rect 229738 212 229744 224
rect 229796 212 229802 264
<< via1 >>
rect 97632 10820 97684 10872
rect 98460 10820 98512 10872
rect 28448 10684 28500 10736
rect 33784 10684 33836 10736
rect 29920 10616 29972 10668
rect 23940 10548 23992 10600
rect 63224 10616 63276 10668
rect 90824 10752 90876 10804
rect 95056 10752 95108 10804
rect 96988 10752 97040 10804
rect 152372 10820 152424 10872
rect 163964 10820 164016 10872
rect 214288 10820 214340 10872
rect 227444 10820 227496 10872
rect 229100 10820 229152 10872
rect 233608 10820 233660 10872
rect 233700 10820 233752 10872
rect 246764 10820 246816 10872
rect 258540 10820 258592 10872
rect 267832 10820 267884 10872
rect 132868 10752 132920 10804
rect 133696 10752 133748 10804
rect 152464 10752 152516 10804
rect 164148 10752 164200 10804
rect 164332 10752 164384 10804
rect 239404 10752 239456 10804
rect 255688 10752 255740 10804
rect 267740 10752 267792 10804
rect 65984 10684 66036 10736
rect 99380 10684 99432 10736
rect 104348 10684 104400 10736
rect 130568 10684 130620 10736
rect 164608 10684 164660 10736
rect 164792 10684 164844 10736
rect 264796 10684 264848 10736
rect 75000 10616 75052 10668
rect 104808 10616 104860 10668
rect 23756 10480 23808 10532
rect 30012 10480 30064 10532
rect 25780 10412 25832 10464
rect 20720 10344 20772 10396
rect 25964 10344 26016 10396
rect 22836 10276 22888 10328
rect 24952 10276 25004 10328
rect 26056 10208 26108 10260
rect 29092 10208 29144 10260
rect 7656 10072 7708 10124
rect 26700 10072 26752 10124
rect 5908 10004 5960 10056
rect 23664 10004 23716 10056
rect 17316 9936 17368 9988
rect 27620 10140 27672 10192
rect 60372 10548 60424 10600
rect 94964 10548 95016 10600
rect 96988 10548 97040 10600
rect 129464 10548 129516 10600
rect 60096 10480 60148 10532
rect 90824 10480 90876 10532
rect 91008 10480 91060 10532
rect 57152 10412 57204 10464
rect 92388 10412 92440 10464
rect 94044 10480 94096 10532
rect 96712 10480 96764 10532
rect 131120 10480 131172 10532
rect 165344 10616 165396 10668
rect 225328 10616 225380 10668
rect 226432 10616 226484 10668
rect 133696 10548 133748 10600
rect 167092 10548 167144 10600
rect 196716 10548 196768 10600
rect 227536 10548 227588 10600
rect 133788 10480 133840 10532
rect 167736 10480 167788 10532
rect 192484 10480 192536 10532
rect 224592 10480 224644 10532
rect 225420 10480 225472 10532
rect 233424 10548 233476 10600
rect 227720 10480 227772 10532
rect 230848 10480 230900 10532
rect 233792 10616 233844 10668
rect 233608 10548 233660 10600
rect 258356 10548 258408 10600
rect 258724 10616 258776 10668
rect 266820 10616 266872 10668
rect 260196 10548 260248 10600
rect 260288 10548 260340 10600
rect 263140 10548 263192 10600
rect 258448 10480 258500 10532
rect 258816 10480 258868 10532
rect 268200 10480 268252 10532
rect 125048 10412 125100 10464
rect 162308 10412 162360 10464
rect 263600 10412 263652 10464
rect 33784 10344 33836 10396
rect 62396 10344 62448 10396
rect 94044 10344 94096 10396
rect 57152 10276 57204 10328
rect 61476 10276 61528 10328
rect 96436 10344 96488 10396
rect 59636 10208 59688 10260
rect 66076 10208 66128 10260
rect 98368 10344 98420 10396
rect 99288 10344 99340 10396
rect 103520 10344 103572 10396
rect 104348 10344 104400 10396
rect 133972 10344 134024 10396
rect 151728 10344 151780 10396
rect 181996 10344 182048 10396
rect 202788 10344 202840 10396
rect 235724 10344 235776 10396
rect 255872 10344 255924 10396
rect 268016 10344 268068 10396
rect 30380 10140 30432 10192
rect 64052 10140 64104 10192
rect 77484 10140 77536 10192
rect 103336 10276 103388 10328
rect 97632 10208 97684 10260
rect 131856 10276 131908 10328
rect 103520 10208 103572 10260
rect 132960 10208 133012 10260
rect 133788 10208 133840 10260
rect 149060 10276 149112 10328
rect 172520 10276 172572 10328
rect 193220 10276 193272 10328
rect 225328 10276 225380 10328
rect 225512 10276 225564 10328
rect 227720 10276 227772 10328
rect 228088 10276 228140 10328
rect 166264 10208 166316 10260
rect 170312 10208 170364 10260
rect 208400 10208 208452 10260
rect 97540 10140 97592 10192
rect 103704 10140 103756 10192
rect 122748 10140 122800 10192
rect 156512 10140 156564 10192
rect 162216 10140 162268 10192
rect 218336 10208 218388 10260
rect 230664 10208 230716 10260
rect 230848 10276 230900 10328
rect 258172 10276 258224 10328
rect 258632 10276 258684 10328
rect 266636 10276 266688 10328
rect 258356 10208 258408 10260
rect 258908 10208 258960 10260
rect 267004 10208 267056 10260
rect 262864 10140 262916 10192
rect 8484 9868 8536 9920
rect 33048 10004 33100 10056
rect 56416 10072 56468 10124
rect 91008 10072 91060 10124
rect 93216 10072 93268 10124
rect 126704 10072 126756 10124
rect 55404 10004 55456 10056
rect 92388 10004 92440 10056
rect 102416 10004 102468 10056
rect 27068 9936 27120 9988
rect 29000 9936 29052 9988
rect 31208 9936 31260 9988
rect 64972 9936 65024 9988
rect 66076 9936 66128 9988
rect 76748 9936 76800 9988
rect 101680 9936 101732 9988
rect 122748 10004 122800 10056
rect 158628 10072 158680 10124
rect 182456 10072 182508 10124
rect 198648 10072 198700 10124
rect 218152 10072 218204 10124
rect 218244 10072 218296 10124
rect 225512 10072 225564 10124
rect 225604 10072 225656 10124
rect 233700 10072 233752 10124
rect 258632 10072 258684 10124
rect 262404 10072 262456 10124
rect 270408 10140 270460 10192
rect 263324 10072 263376 10124
rect 268936 10072 268988 10124
rect 160928 10004 160980 10056
rect 163688 10004 163740 10056
rect 243084 10004 243136 10056
rect 257988 10004 258040 10056
rect 265900 10004 265952 10056
rect 266268 10004 266320 10056
rect 269028 10004 269080 10056
rect 26976 9868 27028 9920
rect 31852 9868 31904 9920
rect 58900 9868 58952 9920
rect 92848 9868 92900 9920
rect 92940 9868 92992 9920
rect 124128 9936 124180 9988
rect 158720 9936 158772 9988
rect 162584 9936 162636 9988
rect 165252 9936 165304 9988
rect 258724 9936 258776 9988
rect 261024 9936 261076 9988
rect 267924 9936 267976 9988
rect 102416 9868 102468 9920
rect 113824 9868 113876 9920
rect 121276 9868 121328 9920
rect 127624 9868 127676 9920
rect 161388 9868 161440 9920
rect 163596 9868 163648 9920
rect 187056 9868 187108 9920
rect 199660 9868 199712 9920
rect 229192 9868 229244 9920
rect 229468 9868 229520 9920
rect 263968 9868 264020 9920
rect 264980 9868 265032 9920
rect 268476 9868 268528 9920
rect 68546 9766 68598 9818
rect 68610 9766 68662 9818
rect 68674 9766 68726 9818
rect 68738 9766 68790 9818
rect 68802 9766 68854 9818
rect 136143 9766 136195 9818
rect 136207 9766 136259 9818
rect 136271 9766 136323 9818
rect 136335 9766 136387 9818
rect 136399 9766 136451 9818
rect 203740 9766 203792 9818
rect 203804 9766 203856 9818
rect 203868 9766 203920 9818
rect 203932 9766 203984 9818
rect 203996 9766 204048 9818
rect 271337 9766 271389 9818
rect 271401 9766 271453 9818
rect 271465 9766 271517 9818
rect 271529 9766 271581 9818
rect 271593 9766 271645 9818
rect 5908 9707 5960 9716
rect 5908 9673 5917 9707
rect 5917 9673 5951 9707
rect 5951 9673 5960 9707
rect 5908 9664 5960 9673
rect 7656 9707 7708 9716
rect 7656 9673 7665 9707
rect 7665 9673 7699 9707
rect 7699 9673 7708 9707
rect 7656 9664 7708 9673
rect 8484 9707 8536 9716
rect 8484 9673 8493 9707
rect 8493 9673 8527 9707
rect 8527 9673 8536 9707
rect 8484 9664 8536 9673
rect 51080 9664 51132 9716
rect 54668 9707 54720 9716
rect 54668 9673 54677 9707
rect 54677 9673 54711 9707
rect 54711 9673 54720 9707
rect 54668 9664 54720 9673
rect 57796 9664 57848 9716
rect 59268 9707 59320 9716
rect 59268 9673 59277 9707
rect 59277 9673 59311 9707
rect 59311 9673 59320 9707
rect 59268 9664 59320 9673
rect 60004 9707 60056 9716
rect 60004 9673 60013 9707
rect 60013 9673 60047 9707
rect 60047 9673 60056 9707
rect 60004 9664 60056 9673
rect 60832 9707 60884 9716
rect 60832 9673 60841 9707
rect 60841 9673 60875 9707
rect 60875 9673 60884 9707
rect 60832 9664 60884 9673
rect 63408 9707 63460 9716
rect 63408 9673 63417 9707
rect 63417 9673 63451 9707
rect 63451 9673 63460 9707
rect 63408 9664 63460 9673
rect 66168 9707 66220 9716
rect 66168 9673 66177 9707
rect 66177 9673 66211 9707
rect 66211 9673 66220 9707
rect 66168 9664 66220 9673
rect 66904 9707 66956 9716
rect 66904 9673 66913 9707
rect 66913 9673 66947 9707
rect 66947 9673 66956 9707
rect 66904 9664 66956 9673
rect 90272 9664 90324 9716
rect 90364 9707 90416 9716
rect 90364 9673 90373 9707
rect 90373 9673 90407 9707
rect 90407 9673 90416 9707
rect 90364 9664 90416 9673
rect 93492 9707 93544 9716
rect 93492 9673 93501 9707
rect 93501 9673 93535 9707
rect 93535 9673 93544 9707
rect 93492 9664 93544 9673
rect 95976 9707 96028 9716
rect 95976 9673 95985 9707
rect 95985 9673 96019 9707
rect 96019 9673 96028 9707
rect 95976 9664 96028 9673
rect 96344 9664 96396 9716
rect 98000 9664 98052 9716
rect 98276 9664 98328 9716
rect 1676 9639 1728 9648
rect 1676 9605 1685 9639
rect 1685 9605 1719 9639
rect 1719 9605 1728 9639
rect 1676 9596 1728 9605
rect 2412 9639 2464 9648
rect 2412 9605 2421 9639
rect 2421 9605 2455 9639
rect 2455 9605 2464 9639
rect 2412 9596 2464 9605
rect 3240 9639 3292 9648
rect 3240 9605 3249 9639
rect 3249 9605 3283 9639
rect 3283 9605 3292 9639
rect 3240 9596 3292 9605
rect 4344 9639 4396 9648
rect 4344 9605 4353 9639
rect 4353 9605 4387 9639
rect 4387 9605 4396 9639
rect 4344 9596 4396 9605
rect 5080 9639 5132 9648
rect 5080 9605 5089 9639
rect 5089 9605 5123 9639
rect 5123 9605 5132 9639
rect 5080 9596 5132 9605
rect 5816 9639 5868 9648
rect 5816 9605 5825 9639
rect 5825 9605 5859 9639
rect 5859 9605 5868 9639
rect 5816 9596 5868 9605
rect 6828 9639 6880 9648
rect 6828 9605 6837 9639
rect 6837 9605 6871 9639
rect 6871 9605 6880 9639
rect 6828 9596 6880 9605
rect 7564 9639 7616 9648
rect 7564 9605 7573 9639
rect 7573 9605 7607 9639
rect 7607 9605 7616 9639
rect 7564 9596 7616 9605
rect 8392 9639 8444 9648
rect 8392 9605 8401 9639
rect 8401 9605 8435 9639
rect 8435 9605 8444 9639
rect 8392 9596 8444 9605
rect 11980 9639 12032 9648
rect 11980 9605 11989 9639
rect 11989 9605 12023 9639
rect 12023 9605 12032 9639
rect 11980 9596 12032 9605
rect 12716 9639 12768 9648
rect 12716 9605 12725 9639
rect 12725 9605 12759 9639
rect 12759 9605 12768 9639
rect 12716 9596 12768 9605
rect 13728 9596 13780 9648
rect 14648 9639 14700 9648
rect 14648 9605 14657 9639
rect 14657 9605 14691 9639
rect 14691 9605 14700 9639
rect 14648 9596 14700 9605
rect 15384 9639 15436 9648
rect 15384 9605 15393 9639
rect 15393 9605 15427 9639
rect 15427 9605 15436 9639
rect 15384 9596 15436 9605
rect 16120 9639 16172 9648
rect 16120 9605 16129 9639
rect 16129 9605 16163 9639
rect 16163 9605 16172 9639
rect 16120 9596 16172 9605
rect 17132 9639 17184 9648
rect 17132 9605 17141 9639
rect 17141 9605 17175 9639
rect 17175 9605 17184 9639
rect 17132 9596 17184 9605
rect 17316 9639 17368 9648
rect 17316 9605 17325 9639
rect 17325 9605 17359 9639
rect 17359 9605 17368 9639
rect 17316 9596 17368 9605
rect 17868 9639 17920 9648
rect 17868 9605 17877 9639
rect 17877 9605 17911 9639
rect 17911 9605 17920 9639
rect 17868 9596 17920 9605
rect 18604 9639 18656 9648
rect 18604 9605 18613 9639
rect 18613 9605 18647 9639
rect 18647 9605 18656 9639
rect 18604 9596 18656 9605
rect 9680 9571 9732 9580
rect 9680 9537 9689 9571
rect 9689 9537 9723 9571
rect 9723 9537 9732 9571
rect 9680 9528 9732 9537
rect 22376 9596 22428 9648
rect 28908 9596 28960 9648
rect 29000 9596 29052 9648
rect 46204 9596 46256 9648
rect 9956 9503 10008 9512
rect 9956 9469 9965 9503
rect 9965 9469 9999 9503
rect 9999 9469 10008 9503
rect 9956 9460 10008 9469
rect 14740 9460 14792 9512
rect 23572 9528 23624 9580
rect 23756 9571 23808 9580
rect 23756 9537 23765 9571
rect 23765 9537 23799 9571
rect 23799 9537 23808 9571
rect 23756 9528 23808 9537
rect 23848 9571 23900 9580
rect 23848 9537 23857 9571
rect 23857 9537 23891 9571
rect 23891 9537 23900 9571
rect 23848 9528 23900 9537
rect 25136 9571 25188 9580
rect 25136 9537 25145 9571
rect 25145 9537 25179 9571
rect 25179 9537 25188 9571
rect 25136 9528 25188 9537
rect 27528 9528 27580 9580
rect 3424 9435 3476 9444
rect 3424 9401 3433 9435
rect 3433 9401 3467 9435
rect 3467 9401 3476 9435
rect 3424 9392 3476 9401
rect 2412 9324 2464 9376
rect 2504 9367 2556 9376
rect 2504 9333 2513 9367
rect 2513 9333 2547 9367
rect 2547 9333 2556 9367
rect 2504 9324 2556 9333
rect 6920 9367 6972 9376
rect 6920 9333 6929 9367
rect 6929 9333 6963 9367
rect 6963 9333 6972 9367
rect 6920 9324 6972 9333
rect 12808 9367 12860 9376
rect 12808 9333 12817 9367
rect 12817 9333 12851 9367
rect 12851 9333 12860 9367
rect 12808 9324 12860 9333
rect 13728 9435 13780 9444
rect 13728 9401 13737 9435
rect 13737 9401 13771 9435
rect 13771 9401 13780 9435
rect 13728 9392 13780 9401
rect 15568 9435 15620 9444
rect 15568 9401 15577 9435
rect 15577 9401 15611 9435
rect 15611 9401 15620 9435
rect 15568 9392 15620 9401
rect 20352 9392 20404 9444
rect 15292 9324 15344 9376
rect 24400 9392 24452 9444
rect 23388 9324 23440 9376
rect 23756 9324 23808 9376
rect 23940 9324 23992 9376
rect 24492 9324 24544 9376
rect 26056 9460 26108 9512
rect 27712 9460 27764 9512
rect 28724 9528 28776 9580
rect 29736 9571 29788 9580
rect 29736 9537 29745 9571
rect 29745 9537 29779 9571
rect 29779 9537 29788 9571
rect 29736 9528 29788 9537
rect 32680 9528 32732 9580
rect 35624 9571 35676 9580
rect 35624 9537 35633 9571
rect 35633 9537 35667 9571
rect 35667 9537 35676 9571
rect 35624 9528 35676 9537
rect 36268 9571 36320 9580
rect 36268 9537 36277 9571
rect 36277 9537 36311 9571
rect 36311 9537 36320 9571
rect 36268 9528 36320 9537
rect 36912 9571 36964 9580
rect 36912 9537 36921 9571
rect 36921 9537 36955 9571
rect 36955 9537 36964 9571
rect 36912 9528 36964 9537
rect 38108 9571 38160 9580
rect 38108 9537 38117 9571
rect 38117 9537 38151 9571
rect 38151 9537 38160 9571
rect 38108 9528 38160 9537
rect 38844 9571 38896 9580
rect 38844 9537 38853 9571
rect 38853 9537 38887 9571
rect 38887 9537 38896 9571
rect 38844 9528 38896 9537
rect 39488 9571 39540 9580
rect 39488 9537 39497 9571
rect 39497 9537 39531 9571
rect 39531 9537 39540 9571
rect 39488 9528 39540 9537
rect 40776 9571 40828 9580
rect 40776 9537 40785 9571
rect 40785 9537 40819 9571
rect 40819 9537 40828 9571
rect 40776 9528 40828 9537
rect 41420 9571 41472 9580
rect 41420 9537 41429 9571
rect 41429 9537 41463 9571
rect 41463 9537 41472 9571
rect 41420 9528 41472 9537
rect 42064 9571 42116 9580
rect 42064 9537 42073 9571
rect 42073 9537 42107 9571
rect 42107 9537 42116 9571
rect 42064 9528 42116 9537
rect 43260 9571 43312 9580
rect 43260 9537 43269 9571
rect 43269 9537 43303 9571
rect 43303 9537 43312 9571
rect 43260 9528 43312 9537
rect 43996 9571 44048 9580
rect 43996 9537 44005 9571
rect 44005 9537 44039 9571
rect 44039 9537 44048 9571
rect 43996 9528 44048 9537
rect 44640 9571 44692 9580
rect 44640 9537 44649 9571
rect 44649 9537 44683 9571
rect 44683 9537 44692 9571
rect 44640 9528 44692 9537
rect 45928 9571 45980 9580
rect 45928 9537 45937 9571
rect 45937 9537 45971 9571
rect 45971 9537 45980 9571
rect 45928 9528 45980 9537
rect 60096 9596 60148 9648
rect 29000 9460 29052 9512
rect 29092 9460 29144 9512
rect 46572 9571 46624 9580
rect 46572 9537 46581 9571
rect 46581 9537 46615 9571
rect 46615 9537 46624 9571
rect 46572 9528 46624 9537
rect 47216 9571 47268 9580
rect 47216 9537 47225 9571
rect 47225 9537 47259 9571
rect 47259 9537 47268 9571
rect 47216 9528 47268 9537
rect 48228 9528 48280 9580
rect 49148 9571 49200 9580
rect 49148 9537 49157 9571
rect 49157 9537 49191 9571
rect 49191 9537 49200 9571
rect 49148 9528 49200 9537
rect 49792 9571 49844 9580
rect 49792 9537 49801 9571
rect 49801 9537 49835 9571
rect 49835 9537 49844 9571
rect 49792 9528 49844 9537
rect 50620 9571 50672 9580
rect 50620 9537 50629 9571
rect 50629 9537 50663 9571
rect 50663 9537 50672 9571
rect 50620 9528 50672 9537
rect 51356 9571 51408 9580
rect 51356 9537 51365 9571
rect 51365 9537 51399 9571
rect 51399 9537 51408 9571
rect 51356 9528 51408 9537
rect 52092 9571 52144 9580
rect 52092 9537 52101 9571
rect 52101 9537 52135 9571
rect 52135 9537 52144 9571
rect 52092 9528 52144 9537
rect 53012 9571 53064 9580
rect 53012 9537 53021 9571
rect 53021 9537 53055 9571
rect 53055 9537 53064 9571
rect 53012 9528 53064 9537
rect 54024 9528 54076 9580
rect 54116 9528 54168 9580
rect 57520 9528 57572 9580
rect 59176 9528 59228 9580
rect 60004 9528 60056 9580
rect 60740 9528 60792 9580
rect 62764 9528 62816 9580
rect 66352 9528 66404 9580
rect 66996 9528 67048 9580
rect 69112 9571 69164 9580
rect 69112 9537 69121 9571
rect 69121 9537 69155 9571
rect 69155 9537 69164 9571
rect 69112 9528 69164 9537
rect 70308 9528 70360 9580
rect 72148 9571 72200 9580
rect 72148 9537 72157 9571
rect 72157 9537 72191 9571
rect 72191 9537 72200 9571
rect 72148 9528 72200 9537
rect 94136 9596 94188 9648
rect 100668 9707 100720 9716
rect 100668 9673 100677 9707
rect 100677 9673 100711 9707
rect 100711 9673 100720 9707
rect 100668 9664 100720 9673
rect 103704 9707 103756 9716
rect 103704 9673 103713 9707
rect 103713 9673 103747 9707
rect 103747 9673 103756 9707
rect 103704 9664 103756 9673
rect 104716 9707 104768 9716
rect 104716 9673 104725 9707
rect 104725 9673 104759 9707
rect 104759 9673 104768 9707
rect 104716 9664 104768 9673
rect 105452 9707 105504 9716
rect 105452 9673 105461 9707
rect 105461 9673 105495 9707
rect 105495 9673 105504 9707
rect 105452 9664 105504 9673
rect 105912 9664 105964 9716
rect 108948 9664 109000 9716
rect 113824 9664 113876 9716
rect 74724 9571 74776 9580
rect 74724 9537 74733 9571
rect 74733 9537 74767 9571
rect 74767 9537 74776 9571
rect 74724 9528 74776 9537
rect 77300 9571 77352 9580
rect 77300 9537 77309 9571
rect 77309 9537 77343 9571
rect 77343 9537 77352 9571
rect 77300 9528 77352 9537
rect 79968 9528 80020 9580
rect 82636 9528 82688 9580
rect 84568 9571 84620 9580
rect 84568 9537 84577 9571
rect 84577 9537 84611 9571
rect 84611 9537 84620 9571
rect 84568 9528 84620 9537
rect 86776 9571 86828 9580
rect 86776 9537 86785 9571
rect 86785 9537 86819 9571
rect 86819 9537 86828 9571
rect 86776 9528 86828 9537
rect 89168 9528 89220 9580
rect 90180 9571 90232 9580
rect 90180 9537 90189 9571
rect 90189 9537 90223 9571
rect 90223 9537 90232 9571
rect 90180 9528 90232 9537
rect 93676 9528 93728 9580
rect 46296 9460 46348 9512
rect 25872 9392 25924 9444
rect 26884 9324 26936 9376
rect 28172 9367 28224 9376
rect 28172 9333 28181 9367
rect 28181 9333 28215 9367
rect 28215 9333 28224 9367
rect 28172 9324 28224 9333
rect 28816 9435 28868 9444
rect 28816 9401 28825 9435
rect 28825 9401 28859 9435
rect 28859 9401 28868 9435
rect 28816 9392 28868 9401
rect 32588 9435 32640 9444
rect 32588 9401 32597 9435
rect 32597 9401 32631 9435
rect 32631 9401 32640 9435
rect 32588 9392 32640 9401
rect 30012 9324 30064 9376
rect 46204 9392 46256 9444
rect 47768 9392 47820 9444
rect 55864 9460 55916 9512
rect 61476 9460 61528 9512
rect 75828 9460 75880 9512
rect 77576 9503 77628 9512
rect 77576 9469 77585 9503
rect 77585 9469 77619 9503
rect 77619 9469 77628 9503
rect 77576 9460 77628 9469
rect 81348 9460 81400 9512
rect 82728 9503 82780 9512
rect 82728 9469 82737 9503
rect 82737 9469 82771 9503
rect 82771 9469 82780 9503
rect 82728 9460 82780 9469
rect 84844 9503 84896 9512
rect 84844 9469 84853 9503
rect 84853 9469 84887 9503
rect 84887 9469 84896 9503
rect 84844 9460 84896 9469
rect 87052 9503 87104 9512
rect 87052 9469 87061 9503
rect 87061 9469 87095 9503
rect 87095 9469 87104 9503
rect 87052 9460 87104 9469
rect 87788 9460 87840 9512
rect 53748 9392 53800 9444
rect 35808 9324 35860 9376
rect 36636 9324 36688 9376
rect 37096 9324 37148 9376
rect 37924 9367 37976 9376
rect 37924 9333 37933 9367
rect 37933 9333 37967 9367
rect 37967 9333 37976 9367
rect 37924 9324 37976 9333
rect 38108 9324 38160 9376
rect 39304 9367 39356 9376
rect 39304 9333 39313 9367
rect 39313 9333 39347 9367
rect 39347 9333 39356 9367
rect 39304 9324 39356 9333
rect 40868 9324 40920 9376
rect 41696 9324 41748 9376
rect 41880 9367 41932 9376
rect 41880 9333 41889 9367
rect 41889 9333 41923 9367
rect 41923 9333 41932 9367
rect 41880 9324 41932 9333
rect 43260 9324 43312 9376
rect 43352 9324 43404 9376
rect 43904 9324 43956 9376
rect 45560 9324 45612 9376
rect 46112 9324 46164 9376
rect 46848 9324 46900 9376
rect 47124 9324 47176 9376
rect 49240 9324 49292 9376
rect 50436 9367 50488 9376
rect 50436 9333 50445 9367
rect 50445 9333 50479 9367
rect 50479 9333 50488 9367
rect 50436 9324 50488 9333
rect 51172 9367 51224 9376
rect 51172 9333 51181 9367
rect 51181 9333 51215 9367
rect 51215 9333 51224 9367
rect 51172 9324 51224 9333
rect 51264 9324 51316 9376
rect 52276 9324 52328 9376
rect 53380 9324 53432 9376
rect 59636 9324 59688 9376
rect 72424 9324 72476 9376
rect 88248 9392 88300 9444
rect 92848 9460 92900 9512
rect 93400 9460 93452 9512
rect 96160 9528 96212 9580
rect 96804 9528 96856 9580
rect 98000 9571 98052 9580
rect 98000 9537 98009 9571
rect 98009 9537 98043 9571
rect 98043 9537 98052 9571
rect 98000 9528 98052 9537
rect 99288 9571 99340 9580
rect 99288 9537 99297 9571
rect 99297 9537 99331 9571
rect 99331 9537 99340 9571
rect 99288 9528 99340 9537
rect 99472 9571 99524 9580
rect 99472 9537 99481 9571
rect 99481 9537 99515 9571
rect 99515 9537 99524 9571
rect 99472 9528 99524 9537
rect 98092 9460 98144 9512
rect 100208 9528 100260 9580
rect 103244 9571 103296 9580
rect 103244 9537 103253 9571
rect 103253 9537 103287 9571
rect 103287 9537 103296 9571
rect 103244 9528 103296 9537
rect 103888 9571 103940 9580
rect 103888 9537 103897 9571
rect 103897 9537 103931 9571
rect 103931 9537 103940 9571
rect 103888 9528 103940 9537
rect 104900 9571 104952 9580
rect 104900 9537 104909 9571
rect 104909 9537 104943 9571
rect 104943 9537 104952 9571
rect 104900 9528 104952 9537
rect 105636 9571 105688 9580
rect 105636 9537 105645 9571
rect 105645 9537 105679 9571
rect 105679 9537 105688 9571
rect 105636 9528 105688 9537
rect 106280 9528 106332 9580
rect 107752 9571 107804 9580
rect 107752 9537 107761 9571
rect 107761 9537 107795 9571
rect 107795 9537 107804 9571
rect 107752 9528 107804 9537
rect 108396 9571 108448 9580
rect 108396 9537 108405 9571
rect 108405 9537 108439 9571
rect 108439 9537 108448 9571
rect 108396 9528 108448 9537
rect 109040 9571 109092 9580
rect 109040 9537 109049 9571
rect 109049 9537 109083 9571
rect 109083 9537 109092 9571
rect 109040 9528 109092 9537
rect 110052 9571 110104 9580
rect 110052 9537 110061 9571
rect 110061 9537 110095 9571
rect 110095 9537 110104 9571
rect 110052 9528 110104 9537
rect 110788 9571 110840 9580
rect 110788 9537 110797 9571
rect 110797 9537 110831 9571
rect 110831 9537 110840 9571
rect 110788 9528 110840 9537
rect 111524 9571 111576 9580
rect 111524 9537 111533 9571
rect 111533 9537 111567 9571
rect 111567 9537 111576 9571
rect 111524 9528 111576 9537
rect 112904 9571 112956 9580
rect 112904 9537 112913 9571
rect 112913 9537 112947 9571
rect 112947 9537 112956 9571
rect 112904 9528 112956 9537
rect 113548 9571 113600 9580
rect 113548 9537 113557 9571
rect 113557 9537 113591 9571
rect 113591 9537 113600 9571
rect 113548 9528 113600 9537
rect 114192 9571 114244 9580
rect 114192 9537 114201 9571
rect 114201 9537 114235 9571
rect 114235 9537 114244 9571
rect 114192 9528 114244 9537
rect 115204 9571 115256 9580
rect 115204 9537 115213 9571
rect 115213 9537 115247 9571
rect 115247 9537 115256 9571
rect 115204 9528 115256 9537
rect 115940 9571 115992 9580
rect 115940 9537 115949 9571
rect 115949 9537 115983 9571
rect 115983 9537 115992 9571
rect 115940 9528 115992 9537
rect 116676 9571 116728 9580
rect 116676 9537 116685 9571
rect 116685 9537 116719 9571
rect 116719 9537 116728 9571
rect 116676 9528 116728 9537
rect 118056 9571 118108 9580
rect 118056 9537 118065 9571
rect 118065 9537 118099 9571
rect 118099 9537 118108 9571
rect 118056 9528 118108 9537
rect 118700 9571 118752 9580
rect 118700 9537 118709 9571
rect 118709 9537 118743 9571
rect 118743 9537 118752 9571
rect 118700 9528 118752 9537
rect 119344 9571 119396 9580
rect 119344 9537 119353 9571
rect 119353 9537 119387 9571
rect 119387 9537 119396 9571
rect 119344 9528 119396 9537
rect 120356 9571 120408 9580
rect 120356 9537 120365 9571
rect 120365 9537 120399 9571
rect 120399 9537 120408 9571
rect 120356 9528 120408 9537
rect 121092 9571 121144 9580
rect 121092 9537 121101 9571
rect 121101 9537 121135 9571
rect 121135 9537 121144 9571
rect 121092 9528 121144 9537
rect 121276 9460 121328 9512
rect 121460 9460 121512 9512
rect 87788 9324 87840 9376
rect 88800 9324 88852 9376
rect 111708 9392 111760 9444
rect 111892 9392 111944 9444
rect 114284 9392 114336 9444
rect 92204 9324 92256 9376
rect 93216 9324 93268 9376
rect 94320 9324 94372 9376
rect 94964 9324 95016 9376
rect 98276 9324 98328 9376
rect 99380 9324 99432 9376
rect 100392 9324 100444 9376
rect 107568 9367 107620 9376
rect 107568 9333 107577 9367
rect 107577 9333 107611 9367
rect 107611 9333 107620 9367
rect 107568 9324 107620 9333
rect 108212 9367 108264 9376
rect 108212 9333 108221 9367
rect 108221 9333 108255 9367
rect 108255 9333 108264 9367
rect 108212 9324 108264 9333
rect 109868 9367 109920 9376
rect 109868 9333 109877 9367
rect 109877 9333 109911 9367
rect 109911 9333 109920 9367
rect 109868 9324 109920 9333
rect 110604 9367 110656 9376
rect 110604 9333 110613 9367
rect 110613 9333 110647 9367
rect 110647 9333 110656 9367
rect 110604 9324 110656 9333
rect 112720 9367 112772 9376
rect 112720 9333 112729 9367
rect 112729 9333 112763 9367
rect 112763 9333 112772 9367
rect 112720 9324 112772 9333
rect 113364 9367 113416 9376
rect 113364 9333 113373 9367
rect 113373 9333 113407 9367
rect 113407 9333 113416 9367
rect 113364 9324 113416 9333
rect 115020 9367 115072 9376
rect 115020 9333 115029 9367
rect 115029 9333 115063 9367
rect 115063 9333 115072 9367
rect 115020 9324 115072 9333
rect 115664 9392 115716 9444
rect 115848 9324 115900 9376
rect 118332 9324 118384 9376
rect 119160 9367 119212 9376
rect 119160 9333 119169 9367
rect 119169 9333 119203 9367
rect 119203 9333 119212 9367
rect 119160 9324 119212 9333
rect 120172 9367 120224 9376
rect 120172 9333 120181 9367
rect 120181 9333 120215 9367
rect 120215 9333 120224 9367
rect 120172 9324 120224 9333
rect 121000 9324 121052 9376
rect 121736 9324 121788 9376
rect 122472 9571 122524 9580
rect 122472 9537 122481 9571
rect 122481 9537 122515 9571
rect 122515 9537 122524 9571
rect 122472 9528 122524 9537
rect 122656 9707 122708 9716
rect 122656 9673 122665 9707
rect 122665 9673 122699 9707
rect 122699 9673 122708 9707
rect 122656 9664 122708 9673
rect 125232 9707 125284 9716
rect 125232 9673 125241 9707
rect 125241 9673 125275 9707
rect 125275 9673 125284 9707
rect 125232 9664 125284 9673
rect 127900 9707 127952 9716
rect 127900 9673 127909 9707
rect 127909 9673 127943 9707
rect 127943 9673 127952 9707
rect 127900 9664 127952 9673
rect 128820 9707 128872 9716
rect 128820 9673 128829 9707
rect 128829 9673 128863 9707
rect 128863 9673 128872 9707
rect 128820 9664 128872 9673
rect 129648 9664 129700 9716
rect 131488 9707 131540 9716
rect 131488 9673 131497 9707
rect 131497 9673 131531 9707
rect 131531 9673 131540 9707
rect 131488 9664 131540 9673
rect 133512 9707 133564 9716
rect 133512 9673 133521 9707
rect 133521 9673 133555 9707
rect 133555 9673 133564 9707
rect 133512 9664 133564 9673
rect 134248 9707 134300 9716
rect 134248 9673 134257 9707
rect 134257 9673 134291 9707
rect 134291 9673 134300 9707
rect 134248 9664 134300 9673
rect 137284 9664 137336 9716
rect 152464 9664 152516 9716
rect 155868 9664 155920 9716
rect 155960 9664 156012 9716
rect 156880 9707 156932 9716
rect 156880 9673 156889 9707
rect 156889 9673 156923 9707
rect 156923 9673 156932 9707
rect 156880 9664 156932 9673
rect 157248 9664 157300 9716
rect 157984 9664 158036 9716
rect 159456 9664 159508 9716
rect 162308 9664 162360 9716
rect 163872 9664 163924 9716
rect 124588 9528 124640 9580
rect 127992 9528 128044 9580
rect 128636 9571 128688 9580
rect 128636 9537 128645 9571
rect 128645 9537 128679 9571
rect 128679 9537 128688 9571
rect 128636 9528 128688 9537
rect 146392 9596 146444 9648
rect 129464 9528 129516 9580
rect 125876 9460 125928 9512
rect 130384 9571 130436 9580
rect 130384 9537 130393 9571
rect 130393 9537 130427 9571
rect 130427 9537 130436 9571
rect 130384 9528 130436 9537
rect 131396 9528 131448 9580
rect 133420 9528 133472 9580
rect 134248 9528 134300 9580
rect 137376 9528 137428 9580
rect 138756 9571 138808 9580
rect 138756 9537 138765 9571
rect 138765 9537 138799 9571
rect 138799 9537 138808 9571
rect 138756 9528 138808 9537
rect 138848 9528 138900 9580
rect 140688 9571 140740 9580
rect 140688 9537 140697 9571
rect 140697 9537 140731 9571
rect 140731 9537 140740 9571
rect 140688 9528 140740 9537
rect 141332 9571 141384 9580
rect 141332 9537 141341 9571
rect 141341 9537 141375 9571
rect 141375 9537 141384 9571
rect 141332 9528 141384 9537
rect 141976 9571 142028 9580
rect 141976 9537 141985 9571
rect 141985 9537 142019 9571
rect 142019 9537 142028 9571
rect 141976 9528 142028 9537
rect 143264 9571 143316 9580
rect 143264 9537 143273 9571
rect 143273 9537 143307 9571
rect 143307 9537 143316 9571
rect 143264 9528 143316 9537
rect 143356 9528 143408 9580
rect 144552 9571 144604 9580
rect 144552 9537 144561 9571
rect 144561 9537 144595 9571
rect 144595 9537 144604 9571
rect 144552 9528 144604 9537
rect 145840 9571 145892 9580
rect 145840 9537 145849 9571
rect 145849 9537 145883 9571
rect 145883 9537 145892 9571
rect 145840 9528 145892 9537
rect 146208 9528 146260 9580
rect 147128 9571 147180 9580
rect 147128 9537 147137 9571
rect 147137 9537 147171 9571
rect 147171 9537 147180 9571
rect 147128 9528 147180 9537
rect 148416 9571 148468 9580
rect 148416 9537 148425 9571
rect 148425 9537 148459 9571
rect 148459 9537 148468 9571
rect 148416 9528 148468 9537
rect 148508 9528 148560 9580
rect 149704 9571 149756 9580
rect 149704 9537 149713 9571
rect 149713 9537 149747 9571
rect 149747 9537 149756 9571
rect 149704 9528 149756 9537
rect 150992 9571 151044 9580
rect 150992 9537 151001 9571
rect 151001 9537 151035 9571
rect 151035 9537 151044 9571
rect 150992 9528 151044 9537
rect 151636 9571 151688 9580
rect 151636 9537 151645 9571
rect 151645 9537 151679 9571
rect 151679 9537 151688 9571
rect 151636 9528 151688 9537
rect 152280 9571 152332 9580
rect 152280 9537 152289 9571
rect 152289 9537 152323 9571
rect 152323 9537 152332 9571
rect 152280 9528 152332 9537
rect 153200 9528 153252 9580
rect 154212 9571 154264 9580
rect 154212 9537 154221 9571
rect 154221 9537 154255 9571
rect 154255 9537 154264 9571
rect 154212 9528 154264 9537
rect 154580 9528 154632 9580
rect 152372 9460 152424 9512
rect 129096 9392 129148 9444
rect 129280 9324 129332 9376
rect 137284 9324 137336 9376
rect 137744 9324 137796 9376
rect 142712 9392 142764 9444
rect 145380 9392 145432 9444
rect 145840 9392 145892 9444
rect 150532 9392 150584 9444
rect 138112 9324 138164 9376
rect 140504 9367 140556 9376
rect 140504 9333 140513 9367
rect 140513 9333 140547 9367
rect 140547 9333 140556 9367
rect 140504 9324 140556 9333
rect 142988 9324 143040 9376
rect 143264 9324 143316 9376
rect 145564 9324 145616 9376
rect 146208 9324 146260 9376
rect 146300 9367 146352 9376
rect 146300 9333 146309 9367
rect 146309 9333 146343 9367
rect 146343 9333 146352 9367
rect 146300 9324 146352 9333
rect 148232 9367 148284 9376
rect 148232 9333 148241 9367
rect 148241 9333 148275 9367
rect 148275 9333 148284 9367
rect 148232 9324 148284 9333
rect 150440 9324 150492 9376
rect 151268 9324 151320 9376
rect 151912 9324 151964 9376
rect 154580 9324 154632 9376
rect 155592 9324 155644 9376
rect 155776 9528 155828 9580
rect 156144 9528 156196 9580
rect 156972 9528 157024 9580
rect 157432 9571 157484 9580
rect 157432 9537 157441 9571
rect 157441 9537 157475 9571
rect 157475 9537 157484 9571
rect 157432 9528 157484 9537
rect 157800 9528 157852 9580
rect 159272 9571 159324 9580
rect 159272 9537 159281 9571
rect 159281 9537 159315 9571
rect 159315 9537 159324 9571
rect 159272 9528 159324 9537
rect 159364 9528 159416 9580
rect 161664 9528 161716 9580
rect 157984 9460 158036 9512
rect 155776 9392 155828 9444
rect 159456 9435 159508 9444
rect 159456 9401 159465 9435
rect 159465 9401 159499 9435
rect 159499 9401 159508 9435
rect 159456 9392 159508 9401
rect 160928 9460 160980 9512
rect 161756 9392 161808 9444
rect 162400 9596 162452 9648
rect 165804 9596 165856 9648
rect 170588 9596 170640 9648
rect 172336 9639 172388 9648
rect 172336 9605 172345 9639
rect 172345 9605 172379 9639
rect 172379 9605 172388 9639
rect 172336 9596 172388 9605
rect 172520 9639 172572 9648
rect 172520 9605 172529 9639
rect 172529 9605 172563 9639
rect 172563 9605 172572 9639
rect 172520 9596 172572 9605
rect 173072 9639 173124 9648
rect 173072 9605 173081 9639
rect 173081 9605 173115 9639
rect 173115 9605 173124 9639
rect 173072 9596 173124 9605
rect 175188 9596 175240 9648
rect 175924 9596 175976 9648
rect 162308 9571 162360 9580
rect 162308 9537 162317 9571
rect 162317 9537 162351 9571
rect 162351 9537 162360 9571
rect 162308 9528 162360 9537
rect 164332 9571 164384 9580
rect 164332 9537 164341 9571
rect 164341 9537 164375 9571
rect 164375 9537 164384 9571
rect 164332 9528 164384 9537
rect 165160 9528 165212 9580
rect 165528 9528 165580 9580
rect 168104 9571 168156 9580
rect 168104 9537 168113 9571
rect 168113 9537 168147 9571
rect 168147 9537 168156 9571
rect 168104 9528 168156 9537
rect 162768 9503 162820 9512
rect 162768 9469 162777 9503
rect 162777 9469 162811 9503
rect 162811 9469 162820 9503
rect 162768 9460 162820 9469
rect 164608 9503 164660 9512
rect 164608 9469 164617 9503
rect 164617 9469 164651 9503
rect 164651 9469 164660 9503
rect 164608 9460 164660 9469
rect 166264 9503 166316 9512
rect 166264 9469 166273 9503
rect 166273 9469 166307 9503
rect 166307 9469 166316 9503
rect 166264 9460 166316 9469
rect 167092 9503 167144 9512
rect 167092 9469 167101 9503
rect 167101 9469 167135 9503
rect 167135 9469 167144 9503
rect 167092 9460 167144 9469
rect 167552 9460 167604 9512
rect 167920 9503 167972 9512
rect 167920 9469 167929 9503
rect 167929 9469 167963 9503
rect 167963 9469 167972 9503
rect 167920 9460 167972 9469
rect 168288 9460 168340 9512
rect 169116 9503 169168 9512
rect 169116 9469 169125 9503
rect 169125 9469 169159 9503
rect 169159 9469 169168 9503
rect 169116 9460 169168 9469
rect 169300 9528 169352 9580
rect 169760 9460 169812 9512
rect 171692 9571 171744 9580
rect 171692 9537 171701 9571
rect 171701 9537 171735 9571
rect 171735 9537 171744 9571
rect 171692 9528 171744 9537
rect 174452 9571 174504 9580
rect 174452 9537 174461 9571
rect 174461 9537 174495 9571
rect 174495 9537 174504 9571
rect 174452 9528 174504 9537
rect 174728 9503 174780 9512
rect 174728 9469 174737 9503
rect 174737 9469 174771 9503
rect 174771 9469 174780 9503
rect 174728 9460 174780 9469
rect 177948 9528 178000 9580
rect 179144 9571 179196 9580
rect 179144 9537 179153 9571
rect 179153 9537 179187 9571
rect 179187 9537 179196 9571
rect 179144 9528 179196 9537
rect 179972 9664 180024 9716
rect 181720 9571 181772 9580
rect 181720 9537 181729 9571
rect 181729 9537 181763 9571
rect 181763 9537 181772 9571
rect 181720 9528 181772 9537
rect 181996 9571 182048 9580
rect 181996 9537 182005 9571
rect 182005 9537 182039 9571
rect 182039 9537 182048 9571
rect 181996 9528 182048 9537
rect 182548 9528 182600 9580
rect 185492 9528 185544 9580
rect 187700 9528 187752 9580
rect 190000 9528 190052 9580
rect 190828 9571 190880 9580
rect 190828 9537 190837 9571
rect 190837 9537 190871 9571
rect 190871 9537 190880 9571
rect 190828 9528 190880 9537
rect 192392 9571 192444 9580
rect 192392 9537 192401 9571
rect 192401 9537 192435 9571
rect 192435 9537 192444 9571
rect 192392 9528 192444 9537
rect 178040 9503 178092 9512
rect 178040 9469 178049 9503
rect 178049 9469 178083 9503
rect 178083 9469 178092 9503
rect 178040 9460 178092 9469
rect 184572 9503 184624 9512
rect 184572 9469 184581 9503
rect 184581 9469 184615 9503
rect 184615 9469 184624 9503
rect 184572 9460 184624 9469
rect 185952 9392 186004 9444
rect 157708 9324 157760 9376
rect 161112 9324 161164 9376
rect 161848 9324 161900 9376
rect 165804 9324 165856 9376
rect 166172 9324 166224 9376
rect 167460 9367 167512 9376
rect 167460 9333 167469 9367
rect 167469 9333 167503 9367
rect 167503 9333 167512 9367
rect 167460 9324 167512 9333
rect 168840 9324 168892 9376
rect 173164 9367 173216 9376
rect 173164 9333 173173 9367
rect 173173 9333 173207 9367
rect 173207 9333 173216 9367
rect 173164 9324 173216 9333
rect 175924 9367 175976 9376
rect 175924 9333 175933 9367
rect 175933 9333 175967 9367
rect 175967 9333 175976 9367
rect 175924 9324 175976 9333
rect 177948 9324 178000 9376
rect 189724 9503 189776 9512
rect 189724 9469 189733 9503
rect 189733 9469 189767 9503
rect 189767 9469 189776 9503
rect 189724 9460 189776 9469
rect 192576 9707 192628 9716
rect 192576 9673 192585 9707
rect 192585 9673 192619 9707
rect 192619 9673 192628 9707
rect 192576 9664 192628 9673
rect 192852 9664 192904 9716
rect 194324 9664 194376 9716
rect 195796 9664 195848 9716
rect 196532 9664 196584 9716
rect 198004 9664 198056 9716
rect 200028 9707 200080 9716
rect 200028 9673 200037 9707
rect 200037 9673 200071 9707
rect 200071 9673 200080 9707
rect 200028 9664 200080 9673
rect 200120 9664 200172 9716
rect 202512 9707 202564 9716
rect 202512 9673 202521 9707
rect 202521 9673 202555 9707
rect 202555 9673 202564 9707
rect 202512 9664 202564 9673
rect 202604 9664 202656 9716
rect 209596 9664 209648 9716
rect 212540 9664 212592 9716
rect 210792 9596 210844 9648
rect 212724 9664 212776 9716
rect 224316 9664 224368 9716
rect 225696 9707 225748 9716
rect 225696 9673 225705 9707
rect 225705 9673 225739 9707
rect 225739 9673 225748 9707
rect 225696 9664 225748 9673
rect 227536 9664 227588 9716
rect 229100 9664 229152 9716
rect 229192 9664 229244 9716
rect 193588 9528 193640 9580
rect 195796 9528 195848 9580
rect 196624 9528 196676 9580
rect 197544 9528 197596 9580
rect 197912 9571 197964 9580
rect 197912 9537 197921 9571
rect 197921 9537 197955 9571
rect 197955 9537 197964 9571
rect 197912 9528 197964 9537
rect 198832 9528 198884 9580
rect 199844 9571 199896 9580
rect 199844 9537 199853 9571
rect 199853 9537 199887 9571
rect 199887 9537 199896 9571
rect 199844 9528 199896 9537
rect 194416 9460 194468 9512
rect 194600 9460 194652 9512
rect 202696 9528 202748 9580
rect 203432 9528 203484 9580
rect 205824 9571 205876 9580
rect 205824 9537 205833 9571
rect 205833 9537 205867 9571
rect 205867 9537 205876 9571
rect 205824 9528 205876 9537
rect 206560 9571 206612 9580
rect 206560 9537 206569 9571
rect 206569 9537 206603 9571
rect 206603 9537 206612 9571
rect 206560 9528 206612 9537
rect 207664 9571 207716 9580
rect 207664 9537 207673 9571
rect 207673 9537 207707 9571
rect 207707 9537 207716 9571
rect 207664 9528 207716 9537
rect 208308 9571 208360 9580
rect 208308 9537 208317 9571
rect 208317 9537 208351 9571
rect 208351 9537 208360 9571
rect 208308 9528 208360 9537
rect 208952 9571 209004 9580
rect 208952 9537 208961 9571
rect 208961 9537 208995 9571
rect 208995 9537 209004 9571
rect 208952 9528 209004 9537
rect 209320 9528 209372 9580
rect 210884 9571 210936 9580
rect 210884 9537 210893 9571
rect 210893 9537 210927 9571
rect 210927 9537 210936 9571
rect 210884 9528 210936 9537
rect 214932 9596 214984 9648
rect 229836 9707 229888 9716
rect 229836 9673 229845 9707
rect 229845 9673 229879 9707
rect 229879 9673 229888 9707
rect 229836 9664 229888 9673
rect 230664 9664 230716 9716
rect 212540 9528 212592 9580
rect 213460 9571 213512 9580
rect 213460 9537 213469 9571
rect 213469 9537 213503 9571
rect 213503 9537 213512 9571
rect 213460 9528 213512 9537
rect 213920 9528 213972 9580
rect 214380 9528 214432 9580
rect 215300 9528 215352 9580
rect 215484 9528 215536 9580
rect 216680 9571 216732 9580
rect 216680 9537 216689 9571
rect 216689 9537 216723 9571
rect 216723 9537 216732 9571
rect 216680 9528 216732 9537
rect 217968 9571 218020 9580
rect 217968 9537 217977 9571
rect 217977 9537 218011 9571
rect 218011 9537 218020 9571
rect 217968 9528 218020 9537
rect 218612 9571 218664 9580
rect 218612 9537 218621 9571
rect 218621 9537 218655 9571
rect 218655 9537 218664 9571
rect 218612 9528 218664 9537
rect 219256 9571 219308 9580
rect 219256 9537 219265 9571
rect 219265 9537 219299 9571
rect 219299 9537 219308 9571
rect 219256 9528 219308 9537
rect 220544 9571 220596 9580
rect 220544 9537 220553 9571
rect 220553 9537 220587 9571
rect 220587 9537 220596 9571
rect 220544 9528 220596 9537
rect 220820 9528 220872 9580
rect 221832 9571 221884 9580
rect 221832 9537 221841 9571
rect 221841 9537 221875 9571
rect 221875 9537 221884 9571
rect 221832 9528 221884 9537
rect 223120 9571 223172 9580
rect 223120 9537 223129 9571
rect 223129 9537 223163 9571
rect 223163 9537 223172 9571
rect 223120 9528 223172 9537
rect 223304 9528 223356 9580
rect 224316 9528 224368 9580
rect 218244 9460 218296 9512
rect 197268 9392 197320 9444
rect 198188 9392 198240 9444
rect 224408 9460 224460 9512
rect 224592 9571 224644 9580
rect 224592 9537 224601 9571
rect 224601 9537 224635 9571
rect 224635 9537 224644 9571
rect 224592 9528 224644 9537
rect 224776 9571 224828 9580
rect 224776 9537 224785 9571
rect 224785 9537 224819 9571
rect 224819 9537 224828 9571
rect 224776 9528 224828 9537
rect 228364 9528 228416 9580
rect 229468 9460 229520 9512
rect 232872 9596 232924 9648
rect 233516 9707 233568 9716
rect 233516 9673 233525 9707
rect 233525 9673 233559 9707
rect 233559 9673 233568 9707
rect 233516 9664 233568 9673
rect 234344 9707 234396 9716
rect 234344 9673 234353 9707
rect 234353 9673 234387 9707
rect 234387 9673 234396 9707
rect 234344 9664 234396 9673
rect 235080 9707 235132 9716
rect 235080 9673 235089 9707
rect 235089 9673 235123 9707
rect 235123 9673 235132 9707
rect 235080 9664 235132 9673
rect 235816 9664 235868 9716
rect 236552 9664 236604 9716
rect 240232 9639 240284 9648
rect 240232 9605 240241 9639
rect 240241 9605 240275 9639
rect 240275 9605 240284 9639
rect 240232 9596 240284 9605
rect 255688 9707 255740 9716
rect 255688 9673 255697 9707
rect 255697 9673 255731 9707
rect 255731 9673 255740 9707
rect 255688 9664 255740 9673
rect 258448 9664 258500 9716
rect 259920 9664 259972 9716
rect 260012 9707 260064 9716
rect 260012 9673 260021 9707
rect 260021 9673 260055 9707
rect 260055 9673 260064 9707
rect 260012 9664 260064 9673
rect 262128 9664 262180 9716
rect 262220 9664 262272 9716
rect 262864 9707 262916 9716
rect 262864 9673 262873 9707
rect 262873 9673 262907 9707
rect 262907 9673 262916 9707
rect 262864 9664 262916 9673
rect 263140 9664 263192 9716
rect 230020 9528 230072 9580
rect 230204 9528 230256 9580
rect 231032 9528 231084 9580
rect 234068 9528 234120 9580
rect 234160 9571 234212 9580
rect 234160 9537 234169 9571
rect 234169 9537 234203 9571
rect 234203 9537 234212 9571
rect 234160 9528 234212 9537
rect 234896 9571 234948 9580
rect 234896 9537 234905 9571
rect 234905 9537 234939 9571
rect 234939 9537 234948 9571
rect 234896 9528 234948 9537
rect 235816 9571 235868 9580
rect 235816 9537 235825 9571
rect 235825 9537 235859 9571
rect 235859 9537 235868 9571
rect 235816 9528 235868 9537
rect 235908 9528 235960 9580
rect 239680 9571 239732 9580
rect 239680 9537 239689 9571
rect 239689 9537 239723 9571
rect 239723 9537 239732 9571
rect 239680 9528 239732 9537
rect 241244 9571 241296 9580
rect 241244 9537 241253 9571
rect 241253 9537 241287 9571
rect 241287 9537 241296 9571
rect 241244 9528 241296 9537
rect 235448 9460 235500 9512
rect 219164 9392 219216 9444
rect 222108 9392 222160 9444
rect 222200 9392 222252 9444
rect 234620 9392 234672 9444
rect 235540 9392 235592 9444
rect 241520 9503 241572 9512
rect 241520 9469 241529 9503
rect 241529 9469 241563 9503
rect 241563 9469 241572 9503
rect 241520 9460 241572 9469
rect 242716 9528 242768 9580
rect 244924 9528 244976 9580
rect 247868 9528 247920 9580
rect 250076 9528 250128 9580
rect 253112 9528 253164 9580
rect 255872 9571 255924 9580
rect 255872 9537 255881 9571
rect 255881 9537 255915 9571
rect 255915 9537 255924 9571
rect 255872 9528 255924 9537
rect 257896 9571 257948 9580
rect 257896 9537 257905 9571
rect 257905 9537 257939 9571
rect 257939 9537 257948 9571
rect 257896 9528 257948 9537
rect 259184 9571 259236 9580
rect 259184 9537 259193 9571
rect 259193 9537 259227 9571
rect 259227 9537 259236 9571
rect 259184 9528 259236 9537
rect 259920 9528 259972 9580
rect 260656 9571 260708 9580
rect 260656 9537 260665 9571
rect 260665 9537 260699 9571
rect 260699 9537 260708 9571
rect 260656 9528 260708 9537
rect 261208 9528 261260 9580
rect 264704 9596 264756 9648
rect 268108 9596 268160 9648
rect 262864 9528 262916 9580
rect 263968 9528 264020 9580
rect 265072 9528 265124 9580
rect 265992 9571 266044 9580
rect 265992 9537 266001 9571
rect 266001 9537 266035 9571
rect 266035 9537 266044 9571
rect 265992 9528 266044 9537
rect 267832 9528 267884 9580
rect 268844 9528 268896 9580
rect 269488 9571 269540 9580
rect 269488 9537 269497 9571
rect 269497 9537 269531 9571
rect 269531 9537 269540 9571
rect 269488 9528 269540 9537
rect 271236 9528 271288 9580
rect 190920 9367 190972 9376
rect 190920 9333 190929 9367
rect 190929 9333 190963 9367
rect 190963 9333 190972 9367
rect 190920 9324 190972 9333
rect 195520 9324 195572 9376
rect 200672 9324 200724 9376
rect 207388 9324 207440 9376
rect 208124 9367 208176 9376
rect 208124 9333 208133 9367
rect 208133 9333 208167 9367
rect 208167 9333 208176 9367
rect 208124 9324 208176 9333
rect 208768 9367 208820 9376
rect 208768 9333 208777 9367
rect 208777 9333 208811 9367
rect 208811 9333 208820 9367
rect 208768 9324 208820 9333
rect 210056 9367 210108 9376
rect 210056 9333 210065 9367
rect 210065 9333 210099 9367
rect 210099 9333 210108 9367
rect 210056 9324 210108 9333
rect 211252 9324 211304 9376
rect 212724 9324 212776 9376
rect 213276 9367 213328 9376
rect 213276 9333 213285 9367
rect 213285 9333 213319 9367
rect 213319 9333 213328 9367
rect 213276 9324 213328 9333
rect 213920 9367 213972 9376
rect 213920 9333 213929 9367
rect 213929 9333 213963 9367
rect 213963 9333 213972 9367
rect 213920 9324 213972 9333
rect 214472 9324 214524 9376
rect 215392 9324 215444 9376
rect 217692 9324 217744 9376
rect 217784 9367 217836 9376
rect 217784 9333 217793 9367
rect 217793 9333 217827 9367
rect 217827 9333 217836 9367
rect 217784 9324 217836 9333
rect 219348 9324 219400 9376
rect 220360 9367 220412 9376
rect 220360 9333 220369 9367
rect 220369 9333 220403 9367
rect 220403 9333 220412 9367
rect 220360 9324 220412 9333
rect 222844 9324 222896 9376
rect 222936 9367 222988 9376
rect 222936 9333 222945 9367
rect 222945 9333 222979 9367
rect 222979 9333 222988 9367
rect 222936 9324 222988 9333
rect 225144 9324 225196 9376
rect 225696 9324 225748 9376
rect 228088 9324 228140 9376
rect 228272 9324 228324 9376
rect 229836 9324 229888 9376
rect 231584 9367 231636 9376
rect 231584 9333 231593 9367
rect 231593 9333 231627 9367
rect 231627 9333 231636 9367
rect 231584 9324 231636 9333
rect 232872 9324 232924 9376
rect 243544 9392 243596 9444
rect 243820 9503 243872 9512
rect 243820 9469 243829 9503
rect 243829 9469 243863 9503
rect 243863 9469 243872 9503
rect 243820 9460 243872 9469
rect 245660 9460 245712 9512
rect 248972 9503 249024 9512
rect 248972 9469 248981 9503
rect 248981 9469 249015 9503
rect 249015 9469 249024 9503
rect 248972 9460 249024 9469
rect 251456 9460 251508 9512
rect 254032 9460 254084 9512
rect 255228 9460 255280 9512
rect 256792 9460 256844 9512
rect 258172 9460 258224 9512
rect 246672 9392 246724 9444
rect 246764 9392 246816 9444
rect 257988 9392 258040 9444
rect 236184 9367 236236 9376
rect 236184 9333 236193 9367
rect 236193 9333 236227 9367
rect 236227 9333 236236 9367
rect 236184 9324 236236 9333
rect 236552 9367 236604 9376
rect 236552 9333 236561 9367
rect 236561 9333 236595 9367
rect 236595 9333 236604 9367
rect 236552 9324 236604 9333
rect 237196 9324 237248 9376
rect 238116 9324 238168 9376
rect 243176 9324 243228 9376
rect 254124 9324 254176 9376
rect 258080 9324 258132 9376
rect 258724 9460 258776 9512
rect 261484 9460 261536 9512
rect 262128 9460 262180 9512
rect 265348 9460 265400 9512
rect 265900 9460 265952 9512
rect 266728 9460 266780 9512
rect 267648 9460 267700 9512
rect 268476 9460 268528 9512
rect 268660 9460 268712 9512
rect 270408 9503 270460 9512
rect 270408 9469 270417 9503
rect 270417 9469 270451 9503
rect 270451 9469 270460 9503
rect 270408 9460 270460 9469
rect 263692 9392 263744 9444
rect 261484 9324 261536 9376
rect 261576 9324 261628 9376
rect 262036 9324 262088 9376
rect 263784 9324 263836 9376
rect 264060 9324 264112 9376
rect 265532 9324 265584 9376
rect 265624 9324 265676 9376
rect 267004 9324 267056 9376
rect 268200 9324 268252 9376
rect 269304 9324 269356 9376
rect 269856 9324 269908 9376
rect 270408 9324 270460 9376
rect 34748 9222 34800 9274
rect 34812 9222 34864 9274
rect 34876 9222 34928 9274
rect 34940 9222 34992 9274
rect 35004 9222 35056 9274
rect 102345 9222 102397 9274
rect 102409 9222 102461 9274
rect 102473 9222 102525 9274
rect 102537 9222 102589 9274
rect 102601 9222 102653 9274
rect 169942 9222 169994 9274
rect 170006 9222 170058 9274
rect 170070 9222 170122 9274
rect 170134 9222 170186 9274
rect 170198 9222 170250 9274
rect 237539 9222 237591 9274
rect 237603 9222 237655 9274
rect 237667 9222 237719 9274
rect 237731 9222 237783 9274
rect 237795 9222 237847 9274
rect 1400 9120 1452 9172
rect 2412 9120 2464 9172
rect 23112 9120 23164 9172
rect 25136 9120 25188 9172
rect 27712 9120 27764 9172
rect 12808 9052 12860 9104
rect 31300 9052 31352 9104
rect 2504 8984 2556 9036
rect 22744 8984 22796 9036
rect 22836 9027 22888 9036
rect 22836 8993 22845 9027
rect 22845 8993 22879 9027
rect 22879 8993 22888 9027
rect 22836 8984 22888 8993
rect 23940 8984 23992 9036
rect 24860 8984 24912 9036
rect 3148 8959 3200 8968
rect 3148 8925 3157 8959
rect 3157 8925 3191 8959
rect 3191 8925 3200 8959
rect 3148 8916 3200 8925
rect 8208 8916 8260 8968
rect 10508 8959 10560 8968
rect 10508 8925 10517 8959
rect 10517 8925 10551 8959
rect 10551 8925 10560 8959
rect 10508 8916 10560 8925
rect 11244 8959 11296 8968
rect 11244 8925 11253 8959
rect 11253 8925 11287 8959
rect 11287 8925 11296 8959
rect 11244 8916 11296 8925
rect 13452 8959 13504 8968
rect 13452 8925 13461 8959
rect 13461 8925 13495 8959
rect 13495 8925 13504 8959
rect 13452 8916 13504 8925
rect 23848 8959 23900 8968
rect 23848 8925 23857 8959
rect 23857 8925 23891 8959
rect 23891 8925 23900 8959
rect 23848 8916 23900 8925
rect 24124 8916 24176 8968
rect 25044 8916 25096 8968
rect 26240 8984 26292 9036
rect 31760 9120 31812 9172
rect 35164 9163 35216 9172
rect 35164 9129 35173 9163
rect 35173 9129 35207 9163
rect 35207 9129 35216 9163
rect 35164 9120 35216 9129
rect 41236 9120 41288 9172
rect 41880 9120 41932 9172
rect 53196 9163 53248 9172
rect 53196 9129 53205 9163
rect 53205 9129 53239 9163
rect 53239 9129 53248 9163
rect 53196 9120 53248 9129
rect 31484 9052 31536 9104
rect 45928 9052 45980 9104
rect 46204 9052 46256 9104
rect 56416 9120 56468 9172
rect 57520 9163 57572 9172
rect 57520 9129 57529 9163
rect 57529 9129 57563 9163
rect 57563 9129 57572 9163
rect 57520 9120 57572 9129
rect 59176 9163 59228 9172
rect 59176 9129 59185 9163
rect 59185 9129 59219 9163
rect 59219 9129 59228 9163
rect 59176 9120 59228 9129
rect 60004 9163 60056 9172
rect 60004 9129 60013 9163
rect 60013 9129 60047 9163
rect 60047 9129 60056 9163
rect 60004 9120 60056 9129
rect 62764 9163 62816 9172
rect 62764 9129 62773 9163
rect 62773 9129 62807 9163
rect 62807 9129 62816 9163
rect 62764 9120 62816 9129
rect 64052 9120 64104 9172
rect 55404 9052 55456 9104
rect 64696 9052 64748 9104
rect 66352 9163 66404 9172
rect 66352 9129 66361 9163
rect 66361 9129 66395 9163
rect 66395 9129 66404 9163
rect 66352 9120 66404 9129
rect 67272 9120 67324 9172
rect 88248 9120 88300 9172
rect 88340 9120 88392 9172
rect 90180 9163 90232 9172
rect 90180 9129 90189 9163
rect 90189 9129 90223 9163
rect 90223 9129 90232 9163
rect 90180 9120 90232 9129
rect 96160 9163 96212 9172
rect 96160 9129 96169 9163
rect 96169 9129 96203 9163
rect 96203 9129 96212 9163
rect 96160 9120 96212 9129
rect 97172 9120 97224 9172
rect 98000 9163 98052 9172
rect 98000 9129 98009 9163
rect 98009 9129 98043 9163
rect 98043 9129 98052 9163
rect 98000 9120 98052 9129
rect 98092 9120 98144 9172
rect 100116 9120 100168 9172
rect 102692 9120 102744 9172
rect 107568 9120 107620 9172
rect 107660 9120 107712 9172
rect 112720 9120 112772 9172
rect 121368 9120 121420 9172
rect 122472 9120 122524 9172
rect 122748 9120 122800 9172
rect 124588 9163 124640 9172
rect 124588 9129 124597 9163
rect 124597 9129 124631 9163
rect 124631 9129 124640 9163
rect 124588 9120 124640 9129
rect 127808 9163 127860 9172
rect 127808 9129 127817 9163
rect 127817 9129 127851 9163
rect 127851 9129 127860 9163
rect 127808 9120 127860 9129
rect 131396 9163 131448 9172
rect 131396 9129 131405 9163
rect 131405 9129 131439 9163
rect 131439 9129 131448 9163
rect 131396 9120 131448 9129
rect 3332 8891 3384 8900
rect 3332 8857 3341 8891
rect 3341 8857 3375 8891
rect 3375 8857 3384 8891
rect 3332 8848 3384 8857
rect 8484 8891 8536 8900
rect 8484 8857 8493 8891
rect 8493 8857 8527 8891
rect 8527 8857 8536 8891
rect 8484 8848 8536 8857
rect 17224 8848 17276 8900
rect 21456 8848 21508 8900
rect 11336 8823 11388 8832
rect 11336 8789 11345 8823
rect 11345 8789 11379 8823
rect 11379 8789 11388 8823
rect 11336 8780 11388 8789
rect 13544 8823 13596 8832
rect 13544 8789 13553 8823
rect 13553 8789 13587 8823
rect 13587 8789 13596 8823
rect 13544 8780 13596 8789
rect 24032 8823 24084 8832
rect 24032 8789 24041 8823
rect 24041 8789 24075 8823
rect 24075 8789 24084 8823
rect 24032 8780 24084 8789
rect 25136 8891 25188 8900
rect 25136 8857 25145 8891
rect 25145 8857 25179 8891
rect 25179 8857 25188 8891
rect 25136 8848 25188 8857
rect 26424 8848 26476 8900
rect 27528 8916 27580 8968
rect 27068 8848 27120 8900
rect 29000 8959 29052 8968
rect 29000 8925 29009 8959
rect 29009 8925 29043 8959
rect 29043 8925 29052 8959
rect 29000 8916 29052 8925
rect 29552 8848 29604 8900
rect 29920 8848 29972 8900
rect 30380 8916 30432 8968
rect 31116 8959 31168 8968
rect 31116 8925 31125 8959
rect 31125 8925 31159 8959
rect 31159 8925 31168 8959
rect 31116 8916 31168 8925
rect 55864 8984 55916 9036
rect 31944 8959 31996 8968
rect 31944 8925 31953 8959
rect 31953 8925 31987 8959
rect 31987 8925 31996 8959
rect 31944 8916 31996 8925
rect 40316 8959 40368 8968
rect 40316 8925 40325 8959
rect 40325 8925 40359 8959
rect 40359 8925 40368 8959
rect 40316 8916 40368 8925
rect 45468 8959 45520 8968
rect 45468 8925 45477 8959
rect 45477 8925 45511 8959
rect 45511 8925 45520 8959
rect 45468 8916 45520 8925
rect 53380 8916 53432 8968
rect 53472 8916 53524 8968
rect 54392 8916 54444 8968
rect 37004 8848 37056 8900
rect 54024 8848 54076 8900
rect 55404 8916 55456 8968
rect 56416 8959 56468 8968
rect 56416 8925 56425 8959
rect 56425 8925 56459 8959
rect 56459 8925 56468 8959
rect 56416 8916 56468 8925
rect 57152 8959 57204 8968
rect 57152 8925 57161 8959
rect 57161 8925 57195 8959
rect 57195 8925 57204 8959
rect 57152 8916 57204 8925
rect 58900 8959 58952 8968
rect 58900 8925 58909 8959
rect 58909 8925 58943 8959
rect 58943 8925 58952 8959
rect 58900 8916 58952 8925
rect 59636 8959 59688 8968
rect 59636 8925 59645 8959
rect 59645 8925 59679 8959
rect 59679 8925 59688 8959
rect 59636 8916 59688 8925
rect 59820 8959 59872 8968
rect 59820 8925 59829 8959
rect 59829 8925 59863 8959
rect 59863 8925 59872 8959
rect 59820 8916 59872 8925
rect 58532 8848 58584 8900
rect 67180 8984 67232 9036
rect 69572 9027 69624 9036
rect 69572 8993 69581 9027
rect 69581 8993 69615 9027
rect 69615 8993 69624 9027
rect 69572 8984 69624 8993
rect 72056 9027 72108 9036
rect 72056 8993 72065 9027
rect 72065 8993 72099 9027
rect 72099 8993 72108 9027
rect 72056 8984 72108 8993
rect 73436 9027 73488 9036
rect 73436 8993 73445 9027
rect 73445 8993 73479 9027
rect 73479 8993 73488 9027
rect 73436 8984 73488 8993
rect 74724 9027 74776 9036
rect 74724 8993 74733 9027
rect 74733 8993 74767 9027
rect 74767 8993 74776 9027
rect 74724 8984 74776 8993
rect 75000 9027 75052 9036
rect 75000 8993 75009 9027
rect 75009 8993 75043 9027
rect 75043 8993 75052 9027
rect 75000 8984 75052 8993
rect 77208 9027 77260 9036
rect 77208 8993 77217 9027
rect 77217 8993 77251 9027
rect 77251 8993 77260 9027
rect 77208 8984 77260 8993
rect 77484 9027 77536 9036
rect 77484 8993 77493 9027
rect 77493 8993 77527 9027
rect 77527 8993 77536 9027
rect 77484 8984 77536 8993
rect 78588 9027 78640 9036
rect 78588 8993 78597 9027
rect 78597 8993 78631 9027
rect 78631 8993 78640 9027
rect 78588 8984 78640 8993
rect 79968 8984 80020 9036
rect 82360 9027 82412 9036
rect 82360 8993 82369 9027
rect 82369 8993 82403 9027
rect 82403 8993 82412 9027
rect 82360 8984 82412 8993
rect 83832 9027 83884 9036
rect 83832 8993 83841 9027
rect 83841 8993 83875 9027
rect 83875 8993 83884 9027
rect 83832 8984 83884 8993
rect 60096 8916 60148 8968
rect 60648 8916 60700 8968
rect 60924 8959 60976 8968
rect 60924 8925 60933 8959
rect 60933 8925 60967 8959
rect 60967 8925 60976 8959
rect 60924 8916 60976 8925
rect 61476 8916 61528 8968
rect 62396 8959 62448 8968
rect 62396 8925 62405 8959
rect 62405 8925 62439 8959
rect 62439 8925 62448 8959
rect 62396 8916 62448 8925
rect 63224 8959 63276 8968
rect 63224 8925 63233 8959
rect 63233 8925 63267 8959
rect 63267 8925 63276 8959
rect 63224 8916 63276 8925
rect 64052 8959 64104 8968
rect 64052 8925 64061 8959
rect 64061 8925 64095 8959
rect 64095 8925 64104 8959
rect 64052 8916 64104 8925
rect 64972 8959 65024 8968
rect 64972 8925 64981 8959
rect 64981 8925 65015 8959
rect 65015 8925 65024 8959
rect 64972 8916 65024 8925
rect 65984 8959 66036 8968
rect 65984 8925 65993 8959
rect 65993 8925 66027 8959
rect 66027 8925 66036 8959
rect 65984 8916 66036 8925
rect 66904 8916 66956 8968
rect 69848 8959 69900 8968
rect 69848 8925 69857 8959
rect 69857 8925 69891 8959
rect 69891 8925 69900 8959
rect 69848 8916 69900 8925
rect 26148 8823 26200 8832
rect 26148 8789 26157 8823
rect 26157 8789 26191 8823
rect 26191 8789 26200 8823
rect 26148 8780 26200 8789
rect 26884 8780 26936 8832
rect 29092 8780 29144 8832
rect 29460 8780 29512 8832
rect 30288 8780 30340 8832
rect 31116 8780 31168 8832
rect 32496 8780 32548 8832
rect 40132 8823 40184 8832
rect 40132 8789 40141 8823
rect 40141 8789 40175 8823
rect 40175 8789 40184 8823
rect 40132 8780 40184 8789
rect 43444 8780 43496 8832
rect 54576 8780 54628 8832
rect 55312 8780 55364 8832
rect 56048 8780 56100 8832
rect 56876 8780 56928 8832
rect 58440 8780 58492 8832
rect 61384 8780 61436 8832
rect 62120 8780 62172 8832
rect 63592 8823 63644 8832
rect 63592 8789 63601 8823
rect 63601 8789 63635 8823
rect 63635 8789 63644 8823
rect 63592 8780 63644 8789
rect 64420 8823 64472 8832
rect 64420 8789 64429 8823
rect 64429 8789 64463 8823
rect 64463 8789 64472 8823
rect 64420 8780 64472 8789
rect 65248 8823 65300 8832
rect 65248 8789 65257 8823
rect 65257 8789 65291 8823
rect 65291 8789 65300 8823
rect 65248 8780 65300 8789
rect 66812 8780 66864 8832
rect 73712 8959 73764 8968
rect 73712 8925 73721 8959
rect 73721 8925 73755 8959
rect 73755 8925 73764 8959
rect 73712 8916 73764 8925
rect 78864 8959 78916 8968
rect 78864 8925 78873 8959
rect 78873 8925 78907 8959
rect 78907 8925 78916 8959
rect 78864 8916 78916 8925
rect 80152 8959 80204 8968
rect 80152 8925 80161 8959
rect 80161 8925 80195 8959
rect 80195 8925 80204 8959
rect 80152 8916 80204 8925
rect 82636 8959 82688 8968
rect 82636 8925 82645 8959
rect 82645 8925 82679 8959
rect 82679 8925 82688 8959
rect 82636 8916 82688 8925
rect 72424 8848 72476 8900
rect 84108 8959 84160 8968
rect 84108 8925 84117 8959
rect 84117 8925 84151 8959
rect 84151 8925 84160 8959
rect 84108 8916 84160 8925
rect 85396 8959 85448 8968
rect 85396 8925 85405 8959
rect 85405 8925 85439 8959
rect 85439 8925 85448 8959
rect 85396 8916 85448 8925
rect 86500 8959 86552 8968
rect 86500 8925 86509 8959
rect 86509 8925 86543 8959
rect 86543 8925 86552 8959
rect 86500 8916 86552 8925
rect 85580 8891 85632 8900
rect 85580 8857 85589 8891
rect 85589 8857 85623 8891
rect 85623 8857 85632 8891
rect 85580 8848 85632 8857
rect 88984 8959 89036 8968
rect 88984 8925 88993 8959
rect 88993 8925 89027 8959
rect 89027 8925 89036 8959
rect 88984 8916 89036 8925
rect 89168 8959 89220 8968
rect 89168 8925 89177 8959
rect 89177 8925 89211 8959
rect 89211 8925 89220 8959
rect 89168 8916 89220 8925
rect 89904 8959 89956 8968
rect 89904 8925 89913 8959
rect 89913 8925 89947 8959
rect 89947 8925 89956 8959
rect 89904 8916 89956 8925
rect 90732 8959 90784 8968
rect 90732 8925 90741 8959
rect 90741 8925 90775 8959
rect 90775 8925 90784 8959
rect 90732 8916 90784 8925
rect 91008 8916 91060 8968
rect 92020 8916 92072 8968
rect 92388 8916 92440 8968
rect 94964 9027 95016 9036
rect 94964 8993 94973 9027
rect 94973 8993 95007 9027
rect 95007 8993 95016 9027
rect 94964 8984 95016 8993
rect 95056 8984 95108 9036
rect 96712 8984 96764 9036
rect 96896 8984 96948 9036
rect 93400 8959 93452 8968
rect 93400 8925 93409 8959
rect 93409 8925 93443 8959
rect 93443 8925 93452 8959
rect 93400 8916 93452 8925
rect 93492 8959 93544 8968
rect 93492 8925 93501 8959
rect 93501 8925 93535 8959
rect 93535 8925 93544 8959
rect 93492 8916 93544 8925
rect 93676 8959 93728 8968
rect 93676 8925 93685 8959
rect 93685 8925 93719 8959
rect 93719 8925 93728 8959
rect 93676 8916 93728 8925
rect 94320 8959 94372 8968
rect 94320 8925 94329 8959
rect 94329 8925 94363 8959
rect 94363 8925 94372 8959
rect 94320 8916 94372 8925
rect 86592 8823 86644 8832
rect 86592 8789 86601 8823
rect 86601 8789 86635 8823
rect 86635 8789 86644 8823
rect 86592 8780 86644 8789
rect 94228 8848 94280 8900
rect 105452 9052 105504 9104
rect 106096 9052 106148 9104
rect 121276 9052 121328 9104
rect 155500 9120 155552 9172
rect 156144 9163 156196 9172
rect 156144 9129 156153 9163
rect 156153 9129 156187 9163
rect 156187 9129 156196 9163
rect 156144 9120 156196 9129
rect 156972 9163 157024 9172
rect 156972 9129 156981 9163
rect 156981 9129 157015 9163
rect 157015 9129 157024 9163
rect 156972 9120 157024 9129
rect 157800 9163 157852 9172
rect 157800 9129 157809 9163
rect 157809 9129 157843 9163
rect 157843 9129 157852 9163
rect 157800 9120 157852 9129
rect 159824 9120 159876 9172
rect 163412 9120 163464 9172
rect 164792 9163 164844 9172
rect 164792 9129 164801 9163
rect 164801 9129 164835 9163
rect 164835 9129 164844 9163
rect 164792 9120 164844 9129
rect 169024 9120 169076 9172
rect 170588 9120 170640 9172
rect 189724 9120 189776 9172
rect 192392 9120 192444 9172
rect 195796 9163 195848 9172
rect 195796 9129 195805 9163
rect 195805 9129 195839 9163
rect 195839 9129 195848 9163
rect 195796 9120 195848 9129
rect 197912 9120 197964 9172
rect 199844 9120 199896 9172
rect 133420 9095 133472 9104
rect 133420 9061 133429 9095
rect 133429 9061 133463 9095
rect 133463 9061 133472 9095
rect 133420 9052 133472 9061
rect 133972 9052 134024 9104
rect 97632 9027 97684 9036
rect 97632 8993 97641 9027
rect 97641 8993 97675 9027
rect 97675 8993 97684 9027
rect 97632 8984 97684 8993
rect 98276 8984 98328 9036
rect 98460 9027 98512 9036
rect 98460 8993 98469 9027
rect 98469 8993 98503 9027
rect 98503 8993 98512 9027
rect 98460 8984 98512 8993
rect 99288 9027 99340 9036
rect 99288 8993 99297 9027
rect 99297 8993 99331 9027
rect 99331 8993 99340 9027
rect 99288 8984 99340 8993
rect 100024 8984 100076 9036
rect 104348 8984 104400 9036
rect 108212 8984 108264 9036
rect 99472 8959 99524 8968
rect 96620 8848 96672 8900
rect 99472 8925 99481 8959
rect 99481 8925 99515 8959
rect 99515 8925 99524 8959
rect 99472 8916 99524 8925
rect 100116 8959 100168 8968
rect 100116 8925 100125 8959
rect 100125 8925 100159 8959
rect 100159 8925 100168 8959
rect 100116 8916 100168 8925
rect 101680 8916 101732 8968
rect 106280 8916 106332 8968
rect 107200 8959 107252 8968
rect 107200 8925 107209 8959
rect 107209 8925 107243 8959
rect 107243 8925 107252 8959
rect 107200 8916 107252 8925
rect 112352 8959 112404 8968
rect 112352 8925 112361 8959
rect 112361 8925 112395 8959
rect 112395 8925 112404 8959
rect 112352 8916 112404 8925
rect 117320 8916 117372 8968
rect 100484 8848 100536 8900
rect 89628 8780 89680 8832
rect 90916 8780 90968 8832
rect 91652 8780 91704 8832
rect 92388 8780 92440 8832
rect 94412 8780 94464 8832
rect 95148 8780 95200 8832
rect 97264 8780 97316 8832
rect 98460 8780 98512 8832
rect 99288 8780 99340 8832
rect 99564 8780 99616 8832
rect 100668 8780 100720 8832
rect 104164 8848 104216 8900
rect 127164 8984 127216 9036
rect 120816 8959 120868 8968
rect 120816 8925 120825 8959
rect 120825 8925 120859 8959
rect 120859 8925 120868 8959
rect 120816 8916 120868 8925
rect 121644 8959 121696 8968
rect 121644 8925 121653 8959
rect 121653 8925 121687 8959
rect 121687 8925 121696 8959
rect 121644 8916 121696 8925
rect 121736 8959 121788 8968
rect 121736 8925 121745 8959
rect 121745 8925 121779 8959
rect 121779 8925 121788 8959
rect 121736 8916 121788 8925
rect 122656 8959 122708 8968
rect 122656 8925 122665 8959
rect 122665 8925 122699 8959
rect 122699 8925 122708 8959
rect 122656 8916 122708 8925
rect 123300 8916 123352 8968
rect 124128 8916 124180 8968
rect 125048 8959 125100 8968
rect 125048 8925 125057 8959
rect 125057 8925 125091 8959
rect 125091 8925 125100 8959
rect 125048 8916 125100 8925
rect 125876 8959 125928 8968
rect 125876 8925 125885 8959
rect 125885 8925 125919 8959
rect 125919 8925 125928 8959
rect 125876 8916 125928 8925
rect 126704 8959 126756 8968
rect 126704 8925 126713 8959
rect 126713 8925 126747 8959
rect 126747 8925 126756 8959
rect 126704 8916 126756 8925
rect 129280 9027 129332 9036
rect 129280 8993 129289 9027
rect 129289 8993 129323 9027
rect 129323 8993 129332 9027
rect 129280 8984 129332 8993
rect 130384 8984 130436 9036
rect 134248 9095 134300 9104
rect 134248 9061 134257 9095
rect 134257 9061 134291 9095
rect 134291 9061 134300 9095
rect 134248 9052 134300 9061
rect 134892 9095 134944 9104
rect 134892 9061 134901 9095
rect 134901 9061 134935 9095
rect 134935 9061 134944 9095
rect 134892 9052 134944 9061
rect 158352 9052 158404 9104
rect 160008 9052 160060 9104
rect 184572 9052 184624 9104
rect 128268 8916 128320 8968
rect 127808 8848 127860 8900
rect 129556 8959 129608 8968
rect 129556 8925 129565 8959
rect 129565 8925 129599 8959
rect 129599 8925 129608 8959
rect 129556 8916 129608 8925
rect 131120 8916 131172 8968
rect 131856 8959 131908 8968
rect 131856 8925 131865 8959
rect 131865 8925 131899 8959
rect 131899 8925 131908 8959
rect 131856 8916 131908 8925
rect 132960 8916 133012 8968
rect 133144 8916 133196 8968
rect 133972 8959 134024 8968
rect 133972 8925 133981 8959
rect 133981 8925 134015 8959
rect 134015 8925 134024 8959
rect 133972 8916 134024 8925
rect 134524 8916 134576 8968
rect 139768 8959 139820 8968
rect 139768 8925 139777 8959
rect 139777 8925 139811 8959
rect 139811 8925 139820 8959
rect 139768 8916 139820 8925
rect 144736 8916 144788 8968
rect 150072 8959 150124 8968
rect 150072 8925 150081 8959
rect 150081 8925 150115 8959
rect 150115 8925 150124 8959
rect 150072 8916 150124 8925
rect 155132 8959 155184 8968
rect 155132 8925 155141 8959
rect 155141 8925 155175 8959
rect 155175 8925 155184 8959
rect 155132 8916 155184 8925
rect 155684 8916 155736 8968
rect 128728 8848 128780 8900
rect 137284 8848 137336 8900
rect 137376 8848 137428 8900
rect 156696 8959 156748 8968
rect 156696 8925 156705 8959
rect 156705 8925 156739 8959
rect 156739 8925 156748 8959
rect 156696 8916 156748 8925
rect 157524 8959 157576 8968
rect 157524 8925 157533 8959
rect 157533 8925 157567 8959
rect 157567 8925 157576 8959
rect 157524 8916 157576 8925
rect 157616 8959 157668 8968
rect 157616 8925 157625 8959
rect 157625 8925 157659 8959
rect 157659 8925 157668 8959
rect 157616 8916 157668 8925
rect 158720 8848 158772 8900
rect 159640 8848 159692 8900
rect 159824 8959 159876 8968
rect 159824 8925 159833 8959
rect 159833 8925 159867 8959
rect 159867 8925 159876 8959
rect 159824 8916 159876 8925
rect 159916 8916 159968 8968
rect 160836 8959 160888 8968
rect 160836 8925 160845 8959
rect 160845 8925 160879 8959
rect 160879 8925 160888 8959
rect 160836 8916 160888 8925
rect 161204 8959 161256 8968
rect 161204 8925 161213 8959
rect 161213 8925 161247 8959
rect 161247 8925 161256 8959
rect 161204 8916 161256 8925
rect 162216 8959 162268 8968
rect 162216 8925 162225 8959
rect 162225 8925 162259 8959
rect 162259 8925 162268 8959
rect 162216 8916 162268 8925
rect 162584 8959 162636 8968
rect 162584 8925 162593 8959
rect 162593 8925 162627 8959
rect 162627 8925 162636 8959
rect 162584 8916 162636 8925
rect 164700 8916 164752 8968
rect 107108 8780 107160 8832
rect 109868 8780 109920 8832
rect 115572 8780 115624 8832
rect 123024 8780 123076 8832
rect 123760 8823 123812 8832
rect 123760 8789 123769 8823
rect 123769 8789 123803 8823
rect 123803 8789 123812 8823
rect 123760 8780 123812 8789
rect 125416 8823 125468 8832
rect 125416 8789 125425 8823
rect 125425 8789 125459 8823
rect 125459 8789 125468 8823
rect 125416 8780 125468 8789
rect 126152 8780 126204 8832
rect 126888 8780 126940 8832
rect 127164 8780 127216 8832
rect 128268 8780 128320 8832
rect 129004 8780 129056 8832
rect 132132 8780 132184 8832
rect 134248 8780 134300 8832
rect 140412 8780 140464 8832
rect 147772 8780 147824 8832
rect 149888 8823 149940 8832
rect 149888 8789 149897 8823
rect 149897 8789 149931 8823
rect 149931 8789 149940 8823
rect 149888 8780 149940 8789
rect 155500 8823 155552 8832
rect 155500 8789 155509 8823
rect 155509 8789 155543 8823
rect 155543 8789 155552 8823
rect 155500 8780 155552 8789
rect 155776 8780 155828 8832
rect 156696 8780 156748 8832
rect 157156 8780 157208 8832
rect 157248 8780 157300 8832
rect 162400 8780 162452 8832
rect 163872 8848 163924 8900
rect 164148 8891 164200 8900
rect 164148 8857 164157 8891
rect 164157 8857 164191 8891
rect 164191 8857 164200 8891
rect 164148 8848 164200 8857
rect 164240 8780 164292 8832
rect 165344 9027 165396 9036
rect 165344 8993 165353 9027
rect 165353 8993 165387 9027
rect 165387 8993 165396 9027
rect 165344 8984 165396 8993
rect 165252 8916 165304 8968
rect 177212 8984 177264 9036
rect 179604 9027 179656 9036
rect 179604 8993 179613 9027
rect 179613 8993 179647 9027
rect 179647 8993 179656 9027
rect 179604 8984 179656 8993
rect 180340 8984 180392 9036
rect 181812 8984 181864 9036
rect 182456 9027 182508 9036
rect 182456 8993 182465 9027
rect 182465 8993 182499 9027
rect 182499 8993 182508 9027
rect 182456 8984 182508 8993
rect 184296 9027 184348 9036
rect 184296 8993 184305 9027
rect 184305 8993 184339 9027
rect 184339 8993 184348 9027
rect 184296 8984 184348 8993
rect 167736 8916 167788 8968
rect 168104 8959 168156 8968
rect 168104 8925 168113 8959
rect 168113 8925 168147 8959
rect 168147 8925 168156 8959
rect 168104 8916 168156 8925
rect 168288 8916 168340 8968
rect 166264 8848 166316 8900
rect 167368 8848 167420 8900
rect 169852 8916 169904 8968
rect 169944 8916 169996 8968
rect 173716 8916 173768 8968
rect 167552 8780 167604 8832
rect 167644 8780 167696 8832
rect 176752 8891 176804 8900
rect 176752 8857 176761 8891
rect 176761 8857 176795 8891
rect 176795 8857 176804 8891
rect 176752 8848 176804 8857
rect 177488 8959 177540 8968
rect 177488 8925 177497 8959
rect 177497 8925 177531 8959
rect 177531 8925 177540 8959
rect 177488 8916 177540 8925
rect 179880 8959 179932 8968
rect 179880 8925 179889 8959
rect 179889 8925 179923 8959
rect 179923 8925 179932 8959
rect 179880 8916 179932 8925
rect 181168 8959 181220 8968
rect 181168 8925 181177 8959
rect 181177 8925 181211 8959
rect 181211 8925 181220 8959
rect 181168 8916 181220 8925
rect 184572 8959 184624 8968
rect 184572 8925 184581 8959
rect 184581 8925 184615 8959
rect 184615 8925 184624 8959
rect 184572 8916 184624 8925
rect 197176 9052 197228 9104
rect 198096 9052 198148 9104
rect 200120 9052 200172 9104
rect 184756 8984 184808 9036
rect 186228 8984 186280 9036
rect 189448 9027 189500 9036
rect 189448 8993 189457 9027
rect 189457 8993 189491 9027
rect 189491 8993 189500 9027
rect 189448 8984 189500 8993
rect 190828 8984 190880 9036
rect 185860 8959 185912 8968
rect 185860 8925 185869 8959
rect 185869 8925 185903 8959
rect 185903 8925 185912 8959
rect 185860 8916 185912 8925
rect 169852 8780 169904 8832
rect 170312 8780 170364 8832
rect 174176 8823 174228 8832
rect 174176 8789 174185 8823
rect 174185 8789 174219 8823
rect 174219 8789 174228 8823
rect 174176 8780 174228 8789
rect 176844 8823 176896 8832
rect 176844 8789 176853 8823
rect 176853 8789 176887 8823
rect 176887 8789 176896 8823
rect 176844 8780 176896 8789
rect 177580 8823 177632 8832
rect 177580 8789 177589 8823
rect 177589 8789 177623 8823
rect 177623 8789 177632 8823
rect 177580 8780 177632 8789
rect 177856 8780 177908 8832
rect 187240 8916 187292 8968
rect 190920 8916 190972 8968
rect 190828 8848 190880 8900
rect 191196 8916 191248 8968
rect 192484 8959 192536 8968
rect 192484 8925 192493 8959
rect 192493 8925 192527 8959
rect 192527 8925 192536 8959
rect 192484 8916 192536 8925
rect 193312 8959 193364 8968
rect 193312 8925 193321 8959
rect 193321 8925 193355 8959
rect 193355 8925 193364 8959
rect 193312 8916 193364 8925
rect 194600 8959 194652 8968
rect 194600 8925 194609 8959
rect 194609 8925 194643 8959
rect 194643 8925 194652 8959
rect 194600 8916 194652 8925
rect 193496 8848 193548 8900
rect 195520 8959 195572 8968
rect 195520 8925 195529 8959
rect 195529 8925 195563 8959
rect 195563 8925 195572 8959
rect 195520 8916 195572 8925
rect 196256 8959 196308 8968
rect 196256 8925 196265 8959
rect 196265 8925 196299 8959
rect 196299 8925 196308 8959
rect 196256 8916 196308 8925
rect 196532 8916 196584 8968
rect 197360 8916 197412 8968
rect 198004 8916 198056 8968
rect 198648 8959 198700 8968
rect 198648 8925 198657 8959
rect 198657 8925 198691 8959
rect 198691 8925 198700 8959
rect 198648 8916 198700 8925
rect 199660 8916 199712 8968
rect 200488 8916 200540 8968
rect 202052 9052 202104 9104
rect 203616 9052 203668 9104
rect 204076 9163 204128 9172
rect 204076 9129 204085 9163
rect 204085 9129 204119 9163
rect 204119 9129 204128 9163
rect 204076 9120 204128 9129
rect 225604 9120 225656 9172
rect 228364 9163 228416 9172
rect 228364 9129 228373 9163
rect 228373 9129 228407 9163
rect 228407 9129 228416 9163
rect 228364 9120 228416 9129
rect 228456 9120 228508 9172
rect 233792 9120 233844 9172
rect 234068 9163 234120 9172
rect 234068 9129 234077 9163
rect 234077 9129 234111 9163
rect 234111 9129 234120 9163
rect 234068 9120 234120 9129
rect 234160 9120 234212 9172
rect 236000 9120 236052 9172
rect 237288 9120 237340 9172
rect 237932 9120 237984 9172
rect 258816 9120 258868 9172
rect 260196 9163 260248 9172
rect 260196 9129 260205 9163
rect 260205 9129 260239 9163
rect 260239 9129 260248 9163
rect 260196 9120 260248 9129
rect 260656 9120 260708 9172
rect 262956 9120 263008 9172
rect 210056 9052 210108 9104
rect 212172 9052 212224 9104
rect 212356 9052 212408 9104
rect 214380 9052 214432 9104
rect 214564 9052 214616 9104
rect 222200 9052 222252 9104
rect 223488 9052 223540 9104
rect 225880 9052 225932 9104
rect 233332 9052 233384 9104
rect 233424 9052 233476 9104
rect 253940 9052 253992 9104
rect 200672 8984 200724 9036
rect 221924 8984 221976 9036
rect 201132 8916 201184 8968
rect 202052 8959 202104 8968
rect 202052 8925 202061 8959
rect 202061 8925 202095 8959
rect 202095 8925 202104 8959
rect 202052 8916 202104 8925
rect 202604 8916 202656 8968
rect 202512 8848 202564 8900
rect 203432 8959 203484 8968
rect 203432 8925 203441 8959
rect 203441 8925 203475 8959
rect 203475 8925 203484 8959
rect 203432 8916 203484 8925
rect 203524 8916 203576 8968
rect 211712 8959 211764 8968
rect 211712 8925 211721 8959
rect 211721 8925 211755 8959
rect 211755 8925 211764 8959
rect 211712 8916 211764 8925
rect 213920 8916 213972 8968
rect 215668 8916 215720 8968
rect 216864 8959 216916 8968
rect 216864 8925 216873 8959
rect 216873 8925 216907 8959
rect 216907 8925 216916 8959
rect 216864 8916 216916 8925
rect 222016 8959 222068 8968
rect 222016 8925 222025 8959
rect 222025 8925 222059 8959
rect 222059 8925 222068 8959
rect 222016 8916 222068 8925
rect 224408 8984 224460 9036
rect 224040 8959 224092 8968
rect 224040 8925 224049 8959
rect 224049 8925 224083 8959
rect 224083 8925 224092 8959
rect 224040 8916 224092 8925
rect 224684 8916 224736 8968
rect 225604 8959 225656 8968
rect 225604 8925 225613 8959
rect 225613 8925 225647 8959
rect 225647 8925 225656 8959
rect 225604 8916 225656 8925
rect 225972 8984 226024 9036
rect 226432 8959 226484 8968
rect 226432 8925 226441 8959
rect 226441 8925 226475 8959
rect 226475 8925 226484 8959
rect 226432 8916 226484 8925
rect 227260 8959 227312 8968
rect 227260 8925 227269 8959
rect 227269 8925 227303 8959
rect 227303 8925 227312 8959
rect 227260 8916 227312 8925
rect 228088 8959 228140 8968
rect 228088 8925 228097 8959
rect 228097 8925 228131 8959
rect 228131 8925 228140 8959
rect 228088 8916 228140 8925
rect 228824 8959 228876 8968
rect 228824 8925 228833 8959
rect 228833 8925 228867 8959
rect 228867 8925 228876 8959
rect 228824 8916 228876 8925
rect 230020 9027 230072 9036
rect 230020 8993 230029 9027
rect 230029 8993 230063 9027
rect 230063 8993 230072 9027
rect 230020 8984 230072 8993
rect 230848 8984 230900 9036
rect 229100 8916 229152 8968
rect 229652 8959 229704 8968
rect 229652 8925 229661 8959
rect 229661 8925 229695 8959
rect 229695 8925 229704 8959
rect 229652 8916 229704 8925
rect 229836 8959 229888 8968
rect 229836 8925 229845 8959
rect 229845 8925 229879 8959
rect 229879 8925 229888 8959
rect 229836 8916 229888 8925
rect 230204 8916 230256 8968
rect 231860 8916 231912 8968
rect 232136 8916 232188 8968
rect 232504 8916 232556 8968
rect 232872 8959 232924 8968
rect 232872 8925 232881 8959
rect 232881 8925 232915 8959
rect 232915 8925 232924 8959
rect 232872 8916 232924 8925
rect 233700 8959 233752 8968
rect 233700 8925 233709 8959
rect 233709 8925 233743 8959
rect 233743 8925 233752 8959
rect 233700 8916 233752 8925
rect 234528 8959 234580 8968
rect 234528 8925 234537 8959
rect 234537 8925 234571 8959
rect 234571 8925 234580 8959
rect 234528 8916 234580 8925
rect 236092 8984 236144 9036
rect 190368 8780 190420 8832
rect 191104 8780 191156 8832
rect 191932 8823 191984 8832
rect 191932 8789 191941 8823
rect 191941 8789 191975 8823
rect 191975 8789 191984 8823
rect 191932 8780 191984 8789
rect 192024 8780 192076 8832
rect 194048 8780 194100 8832
rect 196348 8780 196400 8832
rect 199292 8780 199344 8832
rect 201040 8780 201092 8832
rect 202420 8823 202472 8832
rect 202420 8789 202429 8823
rect 202429 8789 202463 8823
rect 202463 8789 202472 8823
rect 202420 8780 202472 8789
rect 202604 8780 202656 8832
rect 212356 8848 212408 8900
rect 212448 8848 212500 8900
rect 235632 8916 235684 8968
rect 235816 8959 235868 8968
rect 235816 8925 235825 8959
rect 235825 8925 235859 8959
rect 235859 8925 235868 8959
rect 235816 8916 235868 8925
rect 235908 8916 235960 8968
rect 241980 9027 242032 9036
rect 241980 8993 241989 9027
rect 241989 8993 242023 9027
rect 242023 8993 242032 9027
rect 241980 8984 242032 8993
rect 243452 9027 243504 9036
rect 243452 8993 243461 9027
rect 243461 8993 243495 9027
rect 243495 8993 243504 9027
rect 243452 8984 243504 8993
rect 243544 8984 243596 9036
rect 262036 9052 262088 9104
rect 263876 9052 263928 9104
rect 264704 9052 264756 9104
rect 264796 9095 264848 9104
rect 264796 9061 264805 9095
rect 264805 9061 264839 9095
rect 264839 9061 264848 9095
rect 264796 9052 264848 9061
rect 267556 9052 267608 9104
rect 254124 9027 254176 9036
rect 254124 8993 254133 9027
rect 254133 8993 254167 9027
rect 254167 8993 254176 9027
rect 254124 8984 254176 8993
rect 256424 9027 256476 9036
rect 256424 8993 256433 9027
rect 256433 8993 256467 9027
rect 256467 8993 256476 9027
rect 256424 8984 256476 8993
rect 257712 9027 257764 9036
rect 257712 8993 257721 9027
rect 257721 8993 257755 9027
rect 257755 8993 257764 9027
rect 257712 8984 257764 8993
rect 258172 8984 258224 9036
rect 238760 8916 238812 8968
rect 243728 8959 243780 8968
rect 243728 8925 243737 8959
rect 243737 8925 243771 8959
rect 243771 8925 243780 8959
rect 243728 8916 243780 8925
rect 244188 8916 244240 8968
rect 245016 8959 245068 8968
rect 245016 8925 245025 8959
rect 245025 8925 245059 8959
rect 245059 8925 245068 8959
rect 245016 8916 245068 8925
rect 246120 8959 246172 8968
rect 246120 8925 246129 8959
rect 246129 8925 246163 8959
rect 246163 8925 246172 8959
rect 246120 8916 246172 8925
rect 246212 8916 246264 8968
rect 247408 8959 247460 8968
rect 247408 8925 247417 8959
rect 247417 8925 247451 8959
rect 247451 8925 247460 8959
rect 247408 8916 247460 8925
rect 203616 8780 203668 8832
rect 211068 8780 211120 8832
rect 214380 8780 214432 8832
rect 216680 8823 216732 8832
rect 216680 8789 216689 8823
rect 216689 8789 216723 8823
rect 216723 8789 216732 8823
rect 216680 8780 216732 8789
rect 221832 8823 221884 8832
rect 221832 8789 221841 8823
rect 221841 8789 221875 8823
rect 221875 8789 221884 8823
rect 221832 8780 221884 8789
rect 221924 8780 221976 8832
rect 225696 8780 225748 8832
rect 225788 8780 225840 8832
rect 226524 8780 226576 8832
rect 228088 8780 228140 8832
rect 228916 8780 228968 8832
rect 231768 8780 231820 8832
rect 233240 8823 233292 8832
rect 233240 8789 233249 8823
rect 233249 8789 233283 8823
rect 233283 8789 233292 8823
rect 233240 8780 233292 8789
rect 233332 8780 233384 8832
rect 234068 8780 234120 8832
rect 234528 8780 234580 8832
rect 235632 8780 235684 8832
rect 236368 8780 236420 8832
rect 236552 8823 236604 8832
rect 236552 8789 236561 8823
rect 236561 8789 236595 8823
rect 236595 8789 236604 8823
rect 236552 8780 236604 8789
rect 246488 8848 246540 8900
rect 248696 8959 248748 8968
rect 248696 8925 248705 8959
rect 248705 8925 248739 8959
rect 248739 8925 248748 8959
rect 248696 8916 248748 8925
rect 247776 8848 247828 8900
rect 250812 8916 250864 8968
rect 251364 8916 251416 8968
rect 252284 8916 252336 8968
rect 252836 8959 252888 8968
rect 252836 8925 252845 8959
rect 252845 8925 252879 8959
rect 252879 8925 252888 8959
rect 252836 8916 252888 8925
rect 253848 8959 253900 8968
rect 253848 8925 253857 8959
rect 253857 8925 253891 8959
rect 253891 8925 253900 8959
rect 253848 8916 253900 8925
rect 256884 8916 256936 8968
rect 257068 8916 257120 8968
rect 258356 8916 258408 8968
rect 253940 8848 253992 8900
rect 258724 8848 258776 8900
rect 258908 8780 258960 8832
rect 259092 8891 259144 8900
rect 259092 8857 259101 8891
rect 259101 8857 259135 8891
rect 259135 8857 259144 8891
rect 259092 8848 259144 8857
rect 260104 8891 260156 8900
rect 260104 8857 260113 8891
rect 260113 8857 260147 8891
rect 260147 8857 260156 8891
rect 260104 8848 260156 8857
rect 260380 8916 260432 8968
rect 265072 8984 265124 9036
rect 265164 8984 265216 9036
rect 270592 8984 270644 9036
rect 260656 8848 260708 8900
rect 262588 8891 262640 8900
rect 262588 8857 262597 8891
rect 262597 8857 262631 8891
rect 262631 8857 262640 8891
rect 262588 8848 262640 8857
rect 263784 8916 263836 8968
rect 265808 8916 265860 8968
rect 265992 8916 266044 8968
rect 267464 8916 267516 8968
rect 268292 8916 268344 8968
rect 265164 8848 265216 8900
rect 261852 8780 261904 8832
rect 264796 8780 264848 8832
rect 266820 8891 266872 8900
rect 266820 8857 266829 8891
rect 266829 8857 266863 8891
rect 266863 8857 266872 8891
rect 266820 8848 266872 8857
rect 267188 8848 267240 8900
rect 267372 8848 267424 8900
rect 269488 8848 269540 8900
rect 270316 8916 270368 8968
rect 270408 8959 270460 8968
rect 270408 8925 270417 8959
rect 270417 8925 270451 8959
rect 270451 8925 270460 8959
rect 270408 8916 270460 8925
rect 270776 8848 270828 8900
rect 265348 8823 265400 8832
rect 265348 8789 265357 8823
rect 265357 8789 265391 8823
rect 265391 8789 265400 8823
rect 265348 8780 265400 8789
rect 266636 8780 266688 8832
rect 267740 8780 267792 8832
rect 268568 8780 268620 8832
rect 269304 8780 269356 8832
rect 271052 8780 271104 8832
rect 68546 8678 68598 8730
rect 68610 8678 68662 8730
rect 68674 8678 68726 8730
rect 68738 8678 68790 8730
rect 68802 8678 68854 8730
rect 136143 8678 136195 8730
rect 136207 8678 136259 8730
rect 136271 8678 136323 8730
rect 136335 8678 136387 8730
rect 136399 8678 136451 8730
rect 203740 8678 203792 8730
rect 203804 8678 203856 8730
rect 203868 8678 203920 8730
rect 203932 8678 203984 8730
rect 203996 8678 204048 8730
rect 271337 8678 271389 8730
rect 271401 8678 271453 8730
rect 271465 8678 271517 8730
rect 271529 8678 271581 8730
rect 271593 8678 271645 8730
rect 6920 8576 6972 8628
rect 23296 8576 23348 8628
rect 23480 8619 23532 8628
rect 23480 8585 23489 8619
rect 23489 8585 23523 8619
rect 23523 8585 23532 8619
rect 23480 8576 23532 8585
rect 23112 8508 23164 8560
rect 13544 8304 13596 8356
rect 23204 8304 23256 8356
rect 23756 8440 23808 8492
rect 25688 8508 25740 8560
rect 25964 8508 26016 8560
rect 26240 8508 26292 8560
rect 28724 8619 28776 8628
rect 28724 8585 28733 8619
rect 28733 8585 28767 8619
rect 28767 8585 28776 8619
rect 28724 8576 28776 8585
rect 29644 8619 29696 8628
rect 29644 8585 29653 8619
rect 29653 8585 29687 8619
rect 29687 8585 29696 8619
rect 29644 8576 29696 8585
rect 30196 8576 30248 8628
rect 31300 8619 31352 8628
rect 31300 8585 31309 8619
rect 31309 8585 31343 8619
rect 31343 8585 31352 8619
rect 31300 8576 31352 8585
rect 31944 8576 31996 8628
rect 32588 8576 32640 8628
rect 32680 8619 32732 8628
rect 32680 8585 32689 8619
rect 32689 8585 32723 8619
rect 32723 8585 32732 8619
rect 32680 8576 32732 8585
rect 54116 8619 54168 8628
rect 54116 8585 54125 8619
rect 54125 8585 54159 8619
rect 54159 8585 54168 8619
rect 54116 8576 54168 8585
rect 54760 8619 54812 8628
rect 54760 8585 54769 8619
rect 54769 8585 54803 8619
rect 54803 8585 54812 8619
rect 54760 8576 54812 8585
rect 55496 8619 55548 8628
rect 55496 8585 55505 8619
rect 55505 8585 55539 8619
rect 55539 8585 55548 8619
rect 55496 8576 55548 8585
rect 56232 8619 56284 8628
rect 56232 8585 56241 8619
rect 56241 8585 56275 8619
rect 56275 8585 56284 8619
rect 56232 8576 56284 8585
rect 57060 8619 57112 8628
rect 57060 8585 57069 8619
rect 57069 8585 57103 8619
rect 57103 8585 57112 8619
rect 57060 8576 57112 8585
rect 58624 8619 58676 8628
rect 58624 8585 58633 8619
rect 58633 8585 58667 8619
rect 58667 8585 58676 8619
rect 58624 8576 58676 8585
rect 59820 8619 59872 8628
rect 59820 8585 59829 8619
rect 59829 8585 59863 8619
rect 59863 8585 59872 8619
rect 59820 8576 59872 8585
rect 60740 8619 60792 8628
rect 60740 8585 60749 8619
rect 60749 8585 60783 8619
rect 60783 8585 60792 8619
rect 60740 8576 60792 8585
rect 61568 8619 61620 8628
rect 61568 8585 61577 8619
rect 61577 8585 61611 8619
rect 61611 8585 61620 8619
rect 61568 8576 61620 8585
rect 62304 8619 62356 8628
rect 62304 8585 62313 8619
rect 62313 8585 62347 8619
rect 62347 8585 62356 8619
rect 62304 8576 62356 8585
rect 63776 8619 63828 8628
rect 63776 8585 63785 8619
rect 63785 8585 63819 8619
rect 63819 8585 63828 8619
rect 63776 8576 63828 8585
rect 64604 8619 64656 8628
rect 64604 8585 64613 8619
rect 64613 8585 64647 8619
rect 64647 8585 64656 8619
rect 64604 8576 64656 8585
rect 64696 8576 64748 8628
rect 24032 8483 24084 8492
rect 24032 8449 24041 8483
rect 24041 8449 24075 8483
rect 24075 8449 24084 8483
rect 24032 8440 24084 8449
rect 24216 8415 24268 8424
rect 24216 8381 24225 8415
rect 24225 8381 24259 8415
rect 24259 8381 24268 8415
rect 24216 8372 24268 8381
rect 24860 8415 24912 8424
rect 24860 8381 24869 8415
rect 24869 8381 24903 8415
rect 24903 8381 24912 8415
rect 24860 8372 24912 8381
rect 25044 8483 25096 8492
rect 25044 8449 25053 8483
rect 25053 8449 25087 8483
rect 25087 8449 25096 8483
rect 25044 8440 25096 8449
rect 29736 8508 29788 8560
rect 28448 8483 28500 8492
rect 28448 8449 28457 8483
rect 28457 8449 28491 8483
rect 28491 8449 28500 8483
rect 28448 8440 28500 8449
rect 29000 8440 29052 8492
rect 29460 8483 29512 8492
rect 29460 8449 29469 8483
rect 29469 8449 29503 8483
rect 29503 8449 29512 8483
rect 29460 8440 29512 8449
rect 30288 8483 30340 8492
rect 30288 8449 30297 8483
rect 30297 8449 30331 8483
rect 30331 8449 30340 8483
rect 30288 8440 30340 8449
rect 31116 8483 31168 8492
rect 31116 8449 31125 8483
rect 31125 8449 31159 8483
rect 31159 8449 31168 8483
rect 31116 8440 31168 8449
rect 25228 8304 25280 8356
rect 25504 8372 25556 8424
rect 25780 8372 25832 8424
rect 36360 8508 36412 8560
rect 32496 8483 32548 8492
rect 32496 8449 32505 8483
rect 32505 8449 32539 8483
rect 32539 8449 32548 8483
rect 32496 8440 32548 8449
rect 32588 8440 32640 8492
rect 65708 8508 65760 8560
rect 65984 8508 66036 8560
rect 66996 8551 67048 8560
rect 66996 8517 67005 8551
rect 67005 8517 67039 8551
rect 67039 8517 67048 8551
rect 66996 8508 67048 8517
rect 88340 8576 88392 8628
rect 90456 8576 90508 8628
rect 91836 8619 91888 8628
rect 91836 8585 91845 8619
rect 91845 8585 91879 8619
rect 91879 8585 91888 8619
rect 91836 8576 91888 8585
rect 91928 8576 91980 8628
rect 94596 8619 94648 8628
rect 94596 8585 94605 8619
rect 94605 8585 94639 8619
rect 94639 8585 94648 8619
rect 94596 8576 94648 8585
rect 94872 8576 94924 8628
rect 96804 8619 96856 8628
rect 96804 8585 96813 8619
rect 96813 8585 96847 8619
rect 96847 8585 96856 8619
rect 96804 8576 96856 8585
rect 97448 8619 97500 8628
rect 97448 8585 97457 8619
rect 97457 8585 97491 8619
rect 97491 8585 97500 8619
rect 97448 8576 97500 8585
rect 98644 8619 98696 8628
rect 98644 8585 98653 8619
rect 98653 8585 98687 8619
rect 98687 8585 98696 8619
rect 98644 8576 98696 8585
rect 100208 8619 100260 8628
rect 100208 8585 100217 8619
rect 100217 8585 100251 8619
rect 100251 8585 100260 8619
rect 100208 8576 100260 8585
rect 100300 8576 100352 8628
rect 120816 8576 120868 8628
rect 123208 8619 123260 8628
rect 123208 8585 123217 8619
rect 123217 8585 123251 8619
rect 123251 8585 123260 8619
rect 123208 8576 123260 8585
rect 123944 8619 123996 8628
rect 123944 8585 123953 8619
rect 123953 8585 123987 8619
rect 123987 8585 123996 8619
rect 123944 8576 123996 8585
rect 125324 8576 125376 8628
rect 126336 8619 126388 8628
rect 126336 8585 126345 8619
rect 126345 8585 126379 8619
rect 126379 8585 126388 8619
rect 126336 8576 126388 8585
rect 126796 8576 126848 8628
rect 127992 8619 128044 8628
rect 127992 8585 128001 8619
rect 128001 8585 128035 8619
rect 128035 8585 128044 8619
rect 127992 8576 128044 8585
rect 128636 8576 128688 8628
rect 130476 8576 130528 8628
rect 132316 8619 132368 8628
rect 132316 8585 132325 8619
rect 132325 8585 132359 8619
rect 132359 8585 132368 8619
rect 132316 8576 132368 8585
rect 134524 8619 134576 8628
rect 134524 8585 134533 8619
rect 134533 8585 134567 8619
rect 134567 8585 134576 8619
rect 134524 8576 134576 8585
rect 137284 8576 137336 8628
rect 89996 8508 90048 8560
rect 90732 8508 90784 8560
rect 124128 8508 124180 8560
rect 125876 8508 125928 8560
rect 128728 8508 128780 8560
rect 157432 8576 157484 8628
rect 159272 8576 159324 8628
rect 159364 8619 159416 8628
rect 159364 8585 159373 8619
rect 159373 8585 159407 8619
rect 159407 8585 159416 8619
rect 159364 8576 159416 8585
rect 159824 8576 159876 8628
rect 161204 8576 161256 8628
rect 54024 8440 54076 8492
rect 54576 8483 54628 8492
rect 54576 8449 54585 8483
rect 54585 8449 54619 8483
rect 54619 8449 54628 8483
rect 54576 8440 54628 8449
rect 55312 8483 55364 8492
rect 55312 8449 55321 8483
rect 55321 8449 55355 8483
rect 55355 8449 55364 8483
rect 55312 8440 55364 8449
rect 56048 8483 56100 8492
rect 56048 8449 56057 8483
rect 56057 8449 56091 8483
rect 56091 8449 56100 8483
rect 56048 8440 56100 8449
rect 56876 8483 56928 8492
rect 56876 8449 56885 8483
rect 56885 8449 56919 8483
rect 56919 8449 56928 8483
rect 56876 8440 56928 8449
rect 58440 8483 58492 8492
rect 58440 8449 58449 8483
rect 58449 8449 58483 8483
rect 58483 8449 58492 8483
rect 58440 8440 58492 8449
rect 54116 8372 54168 8424
rect 60372 8415 60424 8424
rect 60372 8381 60381 8415
rect 60381 8381 60415 8415
rect 60415 8381 60424 8415
rect 60372 8372 60424 8381
rect 60924 8440 60976 8492
rect 61384 8483 61436 8492
rect 61384 8449 61393 8483
rect 61393 8449 61427 8483
rect 61427 8449 61436 8483
rect 61384 8440 61436 8449
rect 62120 8483 62172 8492
rect 62120 8449 62129 8483
rect 62129 8449 62163 8483
rect 62163 8449 62172 8483
rect 62120 8440 62172 8449
rect 63592 8483 63644 8492
rect 63592 8449 63601 8483
rect 63601 8449 63635 8483
rect 63635 8449 63644 8483
rect 63592 8440 63644 8449
rect 64420 8483 64472 8492
rect 64420 8449 64429 8483
rect 64429 8449 64463 8483
rect 64463 8449 64472 8483
rect 64420 8440 64472 8449
rect 65248 8483 65300 8492
rect 65248 8449 65257 8483
rect 65257 8449 65291 8483
rect 65291 8449 65300 8483
rect 65248 8440 65300 8449
rect 66812 8483 66864 8492
rect 66812 8449 66821 8483
rect 66821 8449 66855 8483
rect 66855 8449 66864 8483
rect 66812 8440 66864 8449
rect 71320 8483 71372 8492
rect 71320 8449 71329 8483
rect 71329 8449 71363 8483
rect 71363 8449 71372 8483
rect 71320 8440 71372 8449
rect 74264 8483 74316 8492
rect 74264 8449 74273 8483
rect 74273 8449 74307 8483
rect 74307 8449 74316 8483
rect 74264 8440 74316 8449
rect 76472 8483 76524 8492
rect 76472 8449 76481 8483
rect 76481 8449 76515 8483
rect 76515 8449 76524 8483
rect 76472 8440 76524 8449
rect 76748 8483 76800 8492
rect 76748 8449 76757 8483
rect 76757 8449 76791 8483
rect 76791 8449 76800 8483
rect 76748 8440 76800 8449
rect 79416 8483 79468 8492
rect 79416 8449 79425 8483
rect 79425 8449 79459 8483
rect 79459 8449 79468 8483
rect 79416 8440 79468 8449
rect 81624 8483 81676 8492
rect 81624 8449 81633 8483
rect 81633 8449 81667 8483
rect 81667 8449 81676 8483
rect 81624 8440 81676 8449
rect 88800 8483 88852 8492
rect 88800 8449 88809 8483
rect 88809 8449 88843 8483
rect 88843 8449 88852 8483
rect 88800 8440 88852 8449
rect 89168 8440 89220 8492
rect 90916 8483 90968 8492
rect 90916 8449 90925 8483
rect 90925 8449 90959 8483
rect 90959 8449 90968 8483
rect 90916 8440 90968 8449
rect 91652 8483 91704 8492
rect 91652 8449 91661 8483
rect 91661 8449 91695 8483
rect 91695 8449 91704 8483
rect 91652 8440 91704 8449
rect 92388 8483 92440 8492
rect 92388 8449 92397 8483
rect 92397 8449 92431 8483
rect 92431 8449 92440 8483
rect 92388 8440 92440 8449
rect 93216 8483 93268 8492
rect 93216 8449 93225 8483
rect 93225 8449 93259 8483
rect 93259 8449 93268 8483
rect 93216 8440 93268 8449
rect 93492 8440 93544 8492
rect 94412 8483 94464 8492
rect 94412 8449 94421 8483
rect 94421 8449 94455 8483
rect 94455 8449 94464 8483
rect 94412 8440 94464 8449
rect 95148 8483 95200 8492
rect 95148 8449 95157 8483
rect 95157 8449 95191 8483
rect 95191 8449 95200 8483
rect 95148 8440 95200 8449
rect 95976 8440 96028 8492
rect 96436 8483 96488 8492
rect 96436 8449 96445 8483
rect 96445 8449 96479 8483
rect 96479 8449 96488 8483
rect 96436 8440 96488 8449
rect 96620 8483 96672 8492
rect 96620 8449 96629 8483
rect 96629 8449 96663 8483
rect 96663 8449 96672 8483
rect 96620 8440 96672 8449
rect 97264 8483 97316 8492
rect 97264 8449 97273 8483
rect 97273 8449 97307 8483
rect 97307 8449 97316 8483
rect 97264 8440 97316 8449
rect 98460 8483 98512 8492
rect 98460 8449 98469 8483
rect 98469 8449 98503 8483
rect 98503 8449 98512 8483
rect 98460 8440 98512 8449
rect 99932 8483 99984 8492
rect 99932 8449 99941 8483
rect 99941 8449 99975 8483
rect 99975 8449 99984 8483
rect 99932 8440 99984 8449
rect 100024 8483 100076 8492
rect 100024 8449 100033 8483
rect 100033 8449 100067 8483
rect 100067 8449 100076 8483
rect 100024 8440 100076 8449
rect 100668 8483 100720 8492
rect 100668 8449 100677 8483
rect 100677 8449 100711 8483
rect 100711 8449 100720 8483
rect 100668 8440 100720 8449
rect 111708 8440 111760 8492
rect 121276 8483 121328 8492
rect 121276 8449 121285 8483
rect 121285 8449 121319 8483
rect 121319 8449 121328 8483
rect 121276 8440 121328 8449
rect 121736 8483 121788 8492
rect 121736 8449 121745 8483
rect 121745 8449 121779 8483
rect 121779 8449 121788 8483
rect 121736 8440 121788 8449
rect 123024 8483 123076 8492
rect 123024 8449 123033 8483
rect 123033 8449 123067 8483
rect 123067 8449 123076 8483
rect 123024 8440 123076 8449
rect 123760 8483 123812 8492
rect 123760 8449 123769 8483
rect 123769 8449 123803 8483
rect 123803 8449 123812 8483
rect 123760 8440 123812 8449
rect 125416 8483 125468 8492
rect 125416 8449 125425 8483
rect 125425 8449 125459 8483
rect 125459 8449 125468 8483
rect 125416 8440 125468 8449
rect 126152 8483 126204 8492
rect 126152 8449 126161 8483
rect 126161 8449 126195 8483
rect 126195 8449 126204 8483
rect 126152 8440 126204 8449
rect 126888 8483 126940 8492
rect 126888 8449 126897 8483
rect 126897 8449 126931 8483
rect 126931 8449 126940 8483
rect 126888 8440 126940 8449
rect 127624 8483 127676 8492
rect 127624 8449 127633 8483
rect 127633 8449 127667 8483
rect 127667 8449 127676 8483
rect 127624 8440 127676 8449
rect 127808 8483 127860 8492
rect 127808 8449 127817 8483
rect 127817 8449 127851 8483
rect 127851 8449 127860 8483
rect 127808 8440 127860 8449
rect 3424 8236 3476 8288
rect 26884 8236 26936 8288
rect 26976 8236 27028 8288
rect 27620 8236 27672 8288
rect 65432 8347 65484 8356
rect 65432 8313 65441 8347
rect 65441 8313 65475 8347
rect 65475 8313 65484 8347
rect 65432 8304 65484 8313
rect 71596 8415 71648 8424
rect 71596 8381 71605 8415
rect 71605 8381 71639 8415
rect 71639 8381 71648 8415
rect 71596 8372 71648 8381
rect 74540 8415 74592 8424
rect 74540 8381 74549 8415
rect 74549 8381 74583 8415
rect 74583 8381 74592 8415
rect 74540 8372 74592 8381
rect 66904 8304 66956 8356
rect 51356 8236 51408 8288
rect 81900 8415 81952 8424
rect 81900 8381 81909 8415
rect 81909 8381 81943 8415
rect 81943 8381 81952 8415
rect 81900 8372 81952 8381
rect 88156 8372 88208 8424
rect 92940 8372 92992 8424
rect 84200 8236 84252 8288
rect 84844 8236 84896 8288
rect 90088 8279 90140 8288
rect 90088 8245 90097 8279
rect 90097 8245 90131 8279
rect 90131 8245 90140 8279
rect 90088 8236 90140 8245
rect 93124 8236 93176 8288
rect 94228 8304 94280 8356
rect 104164 8372 104216 8424
rect 114560 8372 114612 8424
rect 115848 8372 115900 8424
rect 125048 8372 125100 8424
rect 129096 8483 129148 8492
rect 129096 8449 129105 8483
rect 129105 8449 129139 8483
rect 129139 8449 129148 8483
rect 129096 8440 129148 8449
rect 129556 8440 129608 8492
rect 132132 8483 132184 8492
rect 132132 8449 132141 8483
rect 132141 8449 132175 8483
rect 132175 8449 132184 8483
rect 132132 8440 132184 8449
rect 132868 8440 132920 8492
rect 133144 8483 133196 8492
rect 133144 8449 133153 8483
rect 133153 8449 133187 8483
rect 133187 8449 133196 8483
rect 133144 8440 133196 8449
rect 134248 8483 134300 8492
rect 134248 8449 134257 8483
rect 134257 8449 134291 8483
rect 134291 8449 134300 8483
rect 134248 8440 134300 8449
rect 130568 8415 130620 8424
rect 96620 8304 96672 8356
rect 104900 8236 104952 8288
rect 105728 8236 105780 8288
rect 107936 8236 107988 8288
rect 130568 8381 130577 8415
rect 130577 8381 130611 8415
rect 130611 8381 130620 8415
rect 130568 8372 130620 8381
rect 129004 8304 129056 8356
rect 137376 8304 137428 8356
rect 160836 8508 160888 8560
rect 165160 8619 165212 8628
rect 165160 8585 165169 8619
rect 165169 8585 165203 8619
rect 165203 8585 165212 8619
rect 165160 8576 165212 8585
rect 169944 8619 169996 8628
rect 169944 8585 169953 8619
rect 169953 8585 169987 8619
rect 169987 8585 169996 8619
rect 169944 8576 169996 8585
rect 170036 8576 170088 8628
rect 185860 8576 185912 8628
rect 185952 8576 186004 8628
rect 187700 8508 187752 8560
rect 148692 8440 148744 8492
rect 156512 8415 156564 8424
rect 156512 8381 156521 8415
rect 156521 8381 156555 8415
rect 156555 8381 156564 8415
rect 156512 8372 156564 8381
rect 157616 8440 157668 8492
rect 157248 8372 157300 8424
rect 158720 8372 158772 8424
rect 159088 8372 159140 8424
rect 159824 8415 159876 8424
rect 159824 8381 159833 8415
rect 159833 8381 159867 8415
rect 159867 8381 159876 8415
rect 159824 8372 159876 8381
rect 161940 8440 161992 8492
rect 162676 8440 162728 8492
rect 163688 8483 163740 8492
rect 163688 8449 163697 8483
rect 163697 8449 163731 8483
rect 163731 8449 163740 8483
rect 163688 8440 163740 8449
rect 165528 8440 165580 8492
rect 167368 8440 167420 8492
rect 161572 8372 161624 8424
rect 159916 8304 159968 8356
rect 160928 8304 160980 8356
rect 161756 8372 161808 8424
rect 162216 8372 162268 8424
rect 162768 8372 162820 8424
rect 163964 8415 164016 8424
rect 163964 8381 163973 8415
rect 163973 8381 164007 8415
rect 164007 8381 164016 8415
rect 163964 8372 164016 8381
rect 164148 8372 164200 8424
rect 167092 8415 167144 8424
rect 167092 8381 167101 8415
rect 167101 8381 167135 8415
rect 167135 8381 167144 8415
rect 167092 8372 167144 8381
rect 167736 8372 167788 8424
rect 168104 8372 168156 8424
rect 169576 8415 169628 8424
rect 169576 8381 169585 8415
rect 169585 8381 169619 8415
rect 169619 8381 169628 8415
rect 169576 8372 169628 8381
rect 169760 8483 169812 8492
rect 169760 8449 169769 8483
rect 169769 8449 169803 8483
rect 169803 8449 169812 8483
rect 169760 8440 169812 8449
rect 173440 8440 173492 8492
rect 179972 8372 180024 8424
rect 183284 8483 183336 8492
rect 183284 8449 183293 8483
rect 183293 8449 183327 8483
rect 183327 8449 183336 8483
rect 183284 8440 183336 8449
rect 186964 8483 187016 8492
rect 186964 8449 186973 8483
rect 186973 8449 187007 8483
rect 187007 8449 187016 8483
rect 186964 8440 187016 8449
rect 187056 8440 187108 8492
rect 188436 8483 188488 8492
rect 188436 8449 188445 8483
rect 188445 8449 188479 8483
rect 188479 8449 188488 8483
rect 188436 8440 188488 8449
rect 189908 8576 189960 8628
rect 191288 8619 191340 8628
rect 191288 8585 191297 8619
rect 191297 8585 191331 8619
rect 191331 8585 191340 8619
rect 191288 8576 191340 8585
rect 191380 8576 191432 8628
rect 193588 8619 193640 8628
rect 193588 8585 193597 8619
rect 193597 8585 193631 8619
rect 193631 8585 193640 8619
rect 193588 8576 193640 8585
rect 194232 8619 194284 8628
rect 194232 8585 194241 8619
rect 194241 8585 194275 8619
rect 194275 8585 194284 8619
rect 194232 8576 194284 8585
rect 195612 8619 195664 8628
rect 195612 8585 195621 8619
rect 195621 8585 195655 8619
rect 195655 8585 195664 8619
rect 195612 8576 195664 8585
rect 196624 8619 196676 8628
rect 196624 8585 196633 8619
rect 196633 8585 196667 8619
rect 196667 8585 196676 8619
rect 196624 8576 196676 8585
rect 197544 8619 197596 8628
rect 197544 8585 197553 8619
rect 197553 8585 197587 8619
rect 197587 8585 197596 8619
rect 197544 8576 197596 8585
rect 198096 8576 198148 8628
rect 198832 8619 198884 8628
rect 198832 8585 198841 8619
rect 198841 8585 198875 8619
rect 198875 8585 198884 8619
rect 198832 8576 198884 8585
rect 199476 8619 199528 8628
rect 199476 8585 199485 8619
rect 199485 8585 199519 8619
rect 199519 8585 199528 8619
rect 199476 8576 199528 8585
rect 200856 8619 200908 8628
rect 200856 8585 200865 8619
rect 200865 8585 200899 8619
rect 200899 8585 200908 8619
rect 200856 8576 200908 8585
rect 200948 8576 201000 8628
rect 202696 8619 202748 8628
rect 202696 8585 202705 8619
rect 202705 8585 202739 8619
rect 202739 8585 202748 8619
rect 202696 8576 202748 8585
rect 203524 8619 203576 8628
rect 203524 8585 203533 8619
rect 203533 8585 203567 8619
rect 203567 8585 203576 8619
rect 203524 8576 203576 8585
rect 196532 8508 196584 8560
rect 190368 8483 190420 8492
rect 190368 8449 190377 8483
rect 190377 8449 190411 8483
rect 190411 8449 190420 8483
rect 190368 8440 190420 8449
rect 191932 8440 191984 8492
rect 192024 8483 192076 8492
rect 192024 8449 192033 8483
rect 192033 8449 192067 8483
rect 192067 8449 192076 8483
rect 192024 8440 192076 8449
rect 193220 8483 193272 8492
rect 193220 8449 193229 8483
rect 193229 8449 193263 8483
rect 193263 8449 193272 8483
rect 193220 8440 193272 8449
rect 193496 8440 193548 8492
rect 194048 8483 194100 8492
rect 194048 8449 194057 8483
rect 194057 8449 194091 8483
rect 194091 8449 194100 8483
rect 194048 8440 194100 8449
rect 196348 8440 196400 8492
rect 197360 8483 197412 8492
rect 197360 8449 197369 8483
rect 197369 8449 197403 8483
rect 197403 8449 197412 8483
rect 197360 8440 197412 8449
rect 199292 8483 199344 8492
rect 199292 8449 199301 8483
rect 199301 8449 199335 8483
rect 199335 8449 199344 8483
rect 199292 8440 199344 8449
rect 201040 8440 201092 8492
rect 202420 8440 202472 8492
rect 202512 8483 202564 8492
rect 202512 8449 202521 8483
rect 202521 8449 202555 8483
rect 202555 8449 202564 8483
rect 202512 8440 202564 8449
rect 196532 8372 196584 8424
rect 196716 8372 196768 8424
rect 197268 8372 197320 8424
rect 198096 8372 198148 8424
rect 198832 8372 198884 8424
rect 202236 8372 202288 8424
rect 202788 8372 202840 8424
rect 203156 8415 203208 8424
rect 203156 8381 203165 8415
rect 203165 8381 203199 8415
rect 203199 8381 203208 8415
rect 203156 8372 203208 8381
rect 161940 8304 161992 8356
rect 132868 8236 132920 8288
rect 146852 8236 146904 8288
rect 151728 8236 151780 8288
rect 160100 8236 160152 8288
rect 162400 8236 162452 8288
rect 162860 8304 162912 8356
rect 170036 8304 170088 8356
rect 196348 8304 196400 8356
rect 163320 8236 163372 8288
rect 201132 8304 201184 8356
rect 225880 8576 225932 8628
rect 225972 8619 226024 8628
rect 225972 8585 225981 8619
rect 225981 8585 226015 8619
rect 226015 8585 226024 8619
rect 225972 8576 226024 8585
rect 226708 8619 226760 8628
rect 226708 8585 226717 8619
rect 226717 8585 226751 8619
rect 226751 8585 226760 8619
rect 226708 8576 226760 8585
rect 228272 8619 228324 8628
rect 228272 8585 228281 8619
rect 228281 8585 228315 8619
rect 228315 8585 228324 8619
rect 228272 8576 228324 8585
rect 229100 8619 229152 8628
rect 229100 8585 229109 8619
rect 229109 8585 229143 8619
rect 229143 8585 229152 8619
rect 229100 8576 229152 8585
rect 231032 8619 231084 8628
rect 231032 8585 231041 8619
rect 231041 8585 231075 8619
rect 231075 8585 231084 8619
rect 231032 8576 231084 8585
rect 231952 8619 232004 8628
rect 231952 8585 231961 8619
rect 231961 8585 231995 8619
rect 231995 8585 232004 8619
rect 231952 8576 232004 8585
rect 232872 8576 232924 8628
rect 234896 8619 234948 8628
rect 234896 8585 234905 8619
rect 234905 8585 234939 8619
rect 234939 8585 234948 8619
rect 234896 8576 234948 8585
rect 236092 8576 236144 8628
rect 236644 8619 236696 8628
rect 236644 8585 236653 8619
rect 236653 8585 236687 8619
rect 236687 8585 236696 8619
rect 236644 8576 236696 8585
rect 242992 8576 243044 8628
rect 247776 8576 247828 8628
rect 258264 8619 258316 8628
rect 258264 8585 258273 8619
rect 258273 8585 258307 8619
rect 258307 8585 258316 8619
rect 258264 8576 258316 8585
rect 262588 8619 262640 8628
rect 223948 8508 224000 8560
rect 217968 8440 218020 8492
rect 220912 8440 220964 8492
rect 221832 8440 221884 8492
rect 223672 8440 223724 8492
rect 224776 8508 224828 8560
rect 224868 8508 224920 8560
rect 225788 8483 225840 8492
rect 225788 8449 225797 8483
rect 225797 8449 225831 8483
rect 225831 8449 225840 8483
rect 225788 8440 225840 8449
rect 226524 8483 226576 8492
rect 226524 8449 226533 8483
rect 226533 8449 226567 8483
rect 226567 8449 226576 8483
rect 226524 8440 226576 8449
rect 228088 8483 228140 8492
rect 228088 8449 228097 8483
rect 228097 8449 228131 8483
rect 228131 8449 228140 8483
rect 228088 8440 228140 8449
rect 228916 8483 228968 8492
rect 228916 8449 228925 8483
rect 228925 8449 228959 8483
rect 228959 8449 228968 8483
rect 228916 8440 228968 8449
rect 229468 8440 229520 8492
rect 229836 8508 229888 8560
rect 212356 8372 212408 8424
rect 211068 8236 211120 8288
rect 214564 8236 214616 8288
rect 223488 8372 223540 8424
rect 229560 8372 229612 8424
rect 229928 8440 229980 8492
rect 230112 8508 230164 8560
rect 262588 8585 262597 8619
rect 262597 8585 262631 8619
rect 262631 8585 262640 8619
rect 262588 8576 262640 8585
rect 263600 8576 263652 8628
rect 264244 8576 264296 8628
rect 264888 8576 264940 8628
rect 267464 8576 267516 8628
rect 267648 8576 267700 8628
rect 268292 8576 268344 8628
rect 270224 8576 270276 8628
rect 260932 8508 260984 8560
rect 266912 8508 266964 8560
rect 230664 8483 230716 8492
rect 230664 8449 230673 8483
rect 230673 8449 230707 8483
rect 230707 8449 230716 8483
rect 230664 8440 230716 8449
rect 230848 8483 230900 8492
rect 230848 8449 230857 8483
rect 230857 8449 230891 8483
rect 230891 8449 230900 8483
rect 230848 8440 230900 8449
rect 231768 8483 231820 8492
rect 231768 8449 231777 8483
rect 231777 8449 231811 8483
rect 231811 8449 231820 8483
rect 231768 8440 231820 8449
rect 233240 8483 233292 8492
rect 233240 8449 233249 8483
rect 233249 8449 233283 8483
rect 233283 8449 233292 8483
rect 233240 8440 233292 8449
rect 234528 8483 234580 8492
rect 234528 8449 234537 8483
rect 234537 8449 234571 8483
rect 234571 8449 234580 8483
rect 234528 8440 234580 8449
rect 229836 8415 229888 8424
rect 229836 8381 229845 8415
rect 229845 8381 229879 8415
rect 229879 8381 229888 8415
rect 229836 8372 229888 8381
rect 231032 8372 231084 8424
rect 235724 8483 235776 8492
rect 235724 8449 235733 8483
rect 235733 8449 235767 8483
rect 235767 8449 235776 8483
rect 235724 8440 235776 8449
rect 235908 8440 235960 8492
rect 236184 8440 236236 8492
rect 246396 8483 246448 8492
rect 246396 8449 246405 8483
rect 246405 8449 246439 8483
rect 246439 8449 246448 8483
rect 246396 8440 246448 8449
rect 246672 8483 246724 8492
rect 246672 8449 246681 8483
rect 246681 8449 246715 8483
rect 246715 8449 246724 8483
rect 246672 8440 246724 8449
rect 249340 8483 249392 8492
rect 249340 8449 249349 8483
rect 249349 8449 249383 8483
rect 249383 8449 249392 8483
rect 249340 8440 249392 8449
rect 251548 8483 251600 8492
rect 251548 8449 251557 8483
rect 251557 8449 251591 8483
rect 251591 8449 251600 8483
rect 251548 8440 251600 8449
rect 254492 8483 254544 8492
rect 254492 8449 254501 8483
rect 254501 8449 254535 8483
rect 254535 8449 254544 8483
rect 254492 8440 254544 8449
rect 256700 8483 256752 8492
rect 256700 8449 256709 8483
rect 256709 8449 256743 8483
rect 256743 8449 256752 8483
rect 256700 8440 256752 8449
rect 258080 8483 258132 8492
rect 258080 8449 258089 8483
rect 258089 8449 258123 8483
rect 258123 8449 258132 8483
rect 258080 8440 258132 8449
rect 258356 8440 258408 8492
rect 259184 8483 259236 8492
rect 259184 8449 259193 8483
rect 259193 8449 259227 8483
rect 259227 8449 259236 8483
rect 259184 8440 259236 8449
rect 236368 8372 236420 8424
rect 242900 8372 242952 8424
rect 249616 8415 249668 8424
rect 249616 8381 249625 8415
rect 249625 8381 249659 8415
rect 249659 8381 249668 8415
rect 249616 8372 249668 8381
rect 251824 8415 251876 8424
rect 251824 8381 251833 8415
rect 251833 8381 251867 8415
rect 251867 8381 251876 8415
rect 251824 8372 251876 8381
rect 254768 8415 254820 8424
rect 254768 8381 254777 8415
rect 254777 8381 254811 8415
rect 254811 8381 254820 8415
rect 254768 8372 254820 8381
rect 224776 8304 224828 8356
rect 226432 8304 226484 8356
rect 227076 8304 227128 8356
rect 230572 8304 230624 8356
rect 234528 8304 234580 8356
rect 234896 8304 234948 8356
rect 237932 8304 237984 8356
rect 238576 8304 238628 8356
rect 258908 8372 258960 8424
rect 259644 8372 259696 8424
rect 260196 8304 260248 8356
rect 261116 8440 261168 8492
rect 261484 8440 261536 8492
rect 263600 8440 263652 8492
rect 264244 8483 264296 8492
rect 264244 8449 264253 8483
rect 264253 8449 264287 8483
rect 264287 8449 264296 8483
rect 264244 8440 264296 8449
rect 264520 8440 264572 8492
rect 265164 8483 265216 8492
rect 265164 8449 265173 8483
rect 265173 8449 265207 8483
rect 265207 8449 265216 8483
rect 265164 8440 265216 8449
rect 265900 8440 265952 8492
rect 266452 8483 266504 8492
rect 266452 8449 266461 8483
rect 266461 8449 266495 8483
rect 266495 8449 266504 8483
rect 266452 8440 266504 8449
rect 267096 8440 267148 8492
rect 260840 8372 260892 8424
rect 265808 8372 265860 8424
rect 267648 8440 267700 8492
rect 267740 8483 267792 8492
rect 267740 8449 267749 8483
rect 267749 8449 267783 8483
rect 267783 8449 267792 8483
rect 267740 8440 267792 8449
rect 268016 8440 268068 8492
rect 268384 8440 268436 8492
rect 268568 8483 268620 8492
rect 268568 8449 268577 8483
rect 268577 8449 268611 8483
rect 268611 8449 268620 8483
rect 268568 8440 268620 8449
rect 268752 8440 268804 8492
rect 268108 8372 268160 8424
rect 269304 8415 269356 8424
rect 269304 8381 269313 8415
rect 269313 8381 269347 8415
rect 269347 8381 269356 8415
rect 269304 8372 269356 8381
rect 269488 8483 269540 8492
rect 269488 8449 269497 8483
rect 269497 8449 269531 8483
rect 269531 8449 269540 8483
rect 269488 8440 269540 8449
rect 270868 8440 270920 8492
rect 269672 8415 269724 8424
rect 269672 8381 269681 8415
rect 269681 8381 269715 8415
rect 269715 8381 269724 8415
rect 269672 8372 269724 8381
rect 270132 8415 270184 8424
rect 270132 8381 270141 8415
rect 270141 8381 270175 8415
rect 270175 8381 270184 8415
rect 270132 8372 270184 8381
rect 261208 8304 261260 8356
rect 261944 8304 261996 8356
rect 263968 8304 264020 8356
rect 268936 8304 268988 8356
rect 223580 8236 223632 8288
rect 228916 8236 228968 8288
rect 235816 8236 235868 8288
rect 236552 8236 236604 8288
rect 236920 8236 236972 8288
rect 243176 8236 243228 8288
rect 258816 8236 258868 8288
rect 260288 8236 260340 8288
rect 262680 8236 262732 8288
rect 264244 8236 264296 8288
rect 267464 8236 267516 8288
rect 268752 8236 268804 8288
rect 34748 8134 34800 8186
rect 34812 8134 34864 8186
rect 34876 8134 34928 8186
rect 34940 8134 34992 8186
rect 35004 8134 35056 8186
rect 102345 8134 102397 8186
rect 102409 8134 102461 8186
rect 102473 8134 102525 8186
rect 102537 8134 102589 8186
rect 102601 8134 102653 8186
rect 169942 8134 169994 8186
rect 170006 8134 170058 8186
rect 170070 8134 170122 8186
rect 170134 8134 170186 8186
rect 170198 8134 170250 8186
rect 237539 8134 237591 8186
rect 237603 8134 237655 8186
rect 237667 8134 237719 8186
rect 237731 8134 237783 8186
rect 237795 8134 237847 8186
rect 25228 8075 25280 8084
rect 25228 8041 25237 8075
rect 25237 8041 25271 8075
rect 25271 8041 25280 8075
rect 25228 8032 25280 8041
rect 28356 8075 28408 8084
rect 28356 8041 28365 8075
rect 28365 8041 28399 8075
rect 28399 8041 28408 8075
rect 28356 8032 28408 8041
rect 23204 7964 23256 8016
rect 47308 8032 47360 8084
rect 28540 7964 28592 8016
rect 48228 7964 48280 8016
rect 73712 7964 73764 8016
rect 82176 7964 82228 8016
rect 85580 7964 85632 8016
rect 118240 8032 118292 8084
rect 133052 8075 133104 8084
rect 133052 8041 133061 8075
rect 133061 8041 133095 8075
rect 133095 8041 133104 8075
rect 133052 8032 133104 8041
rect 160284 8075 160336 8084
rect 160284 8041 160293 8075
rect 160293 8041 160327 8075
rect 160327 8041 160336 8075
rect 160284 8032 160336 8041
rect 162308 8032 162360 8084
rect 166356 8075 166408 8084
rect 166356 8041 166365 8075
rect 166365 8041 166399 8075
rect 166399 8041 166408 8075
rect 166356 8032 166408 8041
rect 166816 8032 166868 8084
rect 167828 8075 167880 8084
rect 167828 8041 167837 8075
rect 167837 8041 167871 8075
rect 167871 8041 167880 8075
rect 167828 8032 167880 8041
rect 168380 8032 168432 8084
rect 208400 8032 208452 8084
rect 217968 8032 218020 8084
rect 225880 8032 225932 8084
rect 93308 8007 93360 8016
rect 93308 7973 93317 8007
rect 93317 7973 93351 8007
rect 93351 7973 93360 8007
rect 93308 7964 93360 7973
rect 99288 7964 99340 8016
rect 107936 8007 107988 8016
rect 107936 7973 107945 8007
rect 107945 7973 107979 8007
rect 107979 7973 107988 8007
rect 107936 7964 107988 7973
rect 114928 7964 114980 8016
rect 150900 7964 150952 8016
rect 152832 7964 152884 8016
rect 162860 7964 162912 8016
rect 162952 7964 163004 8016
rect 184572 7964 184624 8016
rect 221096 7964 221148 8016
rect 227628 8032 227680 8084
rect 230388 8032 230440 8084
rect 230848 8075 230900 8084
rect 230848 8041 230857 8075
rect 230857 8041 230891 8075
rect 230891 8041 230900 8075
rect 230848 8032 230900 8041
rect 243084 8032 243136 8084
rect 14740 7896 14792 7948
rect 45744 7896 45796 7948
rect 81900 7896 81952 7948
rect 94964 7896 95016 7948
rect 99932 7896 99984 7948
rect 105176 7939 105228 7948
rect 105176 7905 105185 7939
rect 105185 7905 105219 7939
rect 105219 7905 105228 7939
rect 105176 7896 105228 7905
rect 106096 7896 106148 7948
rect 107752 7896 107804 7948
rect 141700 7896 141752 7948
rect 152556 7896 152608 7948
rect 161388 7939 161440 7948
rect 161388 7905 161397 7939
rect 161397 7905 161431 7939
rect 161431 7905 161440 7939
rect 161388 7896 161440 7905
rect 161664 7896 161716 7948
rect 162676 7896 162728 7948
rect 25044 7871 25096 7880
rect 25044 7837 25053 7871
rect 25053 7837 25087 7871
rect 25087 7837 25096 7871
rect 25044 7828 25096 7837
rect 26608 7871 26660 7880
rect 26608 7837 26617 7871
rect 26617 7837 26651 7871
rect 26651 7837 26660 7871
rect 26608 7828 26660 7837
rect 26240 7760 26292 7812
rect 27344 7871 27396 7880
rect 27344 7837 27353 7871
rect 27353 7837 27387 7871
rect 27387 7837 27396 7871
rect 27344 7828 27396 7837
rect 27528 7871 27580 7880
rect 27528 7837 27537 7871
rect 27537 7837 27571 7871
rect 27571 7837 27580 7871
rect 27528 7828 27580 7837
rect 28172 7871 28224 7880
rect 28172 7837 28181 7871
rect 28181 7837 28215 7871
rect 28215 7837 28224 7871
rect 28172 7828 28224 7837
rect 28908 7871 28960 7880
rect 28908 7837 28917 7871
rect 28917 7837 28951 7871
rect 28951 7837 28960 7871
rect 28908 7828 28960 7837
rect 29092 7828 29144 7880
rect 52828 7828 52880 7880
rect 90088 7828 90140 7880
rect 93124 7871 93176 7880
rect 93124 7837 93133 7871
rect 93133 7837 93167 7871
rect 93167 7837 93176 7871
rect 93124 7828 93176 7837
rect 99380 7871 99432 7880
rect 99380 7837 99389 7871
rect 99389 7837 99423 7871
rect 99423 7837 99432 7871
rect 99380 7828 99432 7837
rect 26792 7760 26844 7812
rect 51724 7760 51776 7812
rect 69848 7760 69900 7812
rect 85672 7760 85724 7812
rect 25688 7692 25740 7744
rect 26516 7692 26568 7744
rect 27804 7692 27856 7744
rect 27896 7692 27948 7744
rect 89720 7735 89772 7744
rect 89720 7701 89729 7735
rect 89729 7701 89763 7735
rect 89763 7701 89772 7735
rect 89720 7692 89772 7701
rect 94320 7692 94372 7744
rect 104164 7735 104216 7744
rect 104164 7701 104173 7735
rect 104173 7701 104207 7735
rect 104207 7701 104216 7735
rect 105636 7828 105688 7880
rect 105728 7871 105780 7880
rect 105728 7837 105737 7871
rect 105737 7837 105771 7871
rect 105771 7837 105780 7871
rect 105728 7828 105780 7837
rect 104164 7692 104216 7701
rect 105636 7692 105688 7744
rect 106556 7760 106608 7812
rect 108396 7760 108448 7812
rect 109868 7828 109920 7880
rect 132868 7871 132920 7880
rect 132868 7837 132877 7871
rect 132877 7837 132911 7871
rect 132911 7837 132920 7871
rect 132868 7828 132920 7837
rect 138664 7828 138716 7880
rect 149060 7828 149112 7880
rect 149152 7828 149204 7880
rect 158628 7828 158680 7880
rect 160100 7871 160152 7880
rect 160100 7837 160109 7871
rect 160109 7837 160143 7871
rect 160143 7837 160152 7871
rect 160100 7828 160152 7837
rect 163780 7871 163832 7880
rect 163780 7837 163789 7871
rect 163789 7837 163823 7871
rect 163823 7837 163832 7871
rect 163780 7828 163832 7837
rect 164332 7828 164384 7880
rect 164608 7871 164660 7880
rect 164608 7837 164617 7871
rect 164617 7837 164651 7871
rect 164651 7837 164660 7871
rect 164608 7828 164660 7837
rect 165620 7896 165672 7948
rect 165344 7871 165396 7880
rect 165344 7837 165353 7871
rect 165353 7837 165387 7871
rect 165387 7837 165396 7871
rect 165344 7828 165396 7837
rect 165436 7828 165488 7880
rect 166172 7871 166224 7880
rect 166172 7837 166181 7871
rect 166181 7837 166215 7871
rect 166215 7837 166224 7871
rect 166172 7828 166224 7837
rect 167460 7828 167512 7880
rect 167644 7871 167696 7880
rect 167644 7837 167653 7871
rect 167653 7837 167687 7871
rect 167687 7837 167696 7871
rect 167644 7828 167696 7837
rect 168840 7871 168892 7880
rect 168840 7837 168849 7871
rect 168849 7837 168883 7871
rect 168883 7837 168892 7871
rect 168840 7828 168892 7837
rect 169576 7939 169628 7948
rect 169576 7905 169585 7939
rect 169585 7905 169619 7939
rect 169619 7905 169628 7939
rect 169576 7896 169628 7905
rect 187240 7896 187292 7948
rect 203156 7896 203208 7948
rect 216312 7939 216364 7948
rect 216312 7905 216321 7939
rect 216321 7905 216355 7939
rect 216355 7905 216364 7939
rect 216312 7896 216364 7905
rect 218704 7896 218756 7948
rect 223396 7896 223448 7948
rect 236736 7964 236788 8016
rect 237196 7964 237248 8016
rect 239036 7964 239088 8016
rect 242900 7964 242952 8016
rect 254032 7896 254084 7948
rect 258356 8007 258408 8016
rect 258356 7973 258365 8007
rect 258365 7973 258399 8007
rect 258399 7973 258408 8007
rect 258356 7964 258408 7973
rect 258540 7896 258592 7948
rect 177212 7828 177264 7880
rect 212448 7828 212500 7880
rect 214656 7828 214708 7880
rect 106372 7735 106424 7744
rect 106372 7701 106381 7735
rect 106381 7701 106415 7735
rect 106415 7701 106424 7735
rect 106372 7692 106424 7701
rect 108764 7692 108816 7744
rect 141608 7760 141660 7812
rect 146484 7760 146536 7812
rect 146668 7760 146720 7812
rect 174728 7760 174780 7812
rect 189264 7760 189316 7812
rect 223580 7828 223632 7880
rect 217968 7760 218020 7812
rect 226064 7828 226116 7880
rect 230572 7828 230624 7880
rect 235724 7828 235776 7880
rect 237012 7871 237064 7880
rect 237012 7837 237021 7871
rect 237021 7837 237055 7871
rect 237055 7837 237064 7871
rect 237012 7828 237064 7837
rect 237380 7828 237432 7880
rect 237840 7871 237892 7880
rect 237840 7837 237849 7871
rect 237849 7837 237883 7871
rect 237883 7837 237892 7871
rect 237840 7828 237892 7837
rect 238024 7828 238076 7880
rect 239404 7828 239456 7880
rect 110512 7692 110564 7744
rect 111892 7692 111944 7744
rect 144000 7692 144052 7744
rect 146392 7692 146444 7744
rect 151452 7692 151504 7744
rect 160008 7692 160060 7744
rect 163872 7692 163924 7744
rect 164608 7692 164660 7744
rect 165344 7692 165396 7744
rect 214196 7692 214248 7744
rect 216404 7692 216456 7744
rect 216496 7692 216548 7744
rect 218336 7692 218388 7744
rect 218428 7692 218480 7744
rect 218980 7692 219032 7744
rect 219624 7692 219676 7744
rect 227628 7760 227680 7812
rect 231216 7760 231268 7812
rect 258172 7803 258224 7812
rect 258172 7769 258181 7803
rect 258181 7769 258215 7803
rect 258215 7769 258224 7803
rect 258172 7760 258224 7769
rect 228088 7692 228140 7744
rect 236092 7692 236144 7744
rect 236184 7692 236236 7744
rect 237656 7692 237708 7744
rect 242900 7692 242952 7744
rect 258816 7871 258868 7880
rect 258816 7837 258825 7871
rect 258825 7837 258859 7871
rect 258859 7837 258868 7871
rect 258816 7828 258868 7837
rect 259000 8075 259052 8084
rect 259000 8041 259009 8075
rect 259009 8041 259043 8075
rect 259043 8041 259052 8075
rect 259000 8032 259052 8041
rect 259828 8032 259880 8084
rect 260472 8075 260524 8084
rect 260472 8041 260481 8075
rect 260481 8041 260515 8075
rect 260515 8041 260524 8075
rect 260472 8032 260524 8041
rect 268016 8032 268068 8084
rect 268108 8032 268160 8084
rect 259920 7896 259972 7948
rect 264244 7896 264296 7948
rect 260288 7871 260340 7880
rect 260288 7837 260297 7871
rect 260297 7837 260331 7871
rect 260331 7837 260340 7871
rect 260288 7828 260340 7837
rect 261852 7871 261904 7880
rect 261852 7837 261861 7871
rect 261861 7837 261895 7871
rect 261895 7837 261904 7871
rect 261852 7828 261904 7837
rect 261944 7871 261996 7880
rect 261944 7837 261953 7871
rect 261953 7837 261987 7871
rect 261987 7837 261996 7871
rect 261944 7828 261996 7837
rect 262588 7871 262640 7880
rect 262588 7837 262597 7871
rect 262597 7837 262631 7871
rect 262631 7837 262640 7871
rect 262588 7828 262640 7837
rect 260840 7760 260892 7812
rect 263140 7828 263192 7880
rect 263784 7828 263836 7880
rect 260932 7692 260984 7744
rect 262312 7692 262364 7744
rect 263048 7692 263100 7744
rect 264152 7692 264204 7744
rect 264244 7735 264296 7744
rect 264244 7701 264253 7735
rect 264253 7701 264287 7735
rect 264287 7701 264296 7735
rect 264244 7692 264296 7701
rect 265256 7828 265308 7880
rect 265808 7871 265860 7880
rect 265808 7837 265817 7871
rect 265817 7837 265851 7871
rect 265851 7837 265860 7871
rect 265808 7828 265860 7837
rect 265992 7828 266044 7880
rect 267464 7828 267516 7880
rect 266176 7760 266228 7812
rect 267280 7803 267332 7812
rect 267280 7769 267289 7803
rect 267289 7769 267323 7803
rect 267323 7769 267332 7803
rect 267280 7760 267332 7769
rect 267648 7803 267700 7812
rect 267648 7769 267657 7803
rect 267657 7769 267691 7803
rect 267691 7769 267700 7803
rect 267648 7760 267700 7769
rect 268292 7871 268344 7880
rect 268292 7837 268301 7871
rect 268301 7837 268335 7871
rect 268335 7837 268344 7871
rect 268292 7828 268344 7837
rect 268568 7760 268620 7812
rect 265072 7692 265124 7744
rect 265440 7692 265492 7744
rect 266084 7735 266136 7744
rect 266084 7701 266093 7735
rect 266093 7701 266127 7735
rect 266127 7701 266136 7735
rect 266084 7692 266136 7701
rect 267464 7692 267516 7744
rect 269028 7896 269080 7948
rect 271788 7896 271840 7948
rect 268752 7760 268804 7812
rect 68546 7590 68598 7642
rect 68610 7590 68662 7642
rect 68674 7590 68726 7642
rect 68738 7590 68790 7642
rect 68802 7590 68854 7642
rect 136143 7590 136195 7642
rect 136207 7590 136259 7642
rect 136271 7590 136323 7642
rect 136335 7590 136387 7642
rect 136399 7590 136451 7642
rect 203740 7590 203792 7642
rect 203804 7590 203856 7642
rect 203868 7590 203920 7642
rect 203932 7590 203984 7642
rect 203996 7590 204048 7642
rect 271337 7590 271389 7642
rect 271401 7590 271453 7642
rect 271465 7590 271517 7642
rect 271529 7590 271581 7642
rect 271593 7590 271645 7642
rect 25136 7488 25188 7540
rect 26424 7531 26476 7540
rect 26424 7497 26433 7531
rect 26433 7497 26467 7531
rect 26467 7497 26476 7531
rect 26424 7488 26476 7497
rect 26608 7488 26660 7540
rect 20352 7420 20404 7472
rect 26792 7420 26844 7472
rect 31852 7488 31904 7540
rect 41972 7488 42024 7540
rect 66904 7488 66956 7540
rect 78220 7488 78272 7540
rect 104164 7488 104216 7540
rect 59820 7420 59872 7472
rect 60372 7420 60424 7472
rect 77576 7420 77628 7472
rect 94320 7420 94372 7472
rect 94412 7420 94464 7472
rect 24492 7395 24544 7404
rect 24492 7361 24501 7395
rect 24501 7361 24535 7395
rect 24535 7361 24544 7395
rect 24492 7352 24544 7361
rect 25044 7352 25096 7404
rect 26240 7395 26292 7404
rect 26240 7361 26249 7395
rect 26249 7361 26283 7395
rect 26283 7361 26292 7395
rect 26240 7352 26292 7361
rect 27804 7395 27856 7404
rect 27804 7361 27813 7395
rect 27813 7361 27847 7395
rect 27847 7361 27856 7395
rect 27804 7352 27856 7361
rect 25228 7327 25280 7336
rect 25228 7293 25237 7327
rect 25237 7293 25271 7327
rect 25271 7293 25280 7327
rect 25228 7284 25280 7293
rect 26056 7327 26108 7336
rect 26056 7293 26065 7327
rect 26065 7293 26099 7327
rect 26099 7293 26108 7327
rect 26056 7284 26108 7293
rect 23388 7216 23440 7268
rect 28540 7216 28592 7268
rect 37004 7216 37056 7268
rect 79416 7352 79468 7404
rect 80152 7284 80204 7336
rect 100208 7395 100260 7404
rect 100208 7361 100217 7395
rect 100217 7361 100251 7395
rect 100251 7361 100260 7395
rect 100208 7352 100260 7361
rect 107384 7395 107436 7404
rect 107384 7361 107393 7395
rect 107393 7361 107427 7395
rect 107427 7361 107436 7395
rect 107384 7352 107436 7361
rect 108396 7395 108448 7404
rect 108396 7361 108405 7395
rect 108405 7361 108439 7395
rect 108439 7361 108448 7395
rect 108396 7352 108448 7361
rect 121460 7488 121512 7540
rect 106832 7284 106884 7336
rect 107568 7284 107620 7336
rect 107844 7284 107896 7336
rect 110512 7395 110564 7404
rect 110512 7361 110521 7395
rect 110521 7361 110555 7395
rect 110555 7361 110564 7395
rect 110512 7352 110564 7361
rect 112076 7395 112128 7404
rect 112076 7361 112085 7395
rect 112085 7361 112119 7395
rect 112119 7361 112128 7395
rect 112076 7352 112128 7361
rect 120264 7352 120316 7404
rect 146300 7488 146352 7540
rect 146760 7488 146812 7540
rect 155592 7488 155644 7540
rect 161296 7531 161348 7540
rect 161296 7497 161305 7531
rect 161305 7497 161339 7531
rect 161339 7497 161348 7531
rect 161296 7488 161348 7497
rect 162584 7531 162636 7540
rect 162584 7497 162593 7531
rect 162593 7497 162627 7531
rect 162627 7497 162636 7531
rect 162584 7488 162636 7497
rect 162676 7488 162728 7540
rect 164056 7531 164108 7540
rect 164056 7497 164065 7531
rect 164065 7497 164099 7531
rect 164099 7497 164108 7531
rect 164056 7488 164108 7497
rect 164792 7531 164844 7540
rect 164792 7497 164801 7531
rect 164801 7497 164835 7531
rect 164835 7497 164844 7531
rect 164792 7488 164844 7497
rect 165528 7531 165580 7540
rect 165528 7497 165537 7531
rect 165537 7497 165571 7531
rect 165571 7497 165580 7531
rect 165528 7488 165580 7497
rect 168288 7488 168340 7540
rect 218704 7488 218756 7540
rect 221464 7488 221516 7540
rect 236920 7488 236972 7540
rect 237196 7488 237248 7540
rect 238944 7488 238996 7540
rect 259920 7488 259972 7540
rect 260380 7488 260432 7540
rect 261760 7531 261812 7540
rect 261760 7497 261769 7531
rect 261769 7497 261803 7531
rect 261803 7497 261812 7531
rect 261760 7488 261812 7497
rect 262496 7531 262548 7540
rect 262496 7497 262505 7531
rect 262505 7497 262539 7531
rect 262539 7497 262548 7531
rect 262496 7488 262548 7497
rect 263232 7531 263284 7540
rect 263232 7497 263241 7531
rect 263241 7497 263275 7531
rect 263275 7497 263284 7531
rect 263232 7488 263284 7497
rect 264336 7531 264388 7540
rect 264336 7497 264345 7531
rect 264345 7497 264379 7531
rect 264379 7497 264388 7531
rect 264336 7488 264388 7497
rect 270684 7488 270736 7540
rect 146760 7352 146812 7404
rect 152372 7420 152424 7472
rect 152556 7420 152608 7472
rect 168196 7420 168248 7472
rect 217968 7420 218020 7472
rect 226984 7420 227036 7472
rect 251364 7420 251416 7472
rect 23480 7148 23532 7200
rect 26240 7148 26292 7200
rect 78864 7216 78916 7268
rect 94412 7216 94464 7268
rect 79600 7148 79652 7200
rect 80152 7148 80204 7200
rect 100024 7191 100076 7200
rect 100024 7157 100033 7191
rect 100033 7157 100067 7191
rect 100067 7157 100076 7191
rect 100024 7148 100076 7157
rect 105176 7216 105228 7268
rect 107108 7259 107160 7268
rect 107108 7225 107117 7259
rect 107117 7225 107151 7259
rect 107151 7225 107160 7259
rect 107108 7216 107160 7225
rect 109132 7216 109184 7268
rect 110236 7259 110288 7268
rect 110236 7225 110245 7259
rect 110245 7225 110279 7259
rect 110279 7225 110288 7259
rect 110236 7216 110288 7225
rect 108580 7191 108632 7200
rect 108580 7157 108589 7191
rect 108589 7157 108623 7191
rect 108623 7157 108632 7191
rect 108580 7148 108632 7157
rect 110972 7284 111024 7336
rect 112628 7327 112680 7336
rect 112628 7293 112637 7327
rect 112637 7293 112671 7327
rect 112671 7293 112680 7327
rect 112628 7284 112680 7293
rect 112444 7216 112496 7268
rect 146116 7216 146168 7268
rect 146300 7259 146352 7268
rect 146300 7225 146309 7259
rect 146309 7225 146343 7259
rect 146343 7225 146352 7259
rect 146300 7216 146352 7225
rect 113088 7148 113140 7200
rect 147036 7284 147088 7336
rect 150992 7284 151044 7336
rect 147496 7191 147548 7200
rect 147496 7157 147505 7191
rect 147505 7157 147539 7191
rect 147539 7157 147548 7191
rect 147496 7148 147548 7157
rect 150900 7191 150952 7200
rect 150900 7157 150909 7191
rect 150909 7157 150943 7191
rect 150943 7157 150952 7191
rect 161112 7395 161164 7404
rect 161112 7361 161121 7395
rect 161121 7361 161155 7395
rect 161155 7361 161164 7395
rect 161112 7352 161164 7361
rect 162400 7395 162452 7404
rect 162400 7361 162409 7395
rect 162409 7361 162443 7395
rect 162443 7361 162452 7395
rect 162400 7352 162452 7361
rect 158628 7284 158680 7336
rect 162952 7284 163004 7336
rect 163872 7395 163924 7404
rect 163872 7361 163881 7395
rect 163881 7361 163915 7395
rect 163915 7361 163924 7395
rect 163872 7352 163924 7361
rect 164608 7395 164660 7404
rect 164608 7361 164617 7395
rect 164617 7361 164651 7395
rect 164651 7361 164660 7395
rect 164608 7352 164660 7361
rect 165344 7395 165396 7404
rect 165344 7361 165353 7395
rect 165353 7361 165387 7395
rect 165387 7361 165396 7395
rect 165344 7352 165396 7361
rect 169760 7352 169812 7404
rect 165160 7284 165212 7336
rect 172520 7284 172572 7336
rect 214196 7284 214248 7336
rect 181168 7216 181220 7268
rect 213920 7216 213972 7268
rect 214472 7395 214524 7404
rect 214472 7361 214481 7395
rect 214481 7361 214515 7395
rect 214515 7361 214524 7395
rect 214472 7352 214524 7361
rect 215576 7352 215628 7404
rect 216404 7395 216456 7404
rect 216404 7361 216413 7395
rect 216413 7361 216447 7395
rect 216447 7361 216456 7395
rect 216404 7352 216456 7361
rect 216680 7352 216732 7404
rect 218704 7395 218756 7404
rect 218704 7361 218713 7395
rect 218713 7361 218747 7395
rect 218747 7361 218756 7395
rect 218704 7352 218756 7361
rect 218980 7395 219032 7404
rect 218980 7361 218989 7395
rect 218989 7361 219023 7395
rect 219023 7361 219032 7395
rect 218980 7352 219032 7361
rect 220360 7352 220412 7404
rect 221464 7395 221516 7404
rect 221464 7361 221473 7395
rect 221473 7361 221507 7395
rect 221507 7361 221516 7395
rect 221464 7352 221516 7361
rect 221556 7395 221608 7404
rect 221556 7361 221590 7395
rect 221590 7361 221608 7395
rect 221556 7352 221608 7361
rect 221740 7395 221792 7404
rect 221740 7361 221749 7395
rect 221749 7361 221783 7395
rect 221783 7361 221792 7395
rect 221740 7352 221792 7361
rect 222844 7352 222896 7404
rect 223856 7395 223908 7404
rect 223856 7361 223865 7395
rect 223865 7361 223899 7395
rect 223899 7361 223908 7395
rect 223856 7352 223908 7361
rect 230112 7352 230164 7404
rect 230296 7395 230348 7404
rect 230296 7361 230305 7395
rect 230305 7361 230339 7395
rect 230339 7361 230348 7395
rect 230296 7352 230348 7361
rect 231216 7395 231268 7404
rect 231216 7361 231225 7395
rect 231225 7361 231259 7395
rect 231259 7361 231268 7395
rect 231216 7352 231268 7361
rect 231308 7352 231360 7404
rect 235264 7352 235316 7404
rect 235356 7395 235408 7404
rect 235356 7361 235365 7395
rect 235365 7361 235399 7395
rect 235399 7361 235408 7395
rect 235356 7352 235408 7361
rect 236000 7352 236052 7404
rect 236184 7395 236236 7404
rect 236184 7361 236193 7395
rect 236193 7361 236227 7395
rect 236227 7361 236236 7395
rect 236184 7352 236236 7361
rect 237288 7395 237340 7404
rect 237288 7361 237297 7395
rect 237297 7361 237331 7395
rect 237331 7361 237340 7395
rect 237288 7352 237340 7361
rect 237380 7352 237432 7404
rect 238024 7352 238076 7404
rect 238668 7352 238720 7404
rect 268016 7420 268068 7472
rect 215024 7284 215076 7336
rect 215116 7327 215168 7336
rect 215116 7293 215125 7327
rect 215125 7293 215159 7327
rect 215159 7293 215168 7327
rect 215116 7284 215168 7293
rect 150900 7148 150952 7157
rect 156052 7148 156104 7200
rect 159272 7148 159324 7200
rect 165620 7148 165672 7200
rect 169116 7191 169168 7200
rect 169116 7157 169125 7191
rect 169125 7157 169159 7191
rect 169159 7157 169168 7191
rect 169116 7148 169168 7157
rect 206928 7148 206980 7200
rect 212356 7148 212408 7200
rect 214840 7216 214892 7268
rect 216588 7327 216640 7336
rect 216588 7293 216597 7327
rect 216597 7293 216631 7327
rect 216631 7293 216640 7327
rect 216588 7284 216640 7293
rect 216956 7284 217008 7336
rect 216404 7216 216456 7268
rect 220728 7327 220780 7336
rect 220728 7293 220737 7327
rect 220737 7293 220771 7327
rect 220771 7293 220780 7327
rect 220728 7284 220780 7293
rect 218428 7259 218480 7268
rect 218428 7225 218437 7259
rect 218437 7225 218471 7259
rect 218471 7225 218480 7259
rect 218428 7216 218480 7225
rect 219992 7259 220044 7268
rect 219992 7225 220001 7259
rect 220001 7225 220035 7259
rect 220035 7225 220044 7259
rect 219992 7216 220044 7225
rect 220544 7216 220596 7268
rect 223120 7327 223172 7336
rect 223120 7293 223129 7327
rect 223129 7293 223163 7327
rect 223163 7293 223172 7327
rect 223120 7284 223172 7293
rect 223948 7327 224000 7336
rect 223948 7293 223982 7327
rect 223982 7293 224000 7327
rect 223948 7284 224000 7293
rect 224132 7327 224184 7336
rect 224132 7293 224141 7327
rect 224141 7293 224175 7327
rect 224175 7293 224184 7327
rect 224132 7284 224184 7293
rect 224960 7284 225012 7336
rect 218060 7148 218112 7200
rect 219716 7148 219768 7200
rect 222384 7191 222436 7200
rect 222384 7157 222393 7191
rect 222393 7157 222427 7191
rect 222427 7157 222436 7191
rect 222384 7148 222436 7157
rect 223304 7216 223356 7268
rect 225512 7216 225564 7268
rect 236092 7284 236144 7336
rect 239128 7284 239180 7336
rect 256792 7284 256844 7336
rect 261576 7395 261628 7404
rect 261576 7361 261585 7395
rect 261585 7361 261619 7395
rect 261619 7361 261628 7395
rect 261576 7352 261628 7361
rect 262312 7395 262364 7404
rect 262312 7361 262321 7395
rect 262321 7361 262355 7395
rect 262355 7361 262364 7395
rect 262312 7352 262364 7361
rect 263048 7395 263100 7404
rect 263048 7361 263057 7395
rect 263057 7361 263091 7395
rect 263091 7361 263100 7395
rect 263048 7352 263100 7361
rect 264152 7395 264204 7404
rect 264152 7361 264161 7395
rect 264161 7361 264195 7395
rect 264195 7361 264204 7395
rect 264152 7352 264204 7361
rect 264244 7352 264296 7404
rect 265256 7352 265308 7404
rect 267372 7395 267424 7404
rect 267372 7361 267381 7395
rect 267381 7361 267415 7395
rect 267415 7361 267424 7395
rect 267372 7352 267424 7361
rect 267648 7352 267700 7404
rect 270040 7420 270092 7472
rect 268384 7395 268436 7404
rect 268384 7361 268393 7395
rect 268393 7361 268427 7395
rect 268427 7361 268436 7395
rect 268384 7352 268436 7361
rect 269488 7395 269540 7404
rect 269488 7361 269497 7395
rect 269497 7361 269531 7395
rect 269531 7361 269540 7395
rect 269488 7352 269540 7361
rect 270500 7352 270552 7404
rect 263876 7216 263928 7268
rect 265808 7284 265860 7336
rect 266636 7284 266688 7336
rect 267004 7284 267056 7336
rect 267280 7284 267332 7336
rect 268016 7284 268068 7336
rect 268200 7284 268252 7336
rect 267740 7216 267792 7268
rect 271144 7284 271196 7336
rect 271972 7284 272024 7336
rect 226984 7148 227036 7200
rect 230204 7148 230256 7200
rect 230296 7148 230348 7200
rect 235632 7191 235684 7200
rect 235632 7157 235641 7191
rect 235641 7157 235675 7191
rect 235675 7157 235684 7191
rect 235632 7148 235684 7157
rect 236000 7148 236052 7200
rect 237288 7148 237340 7200
rect 237380 7148 237432 7200
rect 238760 7191 238812 7200
rect 238760 7157 238769 7191
rect 238769 7157 238803 7191
rect 238803 7157 238812 7191
rect 238760 7148 238812 7157
rect 239128 7191 239180 7200
rect 239128 7157 239137 7191
rect 239137 7157 239171 7191
rect 239171 7157 239180 7191
rect 239128 7148 239180 7157
rect 262680 7148 262732 7200
rect 264888 7191 264940 7200
rect 264888 7157 264897 7191
rect 264897 7157 264931 7191
rect 264931 7157 264940 7191
rect 264888 7148 264940 7157
rect 267464 7148 267516 7200
rect 267648 7148 267700 7200
rect 269396 7148 269448 7200
rect 34748 7046 34800 7098
rect 34812 7046 34864 7098
rect 34876 7046 34928 7098
rect 34940 7046 34992 7098
rect 35004 7046 35056 7098
rect 102345 7046 102397 7098
rect 102409 7046 102461 7098
rect 102473 7046 102525 7098
rect 102537 7046 102589 7098
rect 102601 7046 102653 7098
rect 169942 7046 169994 7098
rect 170006 7046 170058 7098
rect 170070 7046 170122 7098
rect 170134 7046 170186 7098
rect 170198 7046 170250 7098
rect 237539 7046 237591 7098
rect 237603 7046 237655 7098
rect 237667 7046 237719 7098
rect 237731 7046 237783 7098
rect 237795 7046 237847 7098
rect 79048 6944 79100 6996
rect 79416 6987 79468 6996
rect 79416 6953 79425 6987
rect 79425 6953 79459 6987
rect 79459 6953 79468 6987
rect 79416 6944 79468 6953
rect 100944 6944 100996 6996
rect 150256 6944 150308 6996
rect 165160 6944 165212 6996
rect 169116 6944 169168 6996
rect 26976 6876 27028 6928
rect 99840 6876 99892 6928
rect 107108 6876 107160 6928
rect 107752 6876 107804 6928
rect 19984 6740 20036 6792
rect 26148 6808 26200 6860
rect 75828 6808 75880 6860
rect 79692 6808 79744 6860
rect 92848 6808 92900 6860
rect 99012 6808 99064 6860
rect 100300 6851 100352 6860
rect 100300 6817 100309 6851
rect 100309 6817 100343 6851
rect 100343 6817 100352 6851
rect 100300 6808 100352 6817
rect 104440 6808 104492 6860
rect 24216 6740 24268 6792
rect 26516 6783 26568 6792
rect 26516 6749 26525 6783
rect 26525 6749 26559 6783
rect 26559 6749 26568 6783
rect 26516 6740 26568 6749
rect 33048 6740 33100 6792
rect 43996 6740 44048 6792
rect 47860 6740 47912 6792
rect 87880 6740 87932 6792
rect 92480 6740 92532 6792
rect 24400 6672 24452 6724
rect 38568 6672 38620 6724
rect 42616 6672 42668 6724
rect 49884 6672 49936 6724
rect 79140 6672 79192 6724
rect 89628 6672 89680 6724
rect 100576 6783 100628 6792
rect 100576 6749 100585 6783
rect 100585 6749 100619 6783
rect 100619 6749 100628 6783
rect 100576 6740 100628 6749
rect 101312 6740 101364 6792
rect 108120 6783 108172 6792
rect 108120 6749 108129 6783
rect 108129 6749 108163 6783
rect 108163 6749 108172 6783
rect 108764 6851 108816 6860
rect 108764 6817 108773 6851
rect 108773 6817 108807 6851
rect 108807 6817 108816 6851
rect 108764 6808 108816 6817
rect 146300 6876 146352 6928
rect 112444 6851 112496 6860
rect 112444 6817 112453 6851
rect 112453 6817 112487 6851
rect 112487 6817 112496 6851
rect 112444 6808 112496 6817
rect 113180 6851 113232 6860
rect 113180 6817 113189 6851
rect 113189 6817 113223 6851
rect 113223 6817 113232 6851
rect 113180 6808 113232 6817
rect 114928 6851 114980 6860
rect 114928 6817 114937 6851
rect 114937 6817 114971 6851
rect 114971 6817 114980 6851
rect 114928 6808 114980 6817
rect 140504 6808 140556 6860
rect 141332 6851 141384 6860
rect 141332 6817 141341 6851
rect 141341 6817 141375 6851
rect 141375 6817 141384 6851
rect 141332 6808 141384 6817
rect 141608 6851 141660 6860
rect 141608 6817 141617 6851
rect 141617 6817 141651 6851
rect 141651 6817 141660 6851
rect 141608 6808 141660 6817
rect 141700 6851 141752 6860
rect 141700 6817 141734 6851
rect 141734 6817 141752 6851
rect 141700 6808 141752 6817
rect 145840 6851 145892 6860
rect 145840 6817 145849 6851
rect 145849 6817 145883 6851
rect 145883 6817 145892 6851
rect 145840 6808 145892 6817
rect 146392 6808 146444 6860
rect 159180 6876 159232 6928
rect 161848 6876 161900 6928
rect 169760 6919 169812 6928
rect 169760 6885 169769 6919
rect 169769 6885 169803 6919
rect 169803 6885 169812 6919
rect 169760 6876 169812 6885
rect 180064 6944 180116 6996
rect 180984 6876 181036 6928
rect 190000 6919 190052 6928
rect 190000 6885 190009 6919
rect 190009 6885 190043 6919
rect 190043 6885 190052 6919
rect 190000 6876 190052 6885
rect 147588 6808 147640 6860
rect 148232 6851 148284 6860
rect 148232 6817 148241 6851
rect 148241 6817 148275 6851
rect 148275 6817 148284 6851
rect 148232 6808 148284 6817
rect 148968 6808 149020 6860
rect 149152 6851 149204 6860
rect 149152 6817 149161 6851
rect 149161 6817 149195 6851
rect 149195 6817 149204 6851
rect 149152 6808 149204 6817
rect 150348 6808 150400 6860
rect 150532 6851 150584 6860
rect 150532 6817 150541 6851
rect 150541 6817 150575 6851
rect 150575 6817 150584 6851
rect 150532 6808 150584 6817
rect 150900 6808 150952 6860
rect 151452 6851 151504 6860
rect 151452 6817 151461 6851
rect 151461 6817 151495 6851
rect 151495 6817 151504 6851
rect 151452 6808 151504 6817
rect 152372 6851 152424 6860
rect 152372 6817 152381 6851
rect 152381 6817 152415 6851
rect 152415 6817 152424 6851
rect 152372 6808 152424 6817
rect 189080 6808 189132 6860
rect 208768 6808 208820 6860
rect 210792 6808 210844 6860
rect 213920 6808 213972 6860
rect 215116 6944 215168 6996
rect 215484 6944 215536 6996
rect 215944 6876 215996 6928
rect 216588 6876 216640 6928
rect 215116 6808 215168 6860
rect 218060 6808 218112 6860
rect 218336 6876 218388 6928
rect 220820 6944 220872 6996
rect 225236 6944 225288 6996
rect 226248 6944 226300 6996
rect 229192 6944 229244 6996
rect 220912 6876 220964 6928
rect 219348 6808 219400 6860
rect 108120 6740 108172 6749
rect 109040 6783 109092 6792
rect 109040 6749 109049 6783
rect 109049 6749 109083 6783
rect 109083 6749 109092 6783
rect 109040 6740 109092 6749
rect 109224 6740 109276 6792
rect 109316 6783 109368 6792
rect 109316 6749 109325 6783
rect 109325 6749 109359 6783
rect 109359 6749 109368 6783
rect 109316 6740 109368 6749
rect 140872 6783 140924 6792
rect 140872 6749 140881 6783
rect 140881 6749 140915 6783
rect 140915 6749 140924 6783
rect 140872 6740 140924 6749
rect 141884 6783 141936 6792
rect 141884 6749 141893 6783
rect 141893 6749 141927 6783
rect 141927 6749 141936 6783
rect 141884 6740 141936 6749
rect 146760 6783 146812 6792
rect 146760 6749 146769 6783
rect 146769 6749 146803 6783
rect 146803 6749 146812 6783
rect 146760 6740 146812 6749
rect 146944 6740 146996 6792
rect 147036 6783 147088 6792
rect 147036 6749 147045 6783
rect 147045 6749 147079 6783
rect 147079 6749 147088 6783
rect 147036 6740 147088 6749
rect 148324 6740 148376 6792
rect 149428 6783 149480 6792
rect 149428 6749 149437 6783
rect 149437 6749 149471 6783
rect 149471 6749 149480 6783
rect 149428 6740 149480 6749
rect 150624 6740 150676 6792
rect 151544 6783 151596 6792
rect 151544 6749 151578 6783
rect 151578 6749 151596 6783
rect 151544 6740 151596 6749
rect 151728 6783 151780 6792
rect 151728 6749 151737 6783
rect 151737 6749 151771 6783
rect 151771 6749 151780 6783
rect 151728 6740 151780 6749
rect 169208 6783 169260 6792
rect 169208 6749 169217 6783
rect 169217 6749 169251 6783
rect 169251 6749 169260 6783
rect 169208 6740 169260 6749
rect 172520 6740 172572 6792
rect 189356 6740 189408 6792
rect 209872 6740 209924 6792
rect 211160 6783 211212 6792
rect 211160 6749 211169 6783
rect 211169 6749 211203 6783
rect 211203 6749 211212 6783
rect 211160 6740 211212 6749
rect 211344 6740 211396 6792
rect 211436 6783 211488 6792
rect 211436 6749 211445 6783
rect 211445 6749 211479 6783
rect 211479 6749 211488 6783
rect 211436 6740 211488 6749
rect 19248 6604 19300 6656
rect 24768 6604 24820 6656
rect 26700 6647 26752 6656
rect 26700 6613 26709 6647
rect 26709 6613 26743 6647
rect 26743 6613 26752 6647
rect 26700 6604 26752 6613
rect 43904 6604 43956 6656
rect 79416 6604 79468 6656
rect 80060 6604 80112 6656
rect 99012 6647 99064 6656
rect 99012 6613 99021 6647
rect 99021 6613 99055 6647
rect 99055 6613 99064 6647
rect 99012 6604 99064 6613
rect 102784 6715 102836 6724
rect 102784 6681 102793 6715
rect 102793 6681 102827 6715
rect 102827 6681 102836 6715
rect 102784 6672 102836 6681
rect 103336 6672 103388 6724
rect 106740 6672 106792 6724
rect 101772 6604 101824 6656
rect 109040 6604 109092 6656
rect 109960 6647 110012 6656
rect 109960 6613 109969 6647
rect 109969 6613 110003 6647
rect 110003 6613 110012 6647
rect 109960 6604 110012 6613
rect 112628 6715 112680 6724
rect 112628 6681 112637 6715
rect 112637 6681 112671 6715
rect 112671 6681 112680 6715
rect 112628 6672 112680 6681
rect 114376 6672 114428 6724
rect 125600 6672 125652 6724
rect 113364 6604 113416 6656
rect 115756 6604 115808 6656
rect 123484 6604 123536 6656
rect 141700 6604 141752 6656
rect 143080 6604 143132 6656
rect 146852 6604 146904 6656
rect 147036 6604 147088 6656
rect 148232 6604 148284 6656
rect 149428 6604 149480 6656
rect 150072 6647 150124 6656
rect 150072 6613 150081 6647
rect 150081 6613 150115 6647
rect 150115 6613 150124 6647
rect 150072 6604 150124 6613
rect 155592 6672 155644 6724
rect 163504 6672 163556 6724
rect 151084 6604 151136 6656
rect 151728 6604 151780 6656
rect 152372 6604 152424 6656
rect 161112 6604 161164 6656
rect 162676 6604 162728 6656
rect 198832 6604 198884 6656
rect 212080 6647 212132 6656
rect 212080 6613 212089 6647
rect 212089 6613 212123 6647
rect 212123 6613 212132 6647
rect 212080 6604 212132 6613
rect 213000 6672 213052 6724
rect 217692 6740 217744 6792
rect 216312 6672 216364 6724
rect 214288 6604 214340 6656
rect 215576 6604 215628 6656
rect 217600 6672 217652 6724
rect 218888 6783 218940 6792
rect 218888 6749 218897 6783
rect 218897 6749 218931 6783
rect 218931 6749 218940 6783
rect 218888 6740 218940 6749
rect 219072 6740 219124 6792
rect 219900 6740 219952 6792
rect 220544 6808 220596 6860
rect 221096 6851 221148 6860
rect 221096 6817 221105 6851
rect 221105 6817 221139 6851
rect 221139 6817 221148 6851
rect 221096 6808 221148 6817
rect 221740 6808 221792 6860
rect 221924 6808 221976 6860
rect 222108 6808 222160 6860
rect 217692 6604 217744 6656
rect 217876 6604 217928 6656
rect 221280 6740 221332 6792
rect 222292 6740 222344 6792
rect 223304 6851 223356 6860
rect 223304 6817 223313 6851
rect 223313 6817 223347 6851
rect 223347 6817 223356 6851
rect 223304 6808 223356 6817
rect 224960 6876 225012 6928
rect 226340 6876 226392 6928
rect 230112 6987 230164 6996
rect 230112 6953 230121 6987
rect 230121 6953 230155 6987
rect 230155 6953 230164 6987
rect 230112 6944 230164 6953
rect 230480 6944 230532 6996
rect 236920 6944 236972 6996
rect 230848 6876 230900 6928
rect 235724 6876 235776 6928
rect 236552 6876 236604 6928
rect 262680 6919 262732 6928
rect 262680 6885 262689 6919
rect 262689 6885 262723 6919
rect 262723 6885 262732 6919
rect 262680 6876 262732 6885
rect 224868 6808 224920 6860
rect 225512 6851 225564 6860
rect 225512 6817 225521 6851
rect 225521 6817 225555 6851
rect 225555 6817 225564 6851
rect 225512 6808 225564 6817
rect 229560 6851 229612 6860
rect 229560 6817 229569 6851
rect 229569 6817 229603 6851
rect 229603 6817 229612 6851
rect 229560 6808 229612 6817
rect 222108 6672 222160 6724
rect 223764 6740 223816 6792
rect 223856 6783 223908 6792
rect 223856 6749 223865 6783
rect 223865 6749 223899 6783
rect 223899 6749 223908 6783
rect 223856 6740 223908 6749
rect 220912 6604 220964 6656
rect 222016 6647 222068 6656
rect 222016 6613 222025 6647
rect 222025 6613 222059 6647
rect 222059 6613 222068 6647
rect 222016 6604 222068 6613
rect 223672 6604 223724 6656
rect 224592 6604 224644 6656
rect 227628 6740 227680 6792
rect 230480 6740 230532 6792
rect 231124 6783 231176 6792
rect 231124 6749 231133 6783
rect 231133 6749 231167 6783
rect 231167 6749 231176 6783
rect 231124 6740 231176 6749
rect 237380 6808 237432 6860
rect 263692 6876 263744 6928
rect 265072 6944 265124 6996
rect 270960 6944 271012 6996
rect 266176 6876 266228 6928
rect 225972 6672 226024 6724
rect 229008 6672 229060 6724
rect 231768 6715 231820 6724
rect 231768 6681 231777 6715
rect 231777 6681 231811 6715
rect 231811 6681 231820 6715
rect 231768 6672 231820 6681
rect 237196 6783 237248 6792
rect 237196 6749 237205 6783
rect 237205 6749 237239 6783
rect 237239 6749 237248 6783
rect 237196 6740 237248 6749
rect 261024 6783 261076 6792
rect 261024 6749 261033 6783
rect 261033 6749 261067 6783
rect 261067 6749 261076 6783
rect 261024 6740 261076 6749
rect 262496 6740 262548 6792
rect 268016 6808 268068 6860
rect 263508 6740 263560 6792
rect 264060 6783 264112 6792
rect 264060 6749 264069 6783
rect 264069 6749 264103 6783
rect 264103 6749 264112 6783
rect 264060 6740 264112 6749
rect 264244 6740 264296 6792
rect 265532 6783 265584 6792
rect 265532 6749 265541 6783
rect 265541 6749 265575 6783
rect 265575 6749 265584 6783
rect 265532 6740 265584 6749
rect 267004 6740 267056 6792
rect 237472 6672 237524 6724
rect 262128 6672 262180 6724
rect 228180 6604 228232 6656
rect 230480 6604 230532 6656
rect 237380 6647 237432 6656
rect 237380 6613 237389 6647
rect 237389 6613 237423 6647
rect 237423 6613 237432 6647
rect 237380 6604 237432 6613
rect 239128 6604 239180 6656
rect 258632 6604 258684 6656
rect 260196 6647 260248 6656
rect 260196 6613 260205 6647
rect 260205 6613 260239 6647
rect 260239 6613 260248 6647
rect 260196 6604 260248 6613
rect 263416 6604 263468 6656
rect 264152 6604 264204 6656
rect 264428 6604 264480 6656
rect 264704 6604 264756 6656
rect 265716 6647 265768 6656
rect 265716 6613 265725 6647
rect 265725 6613 265759 6647
rect 265759 6613 265768 6647
rect 265716 6604 265768 6613
rect 265808 6604 265860 6656
rect 267832 6740 267884 6792
rect 269212 6783 269264 6792
rect 269212 6749 269221 6783
rect 269221 6749 269255 6783
rect 269255 6749 269264 6783
rect 269212 6740 269264 6749
rect 269488 6783 269540 6792
rect 269488 6749 269497 6783
rect 269497 6749 269531 6783
rect 269531 6749 269540 6783
rect 269488 6740 269540 6749
rect 270500 6783 270552 6792
rect 270500 6749 270509 6783
rect 270509 6749 270543 6783
rect 270543 6749 270552 6783
rect 270500 6740 270552 6749
rect 270408 6672 270460 6724
rect 68546 6502 68598 6554
rect 68610 6502 68662 6554
rect 68674 6502 68726 6554
rect 68738 6502 68790 6554
rect 68802 6502 68854 6554
rect 136143 6502 136195 6554
rect 136207 6502 136259 6554
rect 136271 6502 136323 6554
rect 136335 6502 136387 6554
rect 136399 6502 136451 6554
rect 203740 6502 203792 6554
rect 203804 6502 203856 6554
rect 203868 6502 203920 6554
rect 203932 6502 203984 6554
rect 203996 6502 204048 6554
rect 271337 6502 271389 6554
rect 271401 6502 271453 6554
rect 271465 6502 271517 6554
rect 271529 6502 271581 6554
rect 271593 6502 271645 6554
rect 15568 6400 15620 6452
rect 42616 6400 42668 6452
rect 13728 6332 13780 6384
rect 36544 6332 36596 6384
rect 9956 6264 10008 6316
rect 42984 6332 43036 6384
rect 43352 6332 43404 6384
rect 46020 6400 46072 6452
rect 72332 6400 72384 6452
rect 43168 6307 43220 6316
rect 43168 6273 43177 6307
rect 43177 6273 43211 6307
rect 43211 6273 43220 6307
rect 43168 6264 43220 6273
rect 43904 6375 43956 6384
rect 43904 6341 43913 6375
rect 43913 6341 43947 6375
rect 43947 6341 43956 6375
rect 43904 6332 43956 6341
rect 45008 6375 45060 6384
rect 45008 6341 45017 6375
rect 45017 6341 45051 6375
rect 45051 6341 45060 6375
rect 45008 6332 45060 6341
rect 45560 6332 45612 6384
rect 45744 6375 45796 6384
rect 45744 6341 45753 6375
rect 45753 6341 45787 6375
rect 45787 6341 45796 6375
rect 45744 6332 45796 6341
rect 79324 6332 79376 6384
rect 79600 6443 79652 6452
rect 79600 6409 79609 6443
rect 79609 6409 79643 6443
rect 79643 6409 79652 6443
rect 79600 6400 79652 6409
rect 99012 6400 99064 6452
rect 100116 6443 100168 6452
rect 100116 6409 100125 6443
rect 100125 6409 100159 6443
rect 100159 6409 100168 6443
rect 100116 6400 100168 6409
rect 100208 6400 100260 6452
rect 100760 6400 100812 6452
rect 104716 6400 104768 6452
rect 107292 6400 107344 6452
rect 108580 6400 108632 6452
rect 109316 6400 109368 6452
rect 111248 6400 111300 6452
rect 144460 6400 144512 6452
rect 148048 6400 148100 6452
rect 162492 6400 162544 6452
rect 162584 6400 162636 6452
rect 168288 6400 168340 6452
rect 181812 6443 181864 6452
rect 181812 6409 181821 6443
rect 181821 6409 181855 6443
rect 181855 6409 181864 6443
rect 181812 6400 181864 6409
rect 189172 6443 189224 6452
rect 81348 6332 81400 6384
rect 91468 6332 91520 6384
rect 45376 6307 45428 6316
rect 45376 6273 45385 6307
rect 45385 6273 45419 6307
rect 45419 6273 45428 6307
rect 45376 6264 45428 6273
rect 23664 6196 23716 6248
rect 40500 6196 40552 6248
rect 44732 6196 44784 6248
rect 46020 6196 46072 6248
rect 47584 6196 47636 6248
rect 71596 6196 71648 6248
rect 87696 6264 87748 6316
rect 100668 6332 100720 6384
rect 99932 6264 99984 6316
rect 108120 6332 108172 6384
rect 101772 6307 101824 6316
rect 101772 6273 101781 6307
rect 101781 6273 101815 6307
rect 101815 6273 101824 6307
rect 101772 6264 101824 6273
rect 106372 6264 106424 6316
rect 108672 6264 108724 6316
rect 17224 6128 17276 6180
rect 42524 6128 42576 6180
rect 44088 6171 44140 6180
rect 44088 6137 44097 6171
rect 44097 6137 44131 6171
rect 44131 6137 44140 6171
rect 44088 6128 44140 6137
rect 79048 6171 79100 6180
rect 79048 6137 79057 6171
rect 79057 6137 79091 6171
rect 79091 6137 79100 6171
rect 79048 6128 79100 6137
rect 79416 6103 79468 6112
rect 79416 6069 79425 6103
rect 79425 6069 79459 6103
rect 79459 6069 79468 6103
rect 79416 6060 79468 6069
rect 79692 6128 79744 6180
rect 92756 6196 92808 6248
rect 93400 6239 93452 6248
rect 93400 6205 93409 6239
rect 93409 6205 93443 6239
rect 93443 6205 93452 6239
rect 93400 6196 93452 6205
rect 99748 6171 99800 6180
rect 99748 6137 99757 6171
rect 99757 6137 99791 6171
rect 99791 6137 99800 6171
rect 99748 6128 99800 6137
rect 90272 6060 90324 6112
rect 96804 6060 96856 6112
rect 100116 6103 100168 6112
rect 100116 6069 100125 6103
rect 100125 6069 100159 6103
rect 100159 6069 100168 6103
rect 100116 6060 100168 6069
rect 102232 6239 102284 6248
rect 102232 6205 102241 6239
rect 102241 6205 102275 6239
rect 102275 6205 102284 6239
rect 102232 6196 102284 6205
rect 104716 6196 104768 6248
rect 112076 6332 112128 6384
rect 115940 6332 115992 6384
rect 109960 6264 110012 6316
rect 112720 6307 112772 6316
rect 112720 6273 112729 6307
rect 112729 6273 112763 6307
rect 112763 6273 112772 6307
rect 112720 6264 112772 6273
rect 119988 6332 120040 6384
rect 130200 6332 130252 6384
rect 130292 6375 130344 6384
rect 130292 6341 130301 6375
rect 130301 6341 130335 6375
rect 130335 6341 130344 6375
rect 130292 6332 130344 6341
rect 141332 6332 141384 6384
rect 143448 6332 143500 6384
rect 122104 6264 122156 6316
rect 109316 6196 109368 6248
rect 112628 6196 112680 6248
rect 119068 6196 119120 6248
rect 122012 6196 122064 6248
rect 125140 6307 125192 6316
rect 125140 6273 125149 6307
rect 125149 6273 125183 6307
rect 125183 6273 125192 6307
rect 125140 6264 125192 6273
rect 129924 6264 129976 6316
rect 147496 6332 147548 6384
rect 147680 6332 147732 6384
rect 148784 6332 148836 6384
rect 148968 6332 149020 6384
rect 150716 6332 150768 6384
rect 152648 6375 152700 6384
rect 152648 6341 152657 6375
rect 152657 6341 152691 6375
rect 152691 6341 152700 6375
rect 152648 6332 152700 6341
rect 152740 6332 152792 6384
rect 162860 6332 162912 6384
rect 114376 6128 114428 6180
rect 120264 6171 120316 6180
rect 120264 6137 120273 6171
rect 120273 6137 120307 6171
rect 120307 6137 120316 6171
rect 120264 6128 120316 6137
rect 103152 6060 103204 6112
rect 107660 6060 107712 6112
rect 108764 6060 108816 6112
rect 112076 6060 112128 6112
rect 115848 6060 115900 6112
rect 120080 6103 120132 6112
rect 120080 6069 120089 6103
rect 120089 6069 120123 6103
rect 120123 6069 120132 6103
rect 122104 6128 122156 6180
rect 122196 6128 122248 6180
rect 120080 6060 120132 6069
rect 122564 6060 122616 6112
rect 125600 6128 125652 6180
rect 142620 6128 142672 6180
rect 143356 6196 143408 6248
rect 148876 6307 148928 6316
rect 148876 6273 148885 6307
rect 148885 6273 148919 6307
rect 148919 6273 148928 6307
rect 148876 6264 148928 6273
rect 150072 6264 150124 6316
rect 156144 6264 156196 6316
rect 156788 6264 156840 6316
rect 156972 6264 157024 6316
rect 158168 6264 158220 6316
rect 177856 6332 177908 6384
rect 180984 6332 181036 6384
rect 189172 6409 189197 6443
rect 189197 6409 189224 6443
rect 189172 6400 189224 6409
rect 189356 6443 189408 6452
rect 189356 6409 189365 6443
rect 189365 6409 189399 6443
rect 189399 6409 189408 6443
rect 189356 6400 189408 6409
rect 182180 6332 182232 6384
rect 148140 6239 148192 6248
rect 148140 6205 148149 6239
rect 148149 6205 148183 6239
rect 148183 6205 148192 6239
rect 148140 6196 148192 6205
rect 148416 6196 148468 6248
rect 150992 6239 151044 6248
rect 150992 6205 151001 6239
rect 151001 6205 151035 6239
rect 151035 6205 151044 6239
rect 150992 6196 151044 6205
rect 153292 6196 153344 6248
rect 157064 6239 157116 6248
rect 157064 6205 157073 6239
rect 157073 6205 157107 6239
rect 157107 6205 157116 6239
rect 157064 6196 157116 6205
rect 157248 6196 157300 6248
rect 161572 6239 161624 6248
rect 161572 6205 161581 6239
rect 161581 6205 161615 6239
rect 161615 6205 161624 6239
rect 161572 6196 161624 6205
rect 162584 6196 162636 6248
rect 162860 6196 162912 6248
rect 182548 6307 182600 6316
rect 182548 6273 182557 6307
rect 182557 6273 182591 6307
rect 182591 6273 182600 6307
rect 182548 6264 182600 6273
rect 188436 6332 188488 6384
rect 216772 6400 216824 6452
rect 218336 6400 218388 6452
rect 219900 6400 219952 6452
rect 221188 6400 221240 6452
rect 169208 6128 169260 6180
rect 182088 6196 182140 6248
rect 200764 6264 200816 6316
rect 212080 6332 212132 6384
rect 217876 6332 217928 6384
rect 222108 6332 222160 6384
rect 223856 6332 223908 6384
rect 224132 6332 224184 6384
rect 225328 6332 225380 6384
rect 225604 6400 225656 6452
rect 254768 6400 254820 6452
rect 258632 6400 258684 6452
rect 262956 6400 263008 6452
rect 263416 6443 263468 6452
rect 263416 6409 263425 6443
rect 263425 6409 263459 6443
rect 263459 6409 263468 6443
rect 263416 6400 263468 6409
rect 263508 6400 263560 6452
rect 265624 6400 265676 6452
rect 266176 6400 266228 6452
rect 269212 6400 269264 6452
rect 226984 6332 227036 6384
rect 227720 6332 227772 6384
rect 244280 6332 244332 6384
rect 264704 6332 264756 6384
rect 217784 6307 217836 6316
rect 217784 6273 217793 6307
rect 217793 6273 217827 6307
rect 217827 6273 217836 6307
rect 217784 6264 217836 6273
rect 221188 6307 221240 6316
rect 221188 6273 221197 6307
rect 221197 6273 221231 6307
rect 221231 6273 221240 6307
rect 221188 6264 221240 6273
rect 221372 6264 221424 6316
rect 221464 6307 221516 6316
rect 221464 6273 221473 6307
rect 221473 6273 221507 6307
rect 221507 6273 221516 6307
rect 221464 6264 221516 6273
rect 223396 6307 223448 6316
rect 223396 6273 223405 6307
rect 223405 6273 223439 6307
rect 223439 6273 223448 6307
rect 223396 6264 223448 6273
rect 223672 6307 223724 6316
rect 223672 6273 223681 6307
rect 223681 6273 223715 6307
rect 223715 6273 223724 6307
rect 223672 6264 223724 6273
rect 207756 6239 207808 6248
rect 207756 6205 207765 6239
rect 207765 6205 207799 6239
rect 207799 6205 207808 6239
rect 207756 6196 207808 6205
rect 208400 6239 208452 6248
rect 208400 6205 208409 6239
rect 208409 6205 208443 6239
rect 208443 6205 208452 6239
rect 208400 6196 208452 6205
rect 214104 6196 214156 6248
rect 214656 6196 214708 6248
rect 215300 6196 215352 6248
rect 217140 6196 217192 6248
rect 217968 6239 218020 6248
rect 217968 6205 217977 6239
rect 217977 6205 218011 6239
rect 218011 6205 218020 6239
rect 217968 6196 218020 6205
rect 218336 6196 218388 6248
rect 218060 6128 218112 6180
rect 155040 6060 155092 6112
rect 156328 6103 156380 6112
rect 156328 6069 156337 6103
rect 156337 6069 156371 6103
rect 156371 6069 156380 6103
rect 156328 6060 156380 6069
rect 158812 6060 158864 6112
rect 169300 6060 169352 6112
rect 189080 6060 189132 6112
rect 206928 6060 206980 6112
rect 218796 6239 218848 6248
rect 218796 6205 218830 6239
rect 218830 6205 218848 6239
rect 218796 6196 218848 6205
rect 218980 6239 219032 6248
rect 218980 6205 218989 6239
rect 218989 6205 219023 6239
rect 219023 6205 219032 6239
rect 218980 6196 219032 6205
rect 219164 6196 219216 6248
rect 220360 6196 220412 6248
rect 220544 6196 220596 6248
rect 219900 6128 219952 6180
rect 219164 6060 219216 6112
rect 219440 6060 219492 6112
rect 220636 6060 220688 6112
rect 223856 6239 223908 6248
rect 223856 6205 223865 6239
rect 223865 6205 223899 6239
rect 223899 6205 223908 6239
rect 223856 6196 223908 6205
rect 224132 6196 224184 6248
rect 225880 6307 225932 6316
rect 225880 6273 225889 6307
rect 225889 6273 225923 6307
rect 225923 6273 225932 6307
rect 225880 6264 225932 6273
rect 226064 6264 226116 6316
rect 225328 6196 225380 6248
rect 226708 6196 226760 6248
rect 230296 6264 230348 6316
rect 235632 6264 235684 6316
rect 237380 6264 237432 6316
rect 261208 6307 261260 6316
rect 261208 6273 261217 6307
rect 261217 6273 261251 6307
rect 261251 6273 261260 6307
rect 261208 6264 261260 6273
rect 262404 6307 262456 6316
rect 262404 6273 262413 6307
rect 262413 6273 262447 6307
rect 262447 6273 262456 6307
rect 262404 6264 262456 6273
rect 262496 6307 262548 6316
rect 262496 6273 262505 6307
rect 262505 6273 262539 6307
rect 262539 6273 262548 6307
rect 262496 6264 262548 6273
rect 228456 6196 228508 6248
rect 231584 6196 231636 6248
rect 231676 6239 231728 6248
rect 231676 6205 231685 6239
rect 231685 6205 231719 6239
rect 231719 6205 231728 6239
rect 231676 6196 231728 6205
rect 231768 6196 231820 6248
rect 261484 6239 261536 6248
rect 261484 6205 261493 6239
rect 261493 6205 261527 6239
rect 261527 6205 261536 6239
rect 261484 6196 261536 6205
rect 224224 6128 224276 6180
rect 226248 6128 226300 6180
rect 226984 6128 227036 6180
rect 252836 6128 252888 6180
rect 260196 6128 260248 6180
rect 264244 6307 264296 6316
rect 264244 6273 264253 6307
rect 264253 6273 264287 6307
rect 264287 6273 264296 6307
rect 264244 6264 264296 6273
rect 264612 6307 264664 6316
rect 264612 6273 264621 6307
rect 264621 6273 264655 6307
rect 264655 6273 264664 6307
rect 264612 6264 264664 6273
rect 265808 6264 265860 6316
rect 267832 6307 267884 6316
rect 267832 6273 267841 6307
rect 267841 6273 267875 6307
rect 267875 6273 267884 6307
rect 267832 6264 267884 6273
rect 268476 6264 268528 6316
rect 269396 6307 269448 6316
rect 269396 6273 269405 6307
rect 269405 6273 269439 6307
rect 269439 6273 269448 6307
rect 269396 6264 269448 6273
rect 270408 6264 270460 6316
rect 265164 6196 265216 6248
rect 266912 6239 266964 6248
rect 266912 6205 266921 6239
rect 266921 6205 266955 6239
rect 266955 6205 266964 6239
rect 266912 6196 266964 6205
rect 269120 6196 269172 6248
rect 270040 6196 270092 6248
rect 226432 6060 226484 6112
rect 226524 6060 226576 6112
rect 227720 6060 227772 6112
rect 229836 6060 229888 6112
rect 230112 6060 230164 6112
rect 230480 6103 230532 6112
rect 230480 6069 230489 6103
rect 230489 6069 230523 6103
rect 230523 6069 230532 6103
rect 230480 6060 230532 6069
rect 230756 6060 230808 6112
rect 231124 6060 231176 6112
rect 238760 6060 238812 6112
rect 261668 6060 261720 6112
rect 268108 6128 268160 6180
rect 266728 6060 266780 6112
rect 267096 6060 267148 6112
rect 269028 6060 269080 6112
rect 270316 6060 270368 6112
rect 271972 6060 272024 6112
rect 34748 5958 34800 6010
rect 34812 5958 34864 6010
rect 34876 5958 34928 6010
rect 34940 5958 34992 6010
rect 35004 5958 35056 6010
rect 102345 5958 102397 6010
rect 102409 5958 102461 6010
rect 102473 5958 102525 6010
rect 102537 5958 102589 6010
rect 102601 5958 102653 6010
rect 169942 5958 169994 6010
rect 170006 5958 170058 6010
rect 170070 5958 170122 6010
rect 170134 5958 170186 6010
rect 170198 5958 170250 6010
rect 237539 5958 237591 6010
rect 237603 5958 237655 6010
rect 237667 5958 237719 6010
rect 237731 5958 237783 6010
rect 237795 5958 237847 6010
rect 36544 5856 36596 5908
rect 42800 5856 42852 5908
rect 47860 5899 47912 5908
rect 47860 5865 47869 5899
rect 47869 5865 47903 5899
rect 47903 5865 47912 5899
rect 47860 5856 47912 5865
rect 79048 5856 79100 5908
rect 99748 5856 99800 5908
rect 120080 5856 120132 5908
rect 77300 5788 77352 5840
rect 84200 5788 84252 5840
rect 33232 5720 33284 5772
rect 42708 5695 42760 5704
rect 11336 5584 11388 5636
rect 42708 5661 42717 5695
rect 42717 5661 42751 5695
rect 42751 5661 42760 5695
rect 42708 5652 42760 5661
rect 42064 5627 42116 5636
rect 42064 5593 42073 5627
rect 42073 5593 42107 5627
rect 42107 5593 42116 5627
rect 42064 5584 42116 5593
rect 44732 5720 44784 5772
rect 46020 5720 46072 5772
rect 47584 5720 47636 5772
rect 48044 5720 48096 5772
rect 51632 5720 51684 5772
rect 53104 5720 53156 5772
rect 79324 5720 79376 5772
rect 80796 5720 80848 5772
rect 81992 5763 82044 5772
rect 81992 5729 82001 5763
rect 82001 5729 82035 5763
rect 82035 5729 82044 5763
rect 81992 5720 82044 5729
rect 84936 5720 84988 5772
rect 93860 5788 93912 5840
rect 99932 5720 99984 5772
rect 100116 5788 100168 5840
rect 108856 5720 108908 5772
rect 109040 5763 109092 5772
rect 109040 5729 109049 5763
rect 109049 5729 109083 5763
rect 109083 5729 109092 5763
rect 109040 5720 109092 5729
rect 111248 5831 111300 5840
rect 111248 5797 111257 5831
rect 111257 5797 111291 5831
rect 111291 5797 111300 5831
rect 111248 5788 111300 5797
rect 111524 5831 111576 5840
rect 111524 5797 111533 5831
rect 111533 5797 111567 5831
rect 111567 5797 111576 5831
rect 111524 5788 111576 5797
rect 115112 5788 115164 5840
rect 115756 5788 115808 5840
rect 115848 5788 115900 5840
rect 119988 5720 120040 5772
rect 162768 5856 162820 5908
rect 163044 5856 163096 5908
rect 43444 5652 43496 5704
rect 43628 5695 43680 5704
rect 43628 5661 43637 5695
rect 43637 5661 43671 5695
rect 43671 5661 43680 5695
rect 43628 5652 43680 5661
rect 43720 5652 43772 5704
rect 44364 5695 44416 5704
rect 44364 5661 44387 5695
rect 44387 5661 44416 5695
rect 44364 5652 44416 5661
rect 46848 5695 46900 5704
rect 46848 5661 46857 5695
rect 46857 5661 46891 5695
rect 46891 5661 46900 5695
rect 46848 5652 46900 5661
rect 46940 5695 46992 5704
rect 46940 5661 46949 5695
rect 46949 5661 46983 5695
rect 46983 5661 46992 5695
rect 46940 5652 46992 5661
rect 47308 5695 47360 5704
rect 47308 5661 47317 5695
rect 47317 5661 47351 5695
rect 47351 5661 47360 5695
rect 47308 5652 47360 5661
rect 50436 5652 50488 5704
rect 51080 5652 51132 5704
rect 81440 5695 81492 5704
rect 81440 5661 81449 5695
rect 81449 5661 81483 5695
rect 81483 5661 81492 5695
rect 81440 5652 81492 5661
rect 41328 5516 41380 5568
rect 44456 5516 44508 5568
rect 44548 5559 44600 5568
rect 44548 5525 44557 5559
rect 44557 5525 44591 5559
rect 44591 5525 44600 5559
rect 44548 5516 44600 5525
rect 46664 5516 46716 5568
rect 47676 5559 47728 5568
rect 47676 5525 47685 5559
rect 47685 5525 47719 5559
rect 47719 5525 47728 5559
rect 47676 5516 47728 5525
rect 50528 5559 50580 5568
rect 50528 5525 50537 5559
rect 50537 5525 50571 5559
rect 50571 5525 50580 5559
rect 50528 5516 50580 5525
rect 50988 5584 51040 5636
rect 86776 5652 86828 5704
rect 84936 5584 84988 5636
rect 85580 5627 85632 5636
rect 79416 5516 79468 5568
rect 85580 5593 85589 5627
rect 85589 5593 85623 5627
rect 85623 5593 85632 5627
rect 85580 5584 85632 5593
rect 92664 5695 92716 5704
rect 92664 5661 92673 5695
rect 92673 5661 92707 5695
rect 92707 5661 92716 5695
rect 92664 5652 92716 5661
rect 94504 5695 94556 5704
rect 94504 5661 94513 5695
rect 94513 5661 94547 5695
rect 94547 5661 94556 5695
rect 94504 5652 94556 5661
rect 100576 5652 100628 5704
rect 100944 5652 100996 5704
rect 102784 5652 102836 5704
rect 92848 5627 92900 5636
rect 92848 5593 92857 5627
rect 92857 5593 92891 5627
rect 92891 5593 92900 5627
rect 92848 5584 92900 5593
rect 93400 5584 93452 5636
rect 101864 5584 101916 5636
rect 103152 5627 103204 5636
rect 103152 5593 103161 5627
rect 103161 5593 103195 5627
rect 103195 5593 103204 5627
rect 103152 5584 103204 5593
rect 104716 5584 104768 5636
rect 88064 5516 88116 5568
rect 92480 5516 92532 5568
rect 95056 5516 95108 5568
rect 102048 5516 102100 5568
rect 109316 5584 109368 5636
rect 111248 5652 111300 5704
rect 111800 5652 111852 5704
rect 115112 5652 115164 5704
rect 116768 5652 116820 5704
rect 119068 5695 119120 5704
rect 119068 5661 119077 5695
rect 119077 5661 119111 5695
rect 119111 5661 119120 5695
rect 119068 5652 119120 5661
rect 120080 5695 120132 5704
rect 120080 5661 120089 5695
rect 120089 5661 120123 5695
rect 120123 5661 120132 5695
rect 120080 5652 120132 5661
rect 156972 5788 157024 5840
rect 180984 5899 181036 5908
rect 180984 5865 180993 5899
rect 180993 5865 181027 5899
rect 181027 5865 181036 5899
rect 180984 5856 181036 5865
rect 182916 5899 182968 5908
rect 182916 5865 182925 5899
rect 182925 5865 182959 5899
rect 182959 5865 182968 5899
rect 182916 5856 182968 5865
rect 130200 5763 130252 5772
rect 130200 5729 130209 5763
rect 130209 5729 130243 5763
rect 130243 5729 130252 5763
rect 130200 5720 130252 5729
rect 143080 5763 143132 5772
rect 143080 5729 143089 5763
rect 143089 5729 143123 5763
rect 143123 5729 143132 5763
rect 143080 5720 143132 5729
rect 143356 5720 143408 5772
rect 143540 5763 143592 5772
rect 143540 5729 143549 5763
rect 143549 5729 143583 5763
rect 143583 5729 143592 5763
rect 143540 5720 143592 5729
rect 144460 5720 144512 5772
rect 147588 5720 147640 5772
rect 148232 5763 148284 5772
rect 148232 5729 148241 5763
rect 148241 5729 148275 5763
rect 148275 5729 148284 5763
rect 148232 5720 148284 5729
rect 112628 5584 112680 5636
rect 114376 5584 114428 5636
rect 119436 5627 119488 5636
rect 119436 5593 119445 5627
rect 119445 5593 119479 5627
rect 119479 5593 119488 5627
rect 119436 5584 119488 5593
rect 129924 5695 129976 5704
rect 129924 5661 129933 5695
rect 129933 5661 129967 5695
rect 129967 5661 129976 5695
rect 129924 5652 129976 5661
rect 145196 5652 145248 5704
rect 148048 5652 148100 5704
rect 142620 5584 142672 5636
rect 143540 5584 143592 5636
rect 148140 5584 148192 5636
rect 148416 5627 148468 5636
rect 148416 5593 148425 5627
rect 148425 5593 148459 5627
rect 148459 5593 148468 5627
rect 148416 5584 148468 5593
rect 122196 5516 122248 5568
rect 125140 5559 125192 5568
rect 125140 5525 125149 5559
rect 125149 5525 125183 5559
rect 125183 5525 125192 5559
rect 125140 5516 125192 5525
rect 147588 5516 147640 5568
rect 152740 5720 152792 5772
rect 155040 5720 155092 5772
rect 152004 5559 152056 5568
rect 152004 5525 152013 5559
rect 152013 5525 152047 5559
rect 152047 5525 152056 5559
rect 153384 5695 153436 5704
rect 153384 5661 153393 5695
rect 153393 5661 153427 5695
rect 153427 5661 153436 5695
rect 153384 5652 153436 5661
rect 155684 5695 155736 5704
rect 155684 5661 155693 5695
rect 155693 5661 155727 5695
rect 155727 5661 155736 5695
rect 155684 5652 155736 5661
rect 160652 5652 160704 5704
rect 161296 5720 161348 5772
rect 153292 5584 153344 5636
rect 155868 5627 155920 5636
rect 155868 5593 155877 5627
rect 155877 5593 155911 5627
rect 155911 5593 155920 5627
rect 155868 5584 155920 5593
rect 152004 5516 152056 5525
rect 162032 5584 162084 5636
rect 162768 5627 162820 5636
rect 162768 5593 162777 5627
rect 162777 5593 162811 5627
rect 162811 5593 162820 5627
rect 162768 5584 162820 5593
rect 158076 5516 158128 5568
rect 160560 5559 160612 5568
rect 160560 5525 160569 5559
rect 160569 5525 160603 5559
rect 160603 5525 160612 5559
rect 160560 5516 160612 5525
rect 160652 5516 160704 5568
rect 161296 5516 161348 5568
rect 162584 5516 162636 5568
rect 177028 5516 177080 5568
rect 177948 5516 178000 5568
rect 181812 5788 181864 5840
rect 216036 5856 216088 5908
rect 182180 5720 182232 5772
rect 182088 5695 182140 5704
rect 182088 5661 182097 5695
rect 182097 5661 182131 5695
rect 182131 5661 182140 5695
rect 182088 5652 182140 5661
rect 182548 5652 182600 5704
rect 200764 5788 200816 5840
rect 221004 5856 221056 5908
rect 186320 5516 186372 5568
rect 223764 5856 223816 5908
rect 224224 5856 224276 5908
rect 215392 5763 215444 5772
rect 215392 5729 215401 5763
rect 215401 5729 215435 5763
rect 215435 5729 215444 5763
rect 215392 5720 215444 5729
rect 215944 5720 215996 5772
rect 216128 5720 216180 5772
rect 218888 5720 218940 5772
rect 222016 5720 222068 5772
rect 223396 5788 223448 5840
rect 224592 5788 224644 5840
rect 226156 5856 226208 5908
rect 226248 5856 226300 5908
rect 227628 5856 227680 5908
rect 212540 5695 212592 5704
rect 212540 5661 212549 5695
rect 212549 5661 212583 5695
rect 212583 5661 212592 5695
rect 212540 5652 212592 5661
rect 214656 5695 214708 5704
rect 214656 5661 214665 5695
rect 214665 5661 214699 5695
rect 214699 5661 214708 5695
rect 214656 5652 214708 5661
rect 215576 5695 215628 5704
rect 215576 5661 215585 5695
rect 215585 5661 215619 5695
rect 215619 5661 215628 5695
rect 215576 5652 215628 5661
rect 216312 5695 216364 5704
rect 216312 5661 216321 5695
rect 216321 5661 216355 5695
rect 216355 5661 216364 5695
rect 216312 5652 216364 5661
rect 216496 5652 216548 5704
rect 223580 5652 223632 5704
rect 226064 5720 226116 5772
rect 229560 5856 229612 5908
rect 231308 5856 231360 5908
rect 231400 5856 231452 5908
rect 258356 5856 258408 5908
rect 261116 5856 261168 5908
rect 261208 5856 261260 5908
rect 244188 5788 244240 5840
rect 258816 5788 258868 5840
rect 260104 5788 260156 5840
rect 262680 5788 262732 5840
rect 270500 5856 270552 5908
rect 267740 5788 267792 5840
rect 225052 5652 225104 5704
rect 226524 5695 226576 5704
rect 226524 5661 226558 5695
rect 226558 5661 226576 5695
rect 226524 5652 226576 5661
rect 226708 5695 226760 5704
rect 226708 5661 226717 5695
rect 226717 5661 226751 5695
rect 226751 5661 226760 5695
rect 226708 5652 226760 5661
rect 227720 5695 227772 5704
rect 227720 5661 227729 5695
rect 227729 5661 227763 5695
rect 227763 5661 227772 5695
rect 227720 5652 227772 5661
rect 228088 5695 228140 5704
rect 228088 5661 228097 5695
rect 228097 5661 228131 5695
rect 228131 5661 228140 5695
rect 228088 5652 228140 5661
rect 209964 5584 210016 5636
rect 213000 5627 213052 5636
rect 213000 5593 213009 5627
rect 213009 5593 213043 5627
rect 213043 5593 213052 5627
rect 213000 5584 213052 5593
rect 215484 5584 215536 5636
rect 217140 5584 217192 5636
rect 219256 5584 219308 5636
rect 222016 5627 222068 5636
rect 222016 5593 222025 5627
rect 222025 5593 222059 5627
rect 222059 5593 222068 5627
rect 222016 5584 222068 5593
rect 222292 5584 222344 5636
rect 222844 5584 222896 5636
rect 223304 5584 223356 5636
rect 224868 5584 224920 5636
rect 228456 5627 228508 5636
rect 214656 5516 214708 5568
rect 215944 5516 215996 5568
rect 216036 5516 216088 5568
rect 228456 5593 228465 5627
rect 228465 5593 228499 5627
rect 228499 5593 228508 5627
rect 228456 5584 228508 5593
rect 227352 5559 227404 5568
rect 227352 5525 227361 5559
rect 227361 5525 227395 5559
rect 227395 5525 227404 5559
rect 227352 5516 227404 5525
rect 231216 5720 231268 5772
rect 230020 5652 230072 5704
rect 231492 5695 231544 5704
rect 231492 5661 231501 5695
rect 231501 5661 231535 5695
rect 231535 5661 231544 5695
rect 231492 5652 231544 5661
rect 231860 5720 231912 5772
rect 259276 5720 259328 5772
rect 232320 5695 232372 5704
rect 232320 5661 232329 5695
rect 232329 5661 232363 5695
rect 232363 5661 232372 5695
rect 232320 5652 232372 5661
rect 228916 5584 228968 5636
rect 229836 5584 229888 5636
rect 229928 5584 229980 5636
rect 230664 5627 230716 5636
rect 230664 5593 230673 5627
rect 230673 5593 230707 5627
rect 230707 5593 230716 5627
rect 230664 5584 230716 5593
rect 230848 5627 230900 5636
rect 230848 5593 230873 5627
rect 230873 5593 230900 5627
rect 230848 5584 230900 5593
rect 256884 5652 256936 5704
rect 237380 5584 237432 5636
rect 259092 5584 259144 5636
rect 252284 5516 252336 5568
rect 258816 5516 258868 5568
rect 262220 5720 262272 5772
rect 263140 5763 263192 5772
rect 263140 5729 263149 5763
rect 263149 5729 263183 5763
rect 263183 5729 263192 5763
rect 263140 5720 263192 5729
rect 261668 5695 261720 5704
rect 261668 5661 261677 5695
rect 261677 5661 261711 5695
rect 261711 5661 261720 5695
rect 261668 5652 261720 5661
rect 266728 5720 266780 5772
rect 264060 5695 264112 5704
rect 264060 5661 264069 5695
rect 264069 5661 264103 5695
rect 264103 5661 264112 5695
rect 264060 5652 264112 5661
rect 264520 5695 264572 5704
rect 264520 5661 264529 5695
rect 264529 5661 264563 5695
rect 264563 5661 264572 5695
rect 264520 5652 264572 5661
rect 265256 5695 265308 5704
rect 265256 5661 265265 5695
rect 265265 5661 265299 5695
rect 265299 5661 265308 5695
rect 265256 5652 265308 5661
rect 261116 5584 261168 5636
rect 263140 5584 263192 5636
rect 263600 5584 263652 5636
rect 264888 5584 264940 5636
rect 265900 5584 265952 5636
rect 266176 5584 266228 5636
rect 267188 5695 267240 5704
rect 267188 5661 267197 5695
rect 267197 5661 267231 5695
rect 267231 5661 267240 5695
rect 267188 5652 267240 5661
rect 269028 5652 269080 5704
rect 269488 5695 269540 5704
rect 269488 5661 269497 5695
rect 269497 5661 269531 5695
rect 269531 5661 269540 5695
rect 269488 5652 269540 5661
rect 268660 5584 268712 5636
rect 268844 5627 268896 5636
rect 268844 5593 268853 5627
rect 268853 5593 268887 5627
rect 268887 5593 268896 5627
rect 268844 5584 268896 5593
rect 269212 5584 269264 5636
rect 261944 5516 261996 5568
rect 266360 5516 266412 5568
rect 270408 5652 270460 5704
rect 68546 5414 68598 5466
rect 68610 5414 68662 5466
rect 68674 5414 68726 5466
rect 68738 5414 68790 5466
rect 68802 5414 68854 5466
rect 136143 5414 136195 5466
rect 136207 5414 136259 5466
rect 136271 5414 136323 5466
rect 136335 5414 136387 5466
rect 136399 5414 136451 5466
rect 203740 5414 203792 5466
rect 203804 5414 203856 5466
rect 203868 5414 203920 5466
rect 203932 5414 203984 5466
rect 203996 5414 204048 5466
rect 271337 5414 271389 5466
rect 271401 5414 271453 5466
rect 271465 5414 271517 5466
rect 271529 5414 271581 5466
rect 271593 5414 271645 5466
rect 15292 5312 15344 5364
rect 34612 5312 34664 5364
rect 26884 5244 26936 5296
rect 37832 5244 37884 5296
rect 37924 5287 37976 5296
rect 37924 5253 37933 5287
rect 37933 5253 37967 5287
rect 37967 5253 37976 5287
rect 37924 5244 37976 5253
rect 43536 5312 43588 5364
rect 45376 5312 45428 5364
rect 38752 5287 38804 5296
rect 38752 5253 38761 5287
rect 38761 5253 38795 5287
rect 38795 5253 38804 5287
rect 38752 5244 38804 5253
rect 43352 5287 43404 5296
rect 43352 5253 43361 5287
rect 43361 5253 43395 5287
rect 43395 5253 43404 5287
rect 43352 5244 43404 5253
rect 43720 5287 43772 5296
rect 43720 5253 43729 5287
rect 43729 5253 43763 5287
rect 43763 5253 43772 5287
rect 43720 5244 43772 5253
rect 44364 5244 44416 5296
rect 45836 5287 45888 5296
rect 45836 5253 45845 5287
rect 45845 5253 45879 5287
rect 45879 5253 45888 5287
rect 45836 5244 45888 5253
rect 46112 5287 46164 5296
rect 46112 5253 46121 5287
rect 46121 5253 46155 5287
rect 46155 5253 46164 5287
rect 46112 5244 46164 5253
rect 46848 5312 46900 5364
rect 46296 5244 46348 5296
rect 38200 5176 38252 5228
rect 42616 5176 42668 5228
rect 43812 5176 43864 5228
rect 45928 5176 45980 5228
rect 47952 5219 48004 5228
rect 47952 5185 47961 5219
rect 47961 5185 47995 5219
rect 47995 5185 48004 5219
rect 47952 5176 48004 5185
rect 49332 5176 49384 5228
rect 50712 5244 50764 5296
rect 51172 5244 51224 5296
rect 51356 5287 51408 5296
rect 51356 5253 51365 5287
rect 51365 5253 51399 5287
rect 51399 5253 51408 5287
rect 51356 5244 51408 5253
rect 51448 5244 51500 5296
rect 50988 5219 51040 5228
rect 50988 5185 50997 5219
rect 50997 5185 51031 5219
rect 51031 5185 51040 5219
rect 50988 5176 51040 5185
rect 38476 5108 38528 5160
rect 40776 5108 40828 5160
rect 41144 5108 41196 5160
rect 42432 5108 42484 5160
rect 44732 5108 44784 5160
rect 48044 5108 48096 5160
rect 51632 5108 51684 5160
rect 42892 5040 42944 5092
rect 44640 5083 44692 5092
rect 44640 5049 44649 5083
rect 44649 5049 44683 5083
rect 44683 5049 44692 5083
rect 44640 5040 44692 5049
rect 53104 5355 53156 5364
rect 53104 5321 53113 5355
rect 53113 5321 53147 5355
rect 53147 5321 53156 5355
rect 53104 5312 53156 5321
rect 52092 5244 52144 5296
rect 80336 5287 80388 5296
rect 80336 5253 80345 5287
rect 80345 5253 80379 5287
rect 80379 5253 80388 5287
rect 80336 5244 80388 5253
rect 81348 5244 81400 5296
rect 80796 5219 80848 5228
rect 80796 5185 80805 5219
rect 80805 5185 80839 5219
rect 80839 5185 80848 5219
rect 80796 5176 80848 5185
rect 80888 5219 80940 5228
rect 80888 5185 80897 5219
rect 80897 5185 80931 5219
rect 80931 5185 80940 5219
rect 80888 5176 80940 5185
rect 81624 5287 81676 5296
rect 81624 5253 81633 5287
rect 81633 5253 81667 5287
rect 81667 5253 81676 5287
rect 81624 5244 81676 5253
rect 82912 5244 82964 5296
rect 84752 5244 84804 5296
rect 84936 5287 84988 5296
rect 84936 5253 84945 5287
rect 84945 5253 84979 5287
rect 84979 5253 84988 5287
rect 84936 5244 84988 5253
rect 86592 5287 86644 5296
rect 86592 5253 86601 5287
rect 86601 5253 86635 5287
rect 86635 5253 86644 5287
rect 86592 5244 86644 5253
rect 93860 5244 93912 5296
rect 101312 5312 101364 5364
rect 108764 5312 108816 5364
rect 110696 5312 110748 5364
rect 115020 5312 115072 5364
rect 120080 5312 120132 5364
rect 142804 5312 142856 5364
rect 152372 5312 152424 5364
rect 153384 5312 153436 5364
rect 157800 5355 157852 5364
rect 114376 5244 114428 5296
rect 116308 5244 116360 5296
rect 100944 5176 100996 5228
rect 84660 5108 84712 5160
rect 84752 5151 84804 5160
rect 84752 5117 84761 5151
rect 84761 5117 84795 5151
rect 84795 5117 84804 5151
rect 84752 5108 84804 5117
rect 89536 5040 89588 5092
rect 91744 5151 91796 5160
rect 91744 5117 91753 5151
rect 91753 5117 91787 5151
rect 91787 5117 91796 5151
rect 91744 5108 91796 5117
rect 91928 5151 91980 5160
rect 91928 5117 91937 5151
rect 91937 5117 91971 5151
rect 91971 5117 91980 5151
rect 91928 5108 91980 5117
rect 92664 5108 92716 5160
rect 100668 5108 100720 5160
rect 107016 5219 107068 5228
rect 107016 5185 107025 5219
rect 107025 5185 107059 5219
rect 107059 5185 107068 5219
rect 107016 5176 107068 5185
rect 107200 5176 107252 5228
rect 107292 5219 107344 5228
rect 107292 5185 107301 5219
rect 107301 5185 107335 5219
rect 107335 5185 107344 5219
rect 107292 5176 107344 5185
rect 117412 5219 117464 5228
rect 117412 5185 117421 5219
rect 117421 5185 117455 5219
rect 117455 5185 117464 5219
rect 117412 5176 117464 5185
rect 120264 5244 120316 5296
rect 150532 5244 150584 5296
rect 153292 5287 153344 5296
rect 153292 5253 153301 5287
rect 153301 5253 153335 5287
rect 153335 5253 153344 5287
rect 153292 5244 153344 5253
rect 121000 5219 121052 5228
rect 121000 5185 121009 5219
rect 121009 5185 121043 5219
rect 121043 5185 121052 5219
rect 121000 5176 121052 5185
rect 122196 5219 122248 5228
rect 122196 5185 122205 5219
rect 122205 5185 122239 5219
rect 122239 5185 122248 5219
rect 122196 5176 122248 5185
rect 123484 5176 123536 5228
rect 102048 5040 102100 5092
rect 108396 5108 108448 5160
rect 110604 5108 110656 5160
rect 17132 4972 17184 5024
rect 33232 4972 33284 5024
rect 40316 4972 40368 5024
rect 42064 4972 42116 5024
rect 47860 4972 47912 5024
rect 51908 5015 51960 5024
rect 51908 4981 51917 5015
rect 51917 4981 51951 5015
rect 51951 4981 51960 5015
rect 51908 4972 51960 4981
rect 52000 4972 52052 5024
rect 78128 4972 78180 5024
rect 84660 5015 84712 5024
rect 84660 4981 84669 5015
rect 84669 4981 84703 5015
rect 84703 4981 84712 5015
rect 84660 4972 84712 4981
rect 84844 4972 84896 5024
rect 89904 4972 89956 5024
rect 94136 4972 94188 5024
rect 99656 4972 99708 5024
rect 103520 4972 103572 5024
rect 106648 5040 106700 5092
rect 105820 4972 105872 5024
rect 111984 5151 112036 5160
rect 111984 5117 111993 5151
rect 111993 5117 112027 5151
rect 112027 5117 112036 5151
rect 111984 5108 112036 5117
rect 112444 5083 112496 5092
rect 107936 5015 107988 5024
rect 107936 4981 107945 5015
rect 107945 4981 107979 5015
rect 107979 4981 107988 5015
rect 107936 4972 107988 4981
rect 110236 4972 110288 5024
rect 112444 5049 112453 5083
rect 112453 5049 112487 5083
rect 112487 5049 112496 5083
rect 112444 5040 112496 5049
rect 112812 5151 112864 5160
rect 112812 5117 112846 5151
rect 112846 5117 112864 5151
rect 112812 5108 112864 5117
rect 113180 5108 113232 5160
rect 114192 5108 114244 5160
rect 114284 5040 114336 5092
rect 116768 5108 116820 5160
rect 117596 5151 117648 5160
rect 117596 5117 117605 5151
rect 117605 5117 117639 5151
rect 117639 5117 117648 5151
rect 117596 5108 117648 5117
rect 118332 5151 118384 5160
rect 118332 5117 118359 5151
rect 118359 5117 118384 5151
rect 118332 5108 118384 5117
rect 118516 5108 118568 5160
rect 119436 5108 119488 5160
rect 120448 5108 120500 5160
rect 120816 5108 120868 5160
rect 118056 5083 118108 5092
rect 113640 5015 113692 5024
rect 113640 4981 113649 5015
rect 113649 4981 113683 5015
rect 113683 4981 113692 5015
rect 113640 4972 113692 4981
rect 113732 4972 113784 5024
rect 115296 4972 115348 5024
rect 118056 5049 118065 5083
rect 118065 5049 118099 5083
rect 118099 5049 118108 5083
rect 118056 5040 118108 5049
rect 117412 4972 117464 5024
rect 120724 5083 120776 5092
rect 120724 5049 120733 5083
rect 120733 5049 120767 5083
rect 120767 5049 120776 5083
rect 120724 5040 120776 5049
rect 119436 4972 119488 5024
rect 120356 4972 120408 5024
rect 121920 5015 121972 5024
rect 121920 4981 121929 5015
rect 121929 4981 121963 5015
rect 121963 4981 121972 5015
rect 121920 4972 121972 4981
rect 149888 5176 149940 5228
rect 157800 5321 157809 5355
rect 157809 5321 157843 5355
rect 157843 5321 157852 5355
rect 157800 5312 157852 5321
rect 159456 5244 159508 5296
rect 162584 5287 162636 5296
rect 162584 5253 162593 5287
rect 162593 5253 162627 5287
rect 162627 5253 162636 5287
rect 162584 5244 162636 5253
rect 163044 5355 163096 5364
rect 163044 5321 163053 5355
rect 163053 5321 163087 5355
rect 163087 5321 163096 5355
rect 163044 5312 163096 5321
rect 163228 5312 163280 5364
rect 175924 5312 175976 5364
rect 188436 5287 188488 5296
rect 188436 5253 188445 5287
rect 188445 5253 188479 5287
rect 188479 5253 188488 5287
rect 188436 5244 188488 5253
rect 150808 5151 150860 5160
rect 150808 5117 150817 5151
rect 150817 5117 150851 5151
rect 150851 5117 150860 5151
rect 150808 5108 150860 5117
rect 150900 5108 150952 5160
rect 151360 5108 151412 5160
rect 151728 5108 151780 5160
rect 151820 5151 151872 5160
rect 151820 5117 151829 5151
rect 151829 5117 151863 5151
rect 151863 5117 151872 5151
rect 151820 5108 151872 5117
rect 152372 5108 152424 5160
rect 161112 5219 161164 5228
rect 161112 5185 161121 5219
rect 161121 5185 161155 5219
rect 161155 5185 161164 5219
rect 161112 5176 161164 5185
rect 161388 5176 161440 5228
rect 161572 5219 161624 5228
rect 161572 5185 161581 5219
rect 161581 5185 161615 5219
rect 161615 5185 161624 5219
rect 161572 5176 161624 5185
rect 155868 5108 155920 5160
rect 153752 4972 153804 5024
rect 158076 5040 158128 5092
rect 158260 5151 158312 5160
rect 158260 5117 158269 5151
rect 158269 5117 158303 5151
rect 158303 5117 158312 5151
rect 158260 5108 158312 5117
rect 158536 5108 158588 5160
rect 160008 5151 160060 5160
rect 160008 5117 160017 5151
rect 160017 5117 160051 5151
rect 160051 5117 160060 5151
rect 160008 5108 160060 5117
rect 161204 5040 161256 5092
rect 162124 5083 162176 5092
rect 162124 5049 162133 5083
rect 162133 5049 162167 5083
rect 162167 5049 162176 5083
rect 162124 5040 162176 5049
rect 162676 5108 162728 5160
rect 156052 4972 156104 5024
rect 156788 4972 156840 5024
rect 158628 4972 158680 5024
rect 160008 4972 160060 5024
rect 161572 4972 161624 5024
rect 162952 4972 163004 5024
rect 163504 5176 163556 5228
rect 180616 5176 180668 5228
rect 182088 5176 182140 5228
rect 182180 5219 182232 5228
rect 182180 5185 182189 5219
rect 182189 5185 182223 5219
rect 182223 5185 182232 5219
rect 182180 5176 182232 5185
rect 182548 5219 182600 5228
rect 182548 5185 182557 5219
rect 182557 5185 182591 5219
rect 182591 5185 182600 5219
rect 182548 5176 182600 5185
rect 189172 5287 189224 5296
rect 189172 5253 189181 5287
rect 189181 5253 189215 5287
rect 189215 5253 189224 5287
rect 189172 5244 189224 5253
rect 215852 5312 215904 5364
rect 218152 5312 218204 5364
rect 220176 5244 220228 5296
rect 224684 5287 224736 5296
rect 224684 5253 224693 5287
rect 224693 5253 224727 5287
rect 224727 5253 224736 5287
rect 224684 5244 224736 5253
rect 177948 5108 178000 5160
rect 164240 5040 164292 5092
rect 175832 5040 175884 5092
rect 182548 5083 182600 5092
rect 182548 5049 182557 5083
rect 182557 5049 182591 5083
rect 182591 5049 182600 5083
rect 182548 5040 182600 5049
rect 214012 5151 214064 5160
rect 214012 5117 214021 5151
rect 214021 5117 214055 5151
rect 214055 5117 214064 5151
rect 214012 5108 214064 5117
rect 214196 5151 214248 5160
rect 214196 5117 214205 5151
rect 214205 5117 214239 5151
rect 214239 5117 214248 5151
rect 214196 5108 214248 5117
rect 216588 5108 216640 5160
rect 219256 5219 219308 5228
rect 219256 5185 219265 5219
rect 219265 5185 219299 5219
rect 219299 5185 219308 5219
rect 219256 5176 219308 5185
rect 222292 5219 222344 5228
rect 222292 5185 222301 5219
rect 222301 5185 222335 5219
rect 222335 5185 222344 5219
rect 222292 5176 222344 5185
rect 222384 5176 222436 5228
rect 227352 5244 227404 5296
rect 227536 5287 227588 5296
rect 227536 5253 227545 5287
rect 227545 5253 227579 5287
rect 227579 5253 227588 5287
rect 227536 5244 227588 5253
rect 228272 5244 228324 5296
rect 228824 5244 228876 5296
rect 230848 5244 230900 5296
rect 238668 5312 238720 5364
rect 239220 5244 239272 5296
rect 230020 5219 230072 5228
rect 230020 5185 230029 5219
rect 230029 5185 230063 5219
rect 230063 5185 230072 5219
rect 230020 5176 230072 5185
rect 230480 5176 230532 5228
rect 231860 5176 231912 5228
rect 238668 5219 238720 5228
rect 238668 5185 238677 5219
rect 238677 5185 238711 5219
rect 238711 5185 238720 5219
rect 238668 5176 238720 5185
rect 239312 5176 239364 5228
rect 223856 5108 223908 5160
rect 225972 5108 226024 5160
rect 226800 5108 226852 5160
rect 215024 5040 215076 5092
rect 215944 5040 215996 5092
rect 189264 4972 189316 5024
rect 190000 4972 190052 5024
rect 210056 4972 210108 5024
rect 218704 4972 218756 5024
rect 226340 5040 226392 5092
rect 239220 5108 239272 5160
rect 230664 5040 230716 5092
rect 231032 5040 231084 5092
rect 239680 5244 239732 5296
rect 255780 5244 255832 5296
rect 239588 5176 239640 5228
rect 251456 5176 251508 5228
rect 253572 5108 253624 5160
rect 262220 5312 262272 5364
rect 266728 5312 266780 5364
rect 267740 5355 267792 5364
rect 267740 5321 267749 5355
rect 267749 5321 267783 5355
rect 267783 5321 267792 5355
rect 267740 5312 267792 5321
rect 267832 5312 267884 5364
rect 269028 5312 269080 5364
rect 271144 5312 271196 5364
rect 271972 5312 272024 5364
rect 261944 5244 261996 5296
rect 267280 5244 267332 5296
rect 262496 5176 262548 5228
rect 262956 5219 263008 5228
rect 262956 5185 262965 5219
rect 262965 5185 262999 5219
rect 262999 5185 263008 5219
rect 262956 5176 263008 5185
rect 264704 5219 264756 5228
rect 264704 5185 264713 5219
rect 264713 5185 264747 5219
rect 264747 5185 264756 5219
rect 264704 5176 264756 5185
rect 265992 5219 266044 5228
rect 265992 5185 266001 5219
rect 266001 5185 266035 5219
rect 266035 5185 266044 5219
rect 265992 5176 266044 5185
rect 266176 5176 266228 5228
rect 267464 5176 267516 5228
rect 268660 5176 268712 5228
rect 269764 5176 269816 5228
rect 270408 5176 270460 5228
rect 260656 5151 260708 5160
rect 260656 5117 260665 5151
rect 260665 5117 260699 5151
rect 260699 5117 260708 5151
rect 260656 5108 260708 5117
rect 263232 5151 263284 5160
rect 263232 5117 263241 5151
rect 263241 5117 263275 5151
rect 263275 5117 263284 5151
rect 263232 5108 263284 5117
rect 224868 4972 224920 5024
rect 225236 4972 225288 5024
rect 227536 4972 227588 5024
rect 227720 4972 227772 5024
rect 229008 4972 229060 5024
rect 231308 5015 231360 5024
rect 231308 4981 231317 5015
rect 231317 4981 231351 5015
rect 231351 4981 231360 5015
rect 231308 4972 231360 4981
rect 235632 4972 235684 5024
rect 239220 4972 239272 5024
rect 239588 4972 239640 5024
rect 264428 5040 264480 5092
rect 265164 5108 265216 5160
rect 268292 5151 268344 5160
rect 268292 5117 268301 5151
rect 268301 5117 268335 5151
rect 268335 5117 268344 5151
rect 268292 5108 268344 5117
rect 269304 5151 269356 5160
rect 269304 5117 269313 5151
rect 269313 5117 269347 5151
rect 269347 5117 269356 5151
rect 269304 5108 269356 5117
rect 266636 5040 266688 5092
rect 267464 5040 267516 5092
rect 268844 5040 268896 5092
rect 269212 5040 269264 5092
rect 242256 5015 242308 5024
rect 242256 4981 242265 5015
rect 242265 4981 242299 5015
rect 242299 4981 242308 5015
rect 242256 4972 242308 4981
rect 242624 5015 242676 5024
rect 242624 4981 242633 5015
rect 242633 4981 242667 5015
rect 242667 4981 242676 5015
rect 242624 4972 242676 4981
rect 242716 4972 242768 5024
rect 245568 4972 245620 5024
rect 252468 4972 252520 5024
rect 256884 4972 256936 5024
rect 258540 4972 258592 5024
rect 259460 5015 259512 5024
rect 259460 4981 259469 5015
rect 259469 4981 259503 5015
rect 259503 4981 259512 5015
rect 259460 4972 259512 4981
rect 266820 4972 266872 5024
rect 271972 4972 272024 5024
rect 34748 4870 34800 4922
rect 34812 4870 34864 4922
rect 34876 4870 34928 4922
rect 34940 4870 34992 4922
rect 35004 4870 35056 4922
rect 102345 4870 102397 4922
rect 102409 4870 102461 4922
rect 102473 4870 102525 4922
rect 102537 4870 102589 4922
rect 102601 4870 102653 4922
rect 169942 4870 169994 4922
rect 170006 4870 170058 4922
rect 170070 4870 170122 4922
rect 170134 4870 170186 4922
rect 170198 4870 170250 4922
rect 237539 4870 237591 4922
rect 237603 4870 237655 4922
rect 237667 4870 237719 4922
rect 237731 4870 237783 4922
rect 237795 4870 237847 4922
rect 12164 4768 12216 4820
rect 35900 4768 35952 4820
rect 34612 4700 34664 4752
rect 39764 4700 39816 4752
rect 33140 4632 33192 4684
rect 40960 4768 41012 4820
rect 42524 4768 42576 4820
rect 52092 4768 52144 4820
rect 74540 4768 74592 4820
rect 82912 4768 82964 4820
rect 84660 4768 84712 4820
rect 51172 4700 51224 4752
rect 52000 4700 52052 4752
rect 41144 4632 41196 4684
rect 44732 4632 44784 4684
rect 48044 4632 48096 4684
rect 53104 4632 53156 4684
rect 36544 4564 36596 4616
rect 8484 4428 8536 4480
rect 40316 4428 40368 4480
rect 40960 4471 41012 4480
rect 40960 4437 40969 4471
rect 40969 4437 41003 4471
rect 41003 4437 41012 4471
rect 40960 4428 41012 4437
rect 41236 4539 41288 4548
rect 41236 4505 41245 4539
rect 41245 4505 41279 4539
rect 41279 4505 41288 4539
rect 41236 4496 41288 4505
rect 41604 4496 41656 4548
rect 42064 4539 42116 4548
rect 42064 4505 42073 4539
rect 42073 4505 42107 4539
rect 42107 4505 42116 4539
rect 42064 4496 42116 4505
rect 43260 4607 43312 4616
rect 43260 4573 43269 4607
rect 43269 4573 43303 4607
rect 43303 4573 43312 4607
rect 43260 4564 43312 4573
rect 43628 4564 43680 4616
rect 47768 4607 47820 4616
rect 47768 4573 47777 4607
rect 47777 4573 47811 4607
rect 47811 4573 47820 4607
rect 47768 4564 47820 4573
rect 48136 4564 48188 4616
rect 42248 4471 42300 4480
rect 42248 4437 42257 4471
rect 42257 4437 42291 4471
rect 42291 4437 42300 4471
rect 42248 4428 42300 4437
rect 43076 4428 43128 4480
rect 43996 4496 44048 4548
rect 46848 4496 46900 4548
rect 47216 4496 47268 4548
rect 47860 4539 47912 4548
rect 47860 4505 47869 4539
rect 47869 4505 47903 4539
rect 47903 4505 47912 4539
rect 47860 4496 47912 4505
rect 48228 4539 48280 4548
rect 48228 4505 48237 4539
rect 48237 4505 48271 4539
rect 48271 4505 48280 4539
rect 48228 4496 48280 4505
rect 44272 4471 44324 4480
rect 44272 4437 44281 4471
rect 44281 4437 44315 4471
rect 44315 4437 44324 4471
rect 44272 4428 44324 4437
rect 46940 4471 46992 4480
rect 46940 4437 46949 4471
rect 46949 4437 46983 4471
rect 46983 4437 46992 4471
rect 46940 4428 46992 4437
rect 48872 4496 48924 4548
rect 48596 4428 48648 4480
rect 50988 4428 51040 4480
rect 51356 4428 51408 4480
rect 52000 4428 52052 4480
rect 52276 4496 52328 4548
rect 52460 4539 52512 4548
rect 52460 4505 52469 4539
rect 52469 4505 52503 4539
rect 52503 4505 52512 4539
rect 52460 4496 52512 4505
rect 52828 4539 52880 4548
rect 52828 4505 52837 4539
rect 52837 4505 52871 4539
rect 52871 4505 52880 4539
rect 52828 4496 52880 4505
rect 84752 4700 84804 4752
rect 85580 4700 85632 4752
rect 86776 4700 86828 4752
rect 91008 4768 91060 4820
rect 99380 4700 99432 4752
rect 99840 4700 99892 4752
rect 78128 4632 78180 4684
rect 81900 4632 81952 4684
rect 92664 4675 92716 4684
rect 92664 4641 92673 4675
rect 92673 4641 92707 4675
rect 92707 4641 92716 4675
rect 92664 4632 92716 4641
rect 95240 4632 95292 4684
rect 100944 4700 100996 4752
rect 105544 4700 105596 4752
rect 106648 4700 106700 4752
rect 107660 4743 107712 4752
rect 107660 4709 107669 4743
rect 107669 4709 107703 4743
rect 107703 4709 107712 4743
rect 107660 4700 107712 4709
rect 109408 4743 109460 4752
rect 109408 4709 109417 4743
rect 109417 4709 109451 4743
rect 109451 4709 109460 4743
rect 109408 4700 109460 4709
rect 100576 4632 100628 4684
rect 106372 4632 106424 4684
rect 108396 4632 108448 4684
rect 110236 4700 110288 4752
rect 111800 4700 111852 4752
rect 112996 4700 113048 4752
rect 113732 4700 113784 4752
rect 113916 4768 113968 4820
rect 118884 4768 118936 4820
rect 120724 4700 120776 4752
rect 139308 4768 139360 4820
rect 153752 4768 153804 4820
rect 110696 4675 110748 4684
rect 110696 4641 110705 4675
rect 110705 4641 110739 4675
rect 110739 4641 110748 4675
rect 110696 4632 110748 4641
rect 84016 4607 84068 4616
rect 84016 4573 84025 4607
rect 84025 4573 84059 4607
rect 84059 4573 84068 4607
rect 84016 4564 84068 4573
rect 81624 4496 81676 4548
rect 53196 4471 53248 4480
rect 53196 4437 53205 4471
rect 53205 4437 53239 4471
rect 53239 4437 53248 4471
rect 53196 4428 53248 4437
rect 53380 4471 53432 4480
rect 53380 4437 53389 4471
rect 53389 4437 53423 4471
rect 53423 4437 53432 4471
rect 53380 4428 53432 4437
rect 85580 4496 85632 4548
rect 86408 4496 86460 4548
rect 87880 4607 87932 4616
rect 87880 4573 87889 4607
rect 87889 4573 87923 4607
rect 87923 4573 87932 4607
rect 87880 4564 87932 4573
rect 86684 4496 86736 4548
rect 87512 4471 87564 4480
rect 87512 4437 87521 4471
rect 87521 4437 87555 4471
rect 87555 4437 87564 4471
rect 87512 4428 87564 4437
rect 88064 4539 88116 4548
rect 88064 4505 88073 4539
rect 88073 4505 88107 4539
rect 88107 4505 88116 4539
rect 88064 4496 88116 4505
rect 94412 4607 94464 4616
rect 94412 4573 94421 4607
rect 94421 4573 94455 4607
rect 94455 4573 94464 4607
rect 94412 4564 94464 4573
rect 94964 4564 95016 4616
rect 105820 4564 105872 4616
rect 106280 4564 106332 4616
rect 108120 4564 108172 4616
rect 108212 4607 108264 4616
rect 108212 4573 108221 4607
rect 108221 4573 108255 4607
rect 108255 4573 108264 4607
rect 108212 4564 108264 4573
rect 109960 4607 110012 4616
rect 109960 4573 109969 4607
rect 109969 4573 110003 4607
rect 110003 4573 110012 4607
rect 109960 4564 110012 4573
rect 110972 4607 111024 4616
rect 110972 4573 110981 4607
rect 110981 4573 111015 4607
rect 111015 4573 111024 4607
rect 110972 4564 111024 4573
rect 92480 4428 92532 4480
rect 95056 4496 95108 4548
rect 99472 4539 99524 4548
rect 99472 4505 99481 4539
rect 99481 4505 99515 4539
rect 99515 4505 99524 4539
rect 99472 4496 99524 4505
rect 105452 4496 105504 4548
rect 108764 4496 108816 4548
rect 109868 4496 109920 4548
rect 113640 4632 113692 4684
rect 114376 4632 114428 4684
rect 114468 4632 114520 4684
rect 116216 4675 116268 4684
rect 116216 4641 116225 4675
rect 116225 4641 116259 4675
rect 116259 4641 116268 4675
rect 116216 4632 116268 4641
rect 118240 4675 118292 4684
rect 118240 4641 118249 4675
rect 118249 4641 118283 4675
rect 118283 4641 118292 4675
rect 118240 4632 118292 4641
rect 112536 4564 112588 4616
rect 113916 4564 113968 4616
rect 118056 4564 118108 4616
rect 119804 4632 119856 4684
rect 121920 4632 121972 4684
rect 142804 4700 142856 4752
rect 151084 4700 151136 4752
rect 144828 4632 144880 4684
rect 150440 4632 150492 4684
rect 150900 4632 150952 4684
rect 151176 4675 151228 4684
rect 151176 4641 151185 4675
rect 151185 4641 151219 4675
rect 151219 4641 151228 4675
rect 151176 4632 151228 4641
rect 152464 4700 152516 4752
rect 156604 4768 156656 4820
rect 157248 4768 157300 4820
rect 156052 4700 156104 4752
rect 151912 4632 151964 4684
rect 158536 4768 158588 4820
rect 160008 4768 160060 4820
rect 163228 4768 163280 4820
rect 179880 4768 179932 4820
rect 118424 4607 118476 4616
rect 118424 4573 118433 4607
rect 118433 4573 118467 4607
rect 118467 4573 118476 4607
rect 118424 4564 118476 4573
rect 119160 4607 119212 4616
rect 119160 4573 119169 4607
rect 119169 4573 119203 4607
rect 119203 4573 119212 4607
rect 119160 4564 119212 4573
rect 119252 4607 119304 4616
rect 119252 4573 119286 4607
rect 119286 4573 119304 4607
rect 119252 4564 119304 4573
rect 119436 4607 119488 4616
rect 119436 4573 119445 4607
rect 119445 4573 119479 4607
rect 119479 4573 119488 4607
rect 119436 4564 119488 4573
rect 115020 4496 115072 4548
rect 100208 4471 100260 4480
rect 100208 4437 100217 4471
rect 100217 4437 100251 4471
rect 100251 4437 100260 4471
rect 100208 4428 100260 4437
rect 101312 4428 101364 4480
rect 106280 4428 106332 4480
rect 108856 4471 108908 4480
rect 108856 4437 108865 4471
rect 108865 4437 108899 4471
rect 108899 4437 108908 4471
rect 108856 4428 108908 4437
rect 110972 4428 111024 4480
rect 113180 4428 113232 4480
rect 113364 4471 113416 4480
rect 113364 4437 113373 4471
rect 113373 4437 113407 4471
rect 113407 4437 113416 4471
rect 113364 4428 113416 4437
rect 114468 4428 114520 4480
rect 114652 4428 114704 4480
rect 116400 4428 116452 4480
rect 118884 4428 118936 4480
rect 120264 4428 120316 4480
rect 150716 4607 150768 4616
rect 150716 4573 150725 4607
rect 150725 4573 150759 4607
rect 150759 4573 150768 4607
rect 150716 4564 150768 4573
rect 151452 4607 151504 4616
rect 151452 4573 151461 4607
rect 151461 4573 151495 4607
rect 151495 4573 151504 4607
rect 151452 4564 151504 4573
rect 151636 4564 151688 4616
rect 152372 4607 152424 4616
rect 152372 4573 152381 4607
rect 152381 4573 152415 4607
rect 152415 4573 152424 4607
rect 152372 4564 152424 4573
rect 122656 4539 122708 4548
rect 122656 4505 122665 4539
rect 122665 4505 122699 4539
rect 122699 4505 122708 4539
rect 122656 4496 122708 4505
rect 142160 4496 142212 4548
rect 143356 4496 143408 4548
rect 145196 4539 145248 4548
rect 129924 4428 129976 4480
rect 142436 4471 142488 4480
rect 142436 4437 142445 4471
rect 142445 4437 142479 4471
rect 142479 4437 142488 4471
rect 145196 4505 145205 4539
rect 145205 4505 145239 4539
rect 145239 4505 145248 4539
rect 145196 4496 145248 4505
rect 152280 4496 152332 4548
rect 153384 4607 153436 4616
rect 153384 4573 153393 4607
rect 153393 4573 153427 4607
rect 153427 4573 153436 4607
rect 153384 4564 153436 4573
rect 154120 4607 154172 4616
rect 154120 4573 154129 4607
rect 154129 4573 154163 4607
rect 154163 4573 154172 4607
rect 154120 4564 154172 4573
rect 154304 4564 154356 4616
rect 154396 4607 154448 4616
rect 154396 4573 154405 4607
rect 154405 4573 154439 4607
rect 154439 4573 154448 4607
rect 154396 4564 154448 4573
rect 155868 4496 155920 4548
rect 156420 4496 156472 4548
rect 210700 4632 210752 4684
rect 213920 4768 213972 4820
rect 214012 4768 214064 4820
rect 219716 4811 219768 4820
rect 219716 4777 219725 4811
rect 219725 4777 219759 4811
rect 219759 4777 219768 4811
rect 219716 4768 219768 4777
rect 222476 4768 222528 4820
rect 223212 4768 223264 4820
rect 224684 4811 224736 4820
rect 224684 4777 224693 4811
rect 224693 4777 224727 4811
rect 224727 4777 224736 4811
rect 224684 4768 224736 4777
rect 226340 4768 226392 4820
rect 213460 4700 213512 4752
rect 215484 4700 215536 4752
rect 215852 4743 215904 4752
rect 215852 4709 215861 4743
rect 215861 4709 215895 4743
rect 215895 4709 215904 4743
rect 215852 4700 215904 4709
rect 217416 4743 217468 4752
rect 217416 4709 217425 4743
rect 217425 4709 217459 4743
rect 217459 4709 217468 4743
rect 217416 4700 217468 4709
rect 213276 4632 213328 4684
rect 216404 4675 216456 4684
rect 216404 4641 216413 4675
rect 216413 4641 216447 4675
rect 216447 4641 216456 4675
rect 216404 4632 216456 4641
rect 220636 4675 220688 4684
rect 220636 4641 220645 4675
rect 220645 4641 220679 4675
rect 220679 4641 220688 4675
rect 220636 4632 220688 4641
rect 222016 4700 222068 4752
rect 228272 4700 228324 4752
rect 229744 4768 229796 4820
rect 237196 4768 237248 4820
rect 237288 4768 237340 4820
rect 230756 4743 230808 4752
rect 230756 4709 230765 4743
rect 230765 4709 230799 4743
rect 230799 4709 230808 4743
rect 230756 4700 230808 4709
rect 240324 4811 240376 4820
rect 240324 4777 240333 4811
rect 240333 4777 240367 4811
rect 240367 4777 240376 4811
rect 240324 4768 240376 4777
rect 240968 4768 241020 4820
rect 242624 4768 242676 4820
rect 244280 4768 244332 4820
rect 252468 4768 252520 4820
rect 253572 4811 253624 4820
rect 253572 4777 253581 4811
rect 253581 4777 253615 4811
rect 253615 4777 253624 4811
rect 253572 4768 253624 4777
rect 157892 4564 157944 4616
rect 158076 4496 158128 4548
rect 158536 4539 158588 4548
rect 158536 4505 158545 4539
rect 158545 4505 158579 4539
rect 158579 4505 158588 4539
rect 158536 4496 158588 4505
rect 160836 4539 160888 4548
rect 142436 4428 142488 4437
rect 148968 4428 149020 4480
rect 151820 4428 151872 4480
rect 155224 4428 155276 4480
rect 156328 4428 156380 4480
rect 158168 4471 158220 4480
rect 158168 4437 158177 4471
rect 158177 4437 158211 4471
rect 158211 4437 158220 4471
rect 160836 4505 160845 4539
rect 160845 4505 160879 4539
rect 160879 4505 160888 4539
rect 160836 4496 160888 4505
rect 161020 4607 161072 4616
rect 161020 4573 161029 4607
rect 161029 4573 161063 4607
rect 161063 4573 161072 4607
rect 161020 4564 161072 4573
rect 161204 4539 161256 4548
rect 161204 4505 161213 4539
rect 161213 4505 161247 4539
rect 161247 4505 161256 4539
rect 161204 4496 161256 4505
rect 161388 4496 161440 4548
rect 163136 4539 163188 4548
rect 163136 4505 163145 4539
rect 163145 4505 163179 4539
rect 163179 4505 163188 4539
rect 163136 4496 163188 4505
rect 158168 4428 158220 4437
rect 162032 4428 162084 4480
rect 213920 4564 213972 4616
rect 214104 4496 214156 4548
rect 214564 4564 214616 4616
rect 216128 4607 216180 4616
rect 216128 4573 216137 4607
rect 216137 4573 216171 4607
rect 216171 4573 216180 4607
rect 216128 4564 216180 4573
rect 216312 4564 216364 4616
rect 222476 4607 222528 4616
rect 222476 4573 222485 4607
rect 222485 4573 222519 4607
rect 222519 4573 222528 4607
rect 222476 4564 222528 4573
rect 226156 4564 226208 4616
rect 228824 4607 228876 4616
rect 228824 4573 228833 4607
rect 228833 4573 228867 4607
rect 228867 4573 228876 4607
rect 228824 4564 228876 4573
rect 231216 4607 231268 4616
rect 231216 4573 231225 4607
rect 231225 4573 231259 4607
rect 231259 4573 231268 4607
rect 231216 4564 231268 4573
rect 231492 4564 231544 4616
rect 246488 4700 246540 4752
rect 239220 4607 239272 4616
rect 239220 4573 239229 4607
rect 239229 4573 239263 4607
rect 239263 4573 239272 4607
rect 239220 4564 239272 4573
rect 240968 4607 241020 4616
rect 240968 4573 240977 4607
rect 240977 4573 241011 4607
rect 241011 4573 241020 4607
rect 240968 4564 241020 4573
rect 242256 4607 242308 4616
rect 242256 4573 242265 4607
rect 242265 4573 242299 4607
rect 242299 4573 242308 4607
rect 242256 4564 242308 4573
rect 250628 4675 250680 4684
rect 250628 4641 250637 4675
rect 250637 4641 250671 4675
rect 250671 4641 250680 4675
rect 250628 4632 250680 4641
rect 255780 4811 255832 4820
rect 255780 4777 255789 4811
rect 255789 4777 255823 4811
rect 255823 4777 255832 4811
rect 256700 4811 256752 4820
rect 255780 4768 255832 4777
rect 256700 4777 256709 4811
rect 256709 4777 256743 4811
rect 256743 4777 256752 4811
rect 256700 4768 256752 4777
rect 259460 4768 259512 4820
rect 263048 4811 263100 4820
rect 263048 4777 263057 4811
rect 263057 4777 263091 4811
rect 263091 4777 263100 4811
rect 263048 4768 263100 4777
rect 265164 4811 265216 4820
rect 265164 4777 265173 4811
rect 265173 4777 265207 4811
rect 265207 4777 265216 4811
rect 265164 4768 265216 4777
rect 266912 4811 266964 4820
rect 266912 4777 266921 4811
rect 266921 4777 266955 4811
rect 266955 4777 266964 4811
rect 266912 4768 266964 4777
rect 268568 4768 268620 4820
rect 270960 4768 271012 4820
rect 255320 4700 255372 4752
rect 259276 4743 259328 4752
rect 259276 4709 259285 4743
rect 259285 4709 259319 4743
rect 259319 4709 259328 4743
rect 259276 4700 259328 4709
rect 264060 4700 264112 4752
rect 264244 4700 264296 4752
rect 215116 4428 215168 4480
rect 220176 4496 220228 4548
rect 222016 4496 222068 4548
rect 223672 4496 223724 4548
rect 218888 4428 218940 4480
rect 226248 4539 226300 4548
rect 226248 4505 226257 4539
rect 226257 4505 226291 4539
rect 226291 4505 226300 4539
rect 226248 4496 226300 4505
rect 226800 4496 226852 4548
rect 228732 4539 228784 4548
rect 228732 4505 228741 4539
rect 228741 4505 228775 4539
rect 228775 4505 228784 4539
rect 228732 4496 228784 4505
rect 226616 4428 226668 4480
rect 228272 4428 228324 4480
rect 230756 4539 230808 4548
rect 230756 4505 230765 4539
rect 230765 4505 230799 4539
rect 230799 4505 230808 4539
rect 230756 4496 230808 4505
rect 230296 4428 230348 4480
rect 251364 4564 251416 4616
rect 251456 4607 251508 4616
rect 251456 4573 251465 4607
rect 251465 4573 251499 4607
rect 251499 4573 251508 4607
rect 251456 4564 251508 4573
rect 255044 4607 255096 4616
rect 255044 4573 255053 4607
rect 255053 4573 255087 4607
rect 255087 4573 255096 4607
rect 255044 4564 255096 4573
rect 231492 4471 231544 4480
rect 231492 4437 231501 4471
rect 231501 4437 231535 4471
rect 231535 4437 231544 4471
rect 231492 4428 231544 4437
rect 239680 4471 239732 4480
rect 239680 4437 239689 4471
rect 239689 4437 239723 4471
rect 239723 4437 239732 4471
rect 239680 4428 239732 4437
rect 241612 4471 241664 4480
rect 241612 4437 241621 4471
rect 241621 4437 241655 4471
rect 241655 4437 241664 4471
rect 241612 4428 241664 4437
rect 243268 4471 243320 4480
rect 243268 4437 243277 4471
rect 243277 4437 243311 4471
rect 243311 4437 243320 4471
rect 243268 4428 243320 4437
rect 245384 4471 245436 4480
rect 245384 4437 245393 4471
rect 245393 4437 245427 4471
rect 245427 4437 245436 4471
rect 245384 4428 245436 4437
rect 251916 4471 251968 4480
rect 251916 4437 251925 4471
rect 251925 4437 251959 4471
rect 251959 4437 251968 4471
rect 251916 4428 251968 4437
rect 254032 4496 254084 4548
rect 256700 4564 256752 4616
rect 255320 4539 255372 4548
rect 255320 4505 255329 4539
rect 255329 4505 255363 4539
rect 255363 4505 255372 4539
rect 255320 4496 255372 4505
rect 258172 4607 258224 4616
rect 258172 4573 258181 4607
rect 258181 4573 258215 4607
rect 258215 4573 258224 4607
rect 258172 4564 258224 4573
rect 257804 4496 257856 4548
rect 263324 4564 263376 4616
rect 266268 4632 266320 4684
rect 267740 4632 267792 4684
rect 259736 4496 259788 4548
rect 260104 4496 260156 4548
rect 264152 4539 264204 4548
rect 264152 4505 264161 4539
rect 264161 4505 264195 4539
rect 264195 4505 264204 4539
rect 264152 4496 264204 4505
rect 265808 4607 265860 4616
rect 265808 4573 265817 4607
rect 265817 4573 265851 4607
rect 265851 4573 265860 4607
rect 265808 4564 265860 4573
rect 265900 4564 265952 4616
rect 266084 4564 266136 4616
rect 267372 4564 267424 4616
rect 267556 4564 267608 4616
rect 268200 4607 268252 4616
rect 268200 4573 268209 4607
rect 268209 4573 268243 4607
rect 268243 4573 268252 4607
rect 268200 4564 268252 4573
rect 269120 4564 269172 4616
rect 269764 4564 269816 4616
rect 271144 4564 271196 4616
rect 272156 4564 272208 4616
rect 268476 4496 268528 4548
rect 268568 4539 268620 4548
rect 268568 4505 268577 4539
rect 268577 4505 268611 4539
rect 268611 4505 268620 4539
rect 268568 4496 268620 4505
rect 256700 4428 256752 4480
rect 257712 4471 257764 4480
rect 257712 4437 257721 4471
rect 257721 4437 257755 4471
rect 257755 4437 257764 4471
rect 257712 4428 257764 4437
rect 260288 4471 260340 4480
rect 260288 4437 260297 4471
rect 260297 4437 260331 4471
rect 260331 4437 260340 4471
rect 260288 4428 260340 4437
rect 270224 4496 270276 4548
rect 68546 4326 68598 4378
rect 68610 4326 68662 4378
rect 68674 4326 68726 4378
rect 68738 4326 68790 4378
rect 68802 4326 68854 4378
rect 136143 4326 136195 4378
rect 136207 4326 136259 4378
rect 136271 4326 136323 4378
rect 136335 4326 136387 4378
rect 136399 4326 136451 4378
rect 203740 4326 203792 4378
rect 203804 4326 203856 4378
rect 203868 4326 203920 4378
rect 203932 4326 203984 4378
rect 203996 4326 204048 4378
rect 271337 4326 271389 4378
rect 271401 4326 271453 4378
rect 271465 4326 271517 4378
rect 271529 4326 271581 4378
rect 271593 4326 271645 4378
rect 23296 4224 23348 4276
rect 23572 4088 23624 4140
rect 25780 4131 25832 4140
rect 25780 4097 25789 4131
rect 25789 4097 25823 4131
rect 25823 4097 25832 4131
rect 25780 4088 25832 4097
rect 40224 4156 40276 4208
rect 38936 4088 38988 4140
rect 40592 4199 40644 4208
rect 40592 4165 40601 4199
rect 40601 4165 40635 4199
rect 40635 4165 40644 4199
rect 40592 4156 40644 4165
rect 41236 4156 41288 4208
rect 42892 4224 42944 4276
rect 48596 4224 48648 4276
rect 49056 4224 49108 4276
rect 51172 4224 51224 4276
rect 53380 4224 53432 4276
rect 40868 4131 40920 4140
rect 40868 4097 40877 4131
rect 40877 4097 40911 4131
rect 40911 4097 40920 4131
rect 40868 4088 40920 4097
rect 41052 4088 41104 4140
rect 42616 4156 42668 4208
rect 48044 4156 48096 4208
rect 49148 4156 49200 4208
rect 49240 4199 49292 4208
rect 49240 4165 49249 4199
rect 49249 4165 49283 4199
rect 49283 4165 49292 4199
rect 49240 4156 49292 4165
rect 49332 4199 49384 4208
rect 49332 4165 49341 4199
rect 49341 4165 49375 4199
rect 49375 4165 49384 4199
rect 49332 4156 49384 4165
rect 49884 4156 49936 4208
rect 51540 4156 51592 4208
rect 51724 4199 51776 4208
rect 51724 4165 51733 4199
rect 51733 4165 51767 4199
rect 51767 4165 51776 4199
rect 51724 4156 51776 4165
rect 51816 4156 51868 4208
rect 80888 4156 80940 4208
rect 81624 4199 81676 4208
rect 81624 4165 81633 4199
rect 81633 4165 81667 4199
rect 81667 4165 81676 4199
rect 81624 4156 81676 4165
rect 83648 4156 83700 4208
rect 51264 4131 51316 4140
rect 51264 4097 51273 4131
rect 51273 4097 51307 4131
rect 51307 4097 51316 4131
rect 51264 4088 51316 4097
rect 51356 4131 51408 4140
rect 51356 4097 51365 4131
rect 51365 4097 51399 4131
rect 51399 4097 51408 4131
rect 51356 4088 51408 4097
rect 52460 4088 52512 4140
rect 87512 4224 87564 4276
rect 112996 4224 113048 4276
rect 113180 4224 113232 4276
rect 123392 4224 123444 4276
rect 84936 4199 84988 4208
rect 84936 4165 84945 4199
rect 84945 4165 84979 4199
rect 84979 4165 84988 4199
rect 84936 4156 84988 4165
rect 96068 4156 96120 4208
rect 102048 4156 102100 4208
rect 109868 4156 109920 4208
rect 112536 4156 112588 4208
rect 116400 4156 116452 4208
rect 14372 4020 14424 4072
rect 9220 3952 9272 4004
rect 36544 3952 36596 4004
rect 24492 3884 24544 3936
rect 40776 4020 40828 4072
rect 49792 4020 49844 4072
rect 51632 4020 51684 4072
rect 81440 4063 81492 4072
rect 81440 4029 81449 4063
rect 81449 4029 81483 4063
rect 81483 4029 81492 4063
rect 81440 4020 81492 4029
rect 91008 4088 91060 4140
rect 94320 4131 94372 4140
rect 94320 4097 94329 4131
rect 94329 4097 94363 4131
rect 94363 4097 94372 4131
rect 94320 4088 94372 4097
rect 104992 4088 105044 4140
rect 105820 4131 105872 4140
rect 105820 4097 105829 4131
rect 105829 4097 105863 4131
rect 105863 4097 105872 4131
rect 105820 4088 105872 4097
rect 106740 4088 106792 4140
rect 108396 4131 108448 4140
rect 108396 4097 108405 4131
rect 108405 4097 108439 4131
rect 108439 4097 108448 4131
rect 108396 4088 108448 4097
rect 112352 4131 112404 4140
rect 112352 4097 112361 4131
rect 112361 4097 112395 4131
rect 112395 4097 112404 4131
rect 112352 4088 112404 4097
rect 113548 4131 113600 4140
rect 113548 4097 113557 4131
rect 113557 4097 113591 4131
rect 113591 4097 113600 4131
rect 113548 4088 113600 4097
rect 114192 4131 114244 4140
rect 114192 4097 114201 4131
rect 114201 4097 114235 4131
rect 114235 4097 114244 4131
rect 114192 4088 114244 4097
rect 114744 4088 114796 4140
rect 115572 4131 115624 4140
rect 115572 4097 115581 4131
rect 115581 4097 115615 4131
rect 115615 4097 115624 4131
rect 115572 4088 115624 4097
rect 142436 4224 142488 4276
rect 151084 4224 151136 4276
rect 154396 4224 154448 4276
rect 123668 4156 123720 4208
rect 147496 4199 147548 4208
rect 147496 4165 147505 4199
rect 147505 4165 147539 4199
rect 147539 4165 147548 4199
rect 147496 4156 147548 4165
rect 148416 4156 148468 4208
rect 148876 4156 148928 4208
rect 151820 4156 151872 4208
rect 154672 4156 154724 4208
rect 213920 4224 213972 4276
rect 215116 4224 215168 4276
rect 219072 4224 219124 4276
rect 222016 4224 222068 4276
rect 157800 4199 157852 4208
rect 157800 4165 157809 4199
rect 157809 4165 157843 4199
rect 157843 4165 157852 4199
rect 157800 4156 157852 4165
rect 161296 4199 161348 4208
rect 161296 4165 161305 4199
rect 161305 4165 161339 4199
rect 161339 4165 161348 4199
rect 161296 4156 161348 4165
rect 190000 4199 190052 4208
rect 190000 4165 190009 4199
rect 190009 4165 190043 4199
rect 190043 4165 190052 4199
rect 190000 4156 190052 4165
rect 209688 4156 209740 4208
rect 93768 4020 93820 4072
rect 96160 4063 96212 4072
rect 96160 4029 96169 4063
rect 96169 4029 96203 4063
rect 96203 4029 96212 4063
rect 96160 4020 96212 4029
rect 98552 4020 98604 4072
rect 99748 4020 99800 4072
rect 92296 3952 92348 4004
rect 98920 3952 98972 4004
rect 40408 3884 40460 3936
rect 41880 3927 41932 3936
rect 41880 3893 41889 3927
rect 41889 3893 41923 3927
rect 41923 3893 41932 3927
rect 41880 3884 41932 3893
rect 42800 3884 42852 3936
rect 47400 3884 47452 3936
rect 52276 3927 52328 3936
rect 52276 3893 52285 3927
rect 52285 3893 52319 3927
rect 52319 3893 52328 3927
rect 52276 3884 52328 3893
rect 83924 3927 83976 3936
rect 83924 3893 83933 3927
rect 83933 3893 83967 3927
rect 83967 3893 83976 3927
rect 83924 3884 83976 3893
rect 87696 3884 87748 3936
rect 96896 3884 96948 3936
rect 98184 3884 98236 3936
rect 102232 4020 102284 4072
rect 102876 3952 102928 4004
rect 105084 4063 105136 4072
rect 105084 4029 105093 4063
rect 105093 4029 105127 4063
rect 105127 4029 105136 4063
rect 105084 4020 105136 4029
rect 105544 4063 105596 4072
rect 105544 4029 105553 4063
rect 105553 4029 105587 4063
rect 105587 4029 105596 4063
rect 105544 4020 105596 4029
rect 106004 4020 106056 4072
rect 101588 3927 101640 3936
rect 101588 3893 101597 3927
rect 101597 3893 101631 3927
rect 101631 3893 101640 3927
rect 101588 3884 101640 3893
rect 104532 3927 104584 3936
rect 104532 3893 104541 3927
rect 104541 3893 104575 3927
rect 104575 3893 104584 3927
rect 104532 3884 104584 3893
rect 107292 4020 107344 4072
rect 107384 4063 107436 4072
rect 107384 4029 107393 4063
rect 107393 4029 107427 4063
rect 107427 4029 107436 4063
rect 107384 4020 107436 4029
rect 106924 3952 106976 4004
rect 107752 3952 107804 4004
rect 107108 3884 107160 3936
rect 111340 4020 111392 4072
rect 112536 4063 112588 4072
rect 112536 4029 112545 4063
rect 112545 4029 112579 4063
rect 112579 4029 112588 4063
rect 112536 4020 112588 4029
rect 112444 3952 112496 4004
rect 112996 3995 113048 4004
rect 112996 3961 113005 3995
rect 113005 3961 113039 3995
rect 113039 3961 113048 3995
rect 112996 3952 113048 3961
rect 108948 3884 109000 3936
rect 110236 3884 110288 3936
rect 113456 4020 113508 4072
rect 114836 4063 114888 4072
rect 114836 4029 114845 4063
rect 114845 4029 114879 4063
rect 114879 4029 114888 4063
rect 114836 4020 114888 4029
rect 115296 3995 115348 4004
rect 115296 3961 115305 3995
rect 115305 3961 115339 3995
rect 115339 3961 115348 3995
rect 115296 3952 115348 3961
rect 114560 3884 114612 3936
rect 116032 4020 116084 4072
rect 116768 4020 116820 4072
rect 117688 4063 117740 4072
rect 117688 4029 117697 4063
rect 117697 4029 117731 4063
rect 117731 4029 117740 4063
rect 117688 4020 117740 4029
rect 121000 4020 121052 4072
rect 121920 4063 121972 4072
rect 121920 4029 121929 4063
rect 121929 4029 121963 4063
rect 121963 4029 121972 4063
rect 121920 4020 121972 4029
rect 122656 4020 122708 4072
rect 116400 3884 116452 3936
rect 116492 3927 116544 3936
rect 116492 3893 116501 3927
rect 116501 3893 116535 3927
rect 116535 3893 116544 3927
rect 116492 3884 116544 3893
rect 116676 3884 116728 3936
rect 120908 3952 120960 4004
rect 119988 3927 120040 3936
rect 119988 3893 119997 3927
rect 119997 3893 120031 3927
rect 120031 3893 120040 3927
rect 119988 3884 120040 3893
rect 124312 4020 124364 4072
rect 139308 4020 139360 4072
rect 141792 4063 141844 4072
rect 141792 4029 141801 4063
rect 141801 4029 141835 4063
rect 141835 4029 141844 4063
rect 141792 4020 141844 4029
rect 142160 4020 142212 4072
rect 145656 4063 145708 4072
rect 145656 4029 145665 4063
rect 145665 4029 145699 4063
rect 145699 4029 145708 4063
rect 145656 4020 145708 4029
rect 150900 4088 150952 4140
rect 152648 4131 152700 4140
rect 152648 4097 152657 4131
rect 152657 4097 152691 4131
rect 152691 4097 152700 4131
rect 152648 4088 152700 4097
rect 154488 4088 154540 4140
rect 147956 4063 148008 4072
rect 147956 4029 147965 4063
rect 147965 4029 147999 4063
rect 147999 4029 148008 4063
rect 147956 4020 148008 4029
rect 148140 4063 148192 4072
rect 148140 4029 148149 4063
rect 148149 4029 148183 4063
rect 148183 4029 148192 4063
rect 148140 4020 148192 4029
rect 149060 4020 149112 4072
rect 149796 4063 149848 4072
rect 149796 4029 149805 4063
rect 149805 4029 149839 4063
rect 149839 4029 149848 4063
rect 149796 4020 149848 4029
rect 151268 4020 151320 4072
rect 152464 4020 152516 4072
rect 152832 4020 152884 4072
rect 152924 4063 152976 4072
rect 152924 4029 152933 4063
rect 152933 4029 152967 4063
rect 152967 4029 152976 4063
rect 152924 4020 152976 4029
rect 155684 4088 155736 4140
rect 154856 4063 154908 4072
rect 154856 4029 154865 4063
rect 154865 4029 154899 4063
rect 154899 4029 154908 4063
rect 156328 4088 156380 4140
rect 154856 4020 154908 4029
rect 156236 4020 156288 4072
rect 159180 4131 159232 4140
rect 159180 4097 159189 4131
rect 159189 4097 159223 4131
rect 159223 4097 159232 4131
rect 159180 4088 159232 4097
rect 159456 4131 159508 4140
rect 159456 4097 159465 4131
rect 159465 4097 159499 4131
rect 159499 4097 159508 4131
rect 159456 4088 159508 4097
rect 157708 4020 157760 4072
rect 158628 4020 158680 4072
rect 160744 4088 160796 4140
rect 162492 4088 162544 4140
rect 161388 4020 161440 4072
rect 163688 4063 163740 4072
rect 163688 4029 163697 4063
rect 163697 4029 163731 4063
rect 163731 4029 163740 4063
rect 163688 4020 163740 4029
rect 190920 4088 190972 4140
rect 209320 4131 209372 4140
rect 209320 4097 209329 4131
rect 209329 4097 209363 4131
rect 209363 4097 209372 4131
rect 209320 4088 209372 4097
rect 216864 4156 216916 4208
rect 212632 4088 212684 4140
rect 214012 4131 214064 4140
rect 214012 4097 214021 4131
rect 214021 4097 214055 4131
rect 214055 4097 214064 4131
rect 214012 4088 214064 4097
rect 214932 4131 214984 4140
rect 214932 4097 214941 4131
rect 214941 4097 214975 4131
rect 214975 4097 214984 4131
rect 214932 4088 214984 4097
rect 215852 4131 215904 4140
rect 215852 4097 215861 4131
rect 215861 4097 215895 4131
rect 215895 4097 215904 4131
rect 215852 4088 215904 4097
rect 216128 4131 216180 4140
rect 216128 4097 216137 4131
rect 216137 4097 216171 4131
rect 216171 4097 216180 4131
rect 216128 4088 216180 4097
rect 240048 4224 240100 4276
rect 226616 4156 226668 4208
rect 231032 4156 231084 4208
rect 235632 4199 235684 4208
rect 235632 4165 235641 4199
rect 235641 4165 235675 4199
rect 235675 4165 235684 4199
rect 235632 4156 235684 4165
rect 239680 4156 239732 4208
rect 207480 4063 207532 4072
rect 207480 4029 207489 4063
rect 207489 4029 207523 4063
rect 207523 4029 207532 4063
rect 207480 4020 207532 4029
rect 207756 4020 207808 4072
rect 209964 4063 210016 4072
rect 209964 4029 209973 4063
rect 209973 4029 210007 4063
rect 210007 4029 210016 4063
rect 209964 4020 210016 4029
rect 124036 3884 124088 3936
rect 141424 3927 141476 3936
rect 141424 3893 141433 3927
rect 141433 3893 141467 3927
rect 141467 3893 141476 3927
rect 141424 3884 141476 3893
rect 147496 3884 147548 3936
rect 150992 3884 151044 3936
rect 156972 3884 157024 3936
rect 160468 3884 160520 3936
rect 161388 3884 161440 3936
rect 207664 3884 207716 3936
rect 208032 3952 208084 4004
rect 211804 4020 211856 4072
rect 213092 4020 213144 4072
rect 213460 4063 213512 4072
rect 213460 4029 213469 4063
rect 213469 4029 213503 4063
rect 213503 4029 213512 4063
rect 213460 4020 213512 4029
rect 209320 3884 209372 3936
rect 210884 3884 210936 3936
rect 213276 3884 213328 3936
rect 213828 4063 213880 4072
rect 213828 4029 213862 4063
rect 213862 4029 213880 4063
rect 213828 4020 213880 4029
rect 214196 4020 214248 4072
rect 215484 4020 215536 4072
rect 221648 4020 221700 4072
rect 222936 4020 222988 4072
rect 224500 4063 224552 4072
rect 224500 4029 224509 4063
rect 224509 4029 224543 4063
rect 224543 4029 224552 4063
rect 224500 4020 224552 4029
rect 226156 4131 226208 4140
rect 226156 4097 226165 4131
rect 226165 4097 226199 4131
rect 226199 4097 226208 4131
rect 226156 4088 226208 4097
rect 229836 4088 229888 4140
rect 231308 4088 231360 4140
rect 236920 4088 236972 4140
rect 242992 4224 243044 4276
rect 245384 4224 245436 4276
rect 264888 4224 264940 4276
rect 265808 4224 265860 4276
rect 266176 4224 266228 4276
rect 268108 4224 268160 4276
rect 268200 4224 268252 4276
rect 241612 4156 241664 4208
rect 243268 4156 243320 4208
rect 251364 4156 251416 4208
rect 254032 4199 254084 4208
rect 254032 4165 254041 4199
rect 254041 4165 254075 4199
rect 254075 4165 254084 4199
rect 254032 4156 254084 4165
rect 255320 4156 255372 4208
rect 257712 4156 257764 4208
rect 260196 4199 260248 4208
rect 260196 4165 260205 4199
rect 260205 4165 260239 4199
rect 260239 4165 260248 4199
rect 260196 4156 260248 4165
rect 260288 4156 260340 4208
rect 240784 4131 240836 4140
rect 240784 4097 240793 4131
rect 240793 4097 240827 4131
rect 240827 4097 240836 4131
rect 240784 4088 240836 4097
rect 260012 4088 260064 4140
rect 264980 4156 265032 4208
rect 268844 4156 268896 4208
rect 265900 4131 265952 4140
rect 265900 4097 265909 4131
rect 265909 4097 265943 4131
rect 265943 4097 265952 4131
rect 265900 4088 265952 4097
rect 267096 4088 267148 4140
rect 267188 4131 267240 4140
rect 267188 4097 267197 4131
rect 267197 4097 267231 4131
rect 267231 4097 267240 4131
rect 267188 4088 267240 4097
rect 267648 4131 267700 4140
rect 267648 4097 267657 4131
rect 267657 4097 267691 4131
rect 267691 4097 267700 4131
rect 267648 4088 267700 4097
rect 268660 4088 268712 4140
rect 271696 4156 271748 4208
rect 269672 4088 269724 4140
rect 270684 4088 270736 4140
rect 225236 4063 225288 4072
rect 225236 4029 225245 4063
rect 225245 4029 225279 4063
rect 225279 4029 225288 4063
rect 225236 4020 225288 4029
rect 225328 4063 225380 4072
rect 225328 4029 225362 4063
rect 225362 4029 225380 4063
rect 225328 4020 225380 4029
rect 214656 3927 214708 3936
rect 214656 3893 214665 3927
rect 214665 3893 214699 3927
rect 214699 3893 214708 3927
rect 214656 3884 214708 3893
rect 216588 3884 216640 3936
rect 218152 3884 218204 3936
rect 224960 3995 225012 4004
rect 224960 3961 224969 3995
rect 224969 3961 225003 3995
rect 225003 3961 225012 3995
rect 224960 3952 225012 3961
rect 226064 4020 226116 4072
rect 226984 4020 227036 4072
rect 227352 4020 227404 4072
rect 228272 4063 228324 4072
rect 228272 4029 228281 4063
rect 228281 4029 228315 4063
rect 228315 4029 228324 4063
rect 228272 4020 228324 4029
rect 229100 4063 229152 4072
rect 229100 4029 229109 4063
rect 229109 4029 229143 4063
rect 229143 4029 229152 4063
rect 229100 4020 229152 4029
rect 230296 4020 230348 4072
rect 226616 3952 226668 4004
rect 230480 3952 230532 4004
rect 230756 4020 230808 4072
rect 237380 4020 237432 4072
rect 251456 4020 251508 4072
rect 230664 3952 230716 4004
rect 226800 3927 226852 3936
rect 226800 3893 226809 3927
rect 226809 3893 226843 3927
rect 226843 3893 226852 3927
rect 226800 3884 226852 3893
rect 226892 3884 226944 3936
rect 227444 3927 227496 3936
rect 227444 3893 227453 3927
rect 227453 3893 227487 3927
rect 227487 3893 227496 3927
rect 227444 3884 227496 3893
rect 231032 3884 231084 3936
rect 235540 3884 235592 3936
rect 243176 3952 243228 4004
rect 244188 3995 244240 4004
rect 244188 3961 244197 3995
rect 244197 3961 244231 3995
rect 244231 3961 244240 3995
rect 244188 3952 244240 3961
rect 242440 3884 242492 3936
rect 242532 3927 242584 3936
rect 242532 3893 242541 3927
rect 242541 3893 242575 3927
rect 242575 3893 242584 3927
rect 242532 3884 242584 3893
rect 242808 3884 242860 3936
rect 253940 4063 253992 4072
rect 253940 4029 253949 4063
rect 253949 4029 253983 4063
rect 253983 4029 253992 4063
rect 253940 4020 253992 4029
rect 256516 4063 256568 4072
rect 256516 4029 256525 4063
rect 256525 4029 256559 4063
rect 256559 4029 256568 4063
rect 256516 4020 256568 4029
rect 256700 4063 256752 4072
rect 256700 4029 256709 4063
rect 256709 4029 256743 4063
rect 256743 4029 256752 4063
rect 256700 4020 256752 4029
rect 257620 4063 257672 4072
rect 257620 4029 257629 4063
rect 257629 4029 257663 4063
rect 257663 4029 257672 4063
rect 257620 4020 257672 4029
rect 257804 4063 257856 4072
rect 257804 4029 257813 4063
rect 257813 4029 257847 4063
rect 257847 4029 257856 4063
rect 257804 4020 257856 4029
rect 258172 4020 258224 4072
rect 265624 4020 265676 4072
rect 260104 3952 260156 4004
rect 258080 3884 258132 3936
rect 258264 3927 258316 3936
rect 258264 3893 258273 3927
rect 258273 3893 258307 3927
rect 258307 3893 258316 3927
rect 258264 3884 258316 3893
rect 258540 3927 258592 3936
rect 258540 3893 258549 3927
rect 258549 3893 258583 3927
rect 258583 3893 258592 3927
rect 258540 3884 258592 3893
rect 259920 3927 259972 3936
rect 259920 3893 259929 3927
rect 259929 3893 259963 3927
rect 259963 3893 259972 3927
rect 259920 3884 259972 3893
rect 264796 3884 264848 3936
rect 266360 3927 266412 3936
rect 266360 3893 266369 3927
rect 266369 3893 266403 3927
rect 266403 3893 266412 3927
rect 266360 3884 266412 3893
rect 267004 3995 267056 4004
rect 267004 3961 267013 3995
rect 267013 3961 267047 3995
rect 267047 3961 267056 3995
rect 267004 3952 267056 3961
rect 267924 3952 267976 4004
rect 268384 4063 268436 4072
rect 268384 4029 268393 4063
rect 268393 4029 268427 4063
rect 268427 4029 268436 4063
rect 268384 4020 268436 4029
rect 268844 4020 268896 4072
rect 270868 4131 270920 4140
rect 270868 4097 270877 4131
rect 270877 4097 270911 4131
rect 270911 4097 270920 4131
rect 270868 4088 270920 4097
rect 269028 3884 269080 3936
rect 269396 3884 269448 3936
rect 270500 3884 270552 3936
rect 34748 3782 34800 3834
rect 34812 3782 34864 3834
rect 34876 3782 34928 3834
rect 34940 3782 34992 3834
rect 35004 3782 35056 3834
rect 102345 3782 102397 3834
rect 102409 3782 102461 3834
rect 102473 3782 102525 3834
rect 102537 3782 102589 3834
rect 102601 3782 102653 3834
rect 169942 3782 169994 3834
rect 170006 3782 170058 3834
rect 170070 3782 170122 3834
rect 170134 3782 170186 3834
rect 170198 3782 170250 3834
rect 237539 3782 237591 3834
rect 237603 3782 237655 3834
rect 237667 3782 237719 3834
rect 237731 3782 237783 3834
rect 237795 3782 237847 3834
rect 3332 3680 3384 3732
rect 36452 3680 36504 3732
rect 39948 3680 40000 3732
rect 66720 3680 66772 3732
rect 79232 3680 79284 3732
rect 84016 3680 84068 3732
rect 87512 3680 87564 3732
rect 40040 3612 40092 3664
rect 40776 3612 40828 3664
rect 15108 3544 15160 3596
rect 19340 3544 19392 3596
rect 24952 3587 25004 3596
rect 24952 3553 24961 3587
rect 24961 3553 24995 3587
rect 24995 3553 25004 3587
rect 24952 3544 25004 3553
rect 25044 3476 25096 3528
rect 25412 3476 25464 3528
rect 26240 3476 26292 3528
rect 26516 3519 26568 3528
rect 26516 3485 26525 3519
rect 26525 3485 26559 3519
rect 26559 3485 26568 3519
rect 26516 3476 26568 3485
rect 27528 3476 27580 3528
rect 36636 3476 36688 3528
rect 37280 3476 37332 3528
rect 11152 3408 11204 3460
rect 20720 3408 20772 3460
rect 22744 3408 22796 3460
rect 27620 3408 27672 3460
rect 37556 3544 37608 3596
rect 48044 3544 48096 3596
rect 38476 3408 38528 3460
rect 40960 3408 41012 3460
rect 23756 3340 23808 3392
rect 25964 3383 26016 3392
rect 25964 3349 25973 3383
rect 25973 3349 26007 3383
rect 26007 3349 26016 3383
rect 25964 3340 26016 3349
rect 26700 3383 26752 3392
rect 26700 3349 26709 3383
rect 26709 3349 26743 3383
rect 26743 3349 26752 3383
rect 26700 3340 26752 3349
rect 27436 3383 27488 3392
rect 27436 3349 27445 3383
rect 27445 3349 27479 3383
rect 27479 3349 27488 3383
rect 27436 3340 27488 3349
rect 35900 3383 35952 3392
rect 35900 3349 35909 3383
rect 35909 3349 35943 3383
rect 35943 3349 35952 3383
rect 35900 3340 35952 3349
rect 36084 3340 36136 3392
rect 37556 3383 37608 3392
rect 37556 3349 37565 3383
rect 37565 3349 37599 3383
rect 37599 3349 37608 3383
rect 37556 3340 37608 3349
rect 38660 3340 38712 3392
rect 40408 3340 40460 3392
rect 41236 3383 41288 3392
rect 41236 3349 41245 3383
rect 41245 3349 41279 3383
rect 41279 3349 41288 3383
rect 41236 3340 41288 3349
rect 41512 3451 41564 3460
rect 41512 3417 41521 3451
rect 41521 3417 41555 3451
rect 41555 3417 41564 3451
rect 41512 3408 41564 3417
rect 41604 3451 41656 3460
rect 41604 3417 41613 3451
rect 41613 3417 41647 3451
rect 41647 3417 41656 3451
rect 41604 3408 41656 3417
rect 41972 3451 42024 3460
rect 41972 3417 41981 3451
rect 41981 3417 42015 3451
rect 42015 3417 42024 3451
rect 41972 3408 42024 3417
rect 46664 3451 46716 3460
rect 46664 3417 46673 3451
rect 46673 3417 46707 3451
rect 46707 3417 46716 3451
rect 46664 3408 46716 3417
rect 46940 3451 46992 3460
rect 46940 3417 46949 3451
rect 46949 3417 46983 3451
rect 46983 3417 46992 3451
rect 46940 3408 46992 3417
rect 47216 3408 47268 3460
rect 47400 3451 47452 3460
rect 47400 3417 47409 3451
rect 47409 3417 47443 3451
rect 47443 3417 47452 3451
rect 47400 3408 47452 3417
rect 60740 3612 60792 3664
rect 94228 3612 94280 3664
rect 51908 3476 51960 3528
rect 66996 3476 67048 3528
rect 77300 3544 77352 3596
rect 67180 3476 67232 3528
rect 79232 3408 79284 3460
rect 83648 3451 83700 3460
rect 83648 3417 83657 3451
rect 83657 3417 83691 3451
rect 83691 3417 83700 3451
rect 83648 3408 83700 3417
rect 84476 3408 84528 3460
rect 84936 3408 84988 3460
rect 85396 3408 85448 3460
rect 88248 3476 88300 3528
rect 85672 3383 85724 3392
rect 85672 3349 85681 3383
rect 85681 3349 85715 3383
rect 85715 3349 85724 3383
rect 85672 3340 85724 3349
rect 86040 3340 86092 3392
rect 95884 3519 95936 3528
rect 95884 3485 95893 3519
rect 95893 3485 95927 3519
rect 95927 3485 95936 3519
rect 95884 3476 95936 3485
rect 91652 3408 91704 3460
rect 91928 3451 91980 3460
rect 91928 3417 91937 3451
rect 91937 3417 91971 3451
rect 91971 3417 91980 3451
rect 91928 3408 91980 3417
rect 89812 3340 89864 3392
rect 95056 3408 95108 3460
rect 98828 3680 98880 3732
rect 98920 3680 98972 3732
rect 98644 3612 98696 3664
rect 99104 3655 99156 3664
rect 99104 3621 99113 3655
rect 99113 3621 99147 3655
rect 99147 3621 99156 3655
rect 99104 3612 99156 3621
rect 99472 3612 99524 3664
rect 104164 3612 104216 3664
rect 104532 3680 104584 3732
rect 96620 3587 96672 3596
rect 96620 3553 96629 3587
rect 96629 3553 96663 3587
rect 96663 3553 96672 3587
rect 96620 3544 96672 3553
rect 97264 3587 97316 3596
rect 97264 3553 97273 3587
rect 97273 3553 97307 3587
rect 97307 3553 97316 3587
rect 97264 3544 97316 3553
rect 97540 3587 97592 3596
rect 97540 3553 97549 3587
rect 97549 3553 97583 3587
rect 97583 3553 97592 3587
rect 97540 3544 97592 3553
rect 100576 3544 100628 3596
rect 101312 3587 101364 3596
rect 101312 3553 101321 3587
rect 101321 3553 101355 3587
rect 101355 3553 101364 3587
rect 101312 3544 101364 3553
rect 101404 3544 101456 3596
rect 102876 3544 102928 3596
rect 103796 3587 103848 3596
rect 103796 3553 103805 3587
rect 103805 3553 103839 3587
rect 103839 3553 103848 3587
rect 103796 3544 103848 3553
rect 104532 3544 104584 3596
rect 105268 3544 105320 3596
rect 105452 3612 105504 3664
rect 112720 3612 112772 3664
rect 96712 3476 96764 3528
rect 97816 3519 97868 3528
rect 97816 3485 97825 3519
rect 97825 3485 97859 3519
rect 97859 3485 97868 3519
rect 97816 3476 97868 3485
rect 98736 3476 98788 3528
rect 101496 3476 101548 3528
rect 104164 3476 104216 3528
rect 97264 3340 97316 3392
rect 98460 3383 98512 3392
rect 98460 3349 98469 3383
rect 98469 3349 98503 3383
rect 98503 3349 98512 3383
rect 98460 3340 98512 3349
rect 98644 3340 98696 3392
rect 99104 3408 99156 3460
rect 99472 3340 99524 3392
rect 99748 3408 99800 3460
rect 101312 3340 101364 3392
rect 103152 3340 103204 3392
rect 104624 3340 104676 3392
rect 104900 3408 104952 3460
rect 106924 3340 106976 3392
rect 108856 3544 108908 3596
rect 110512 3587 110564 3596
rect 110512 3553 110521 3587
rect 110521 3553 110555 3587
rect 110555 3553 110564 3587
rect 110512 3544 110564 3553
rect 110972 3544 111024 3596
rect 113456 3680 113508 3732
rect 115848 3680 115900 3732
rect 115940 3680 115992 3732
rect 116768 3723 116820 3732
rect 116768 3689 116777 3723
rect 116777 3689 116811 3723
rect 116811 3689 116820 3723
rect 116768 3680 116820 3689
rect 152372 3680 152424 3732
rect 152832 3680 152884 3732
rect 155684 3680 155736 3732
rect 158260 3680 158312 3732
rect 158628 3680 158680 3732
rect 119804 3655 119856 3664
rect 119804 3621 119813 3655
rect 119813 3621 119847 3655
rect 119847 3621 119856 3655
rect 119804 3612 119856 3621
rect 121000 3655 121052 3664
rect 121000 3621 121009 3655
rect 121009 3621 121043 3655
rect 121043 3621 121052 3655
rect 121000 3612 121052 3621
rect 143448 3612 143500 3664
rect 144736 3612 144788 3664
rect 144828 3612 144880 3664
rect 112996 3544 113048 3596
rect 115296 3544 115348 3596
rect 115664 3544 115716 3596
rect 117228 3544 117280 3596
rect 118976 3544 119028 3596
rect 120080 3587 120132 3596
rect 120080 3553 120089 3587
rect 120089 3553 120123 3587
rect 120123 3553 120132 3587
rect 120080 3544 120132 3553
rect 120356 3587 120408 3596
rect 120356 3553 120365 3587
rect 120365 3553 120399 3587
rect 120399 3553 120408 3587
rect 120356 3544 120408 3553
rect 109316 3451 109368 3460
rect 109316 3417 109325 3451
rect 109325 3417 109359 3451
rect 109359 3417 109368 3451
rect 109316 3408 109368 3417
rect 113180 3340 113232 3392
rect 114928 3519 114980 3528
rect 114928 3485 114937 3519
rect 114937 3485 114971 3519
rect 114971 3485 114980 3519
rect 114928 3476 114980 3485
rect 115112 3519 115164 3528
rect 115112 3485 115121 3519
rect 115121 3485 115155 3519
rect 115155 3485 115164 3519
rect 115112 3476 115164 3485
rect 116124 3519 116176 3528
rect 116124 3485 116133 3519
rect 116133 3485 116167 3519
rect 116167 3485 116176 3519
rect 116124 3476 116176 3485
rect 119344 3519 119396 3528
rect 119344 3485 119353 3519
rect 119353 3485 119387 3519
rect 119387 3485 119396 3519
rect 119344 3476 119396 3485
rect 120172 3519 120224 3528
rect 120172 3485 120206 3519
rect 120206 3485 120224 3519
rect 120172 3476 120224 3485
rect 141424 3544 141476 3596
rect 142988 3544 143040 3596
rect 144000 3587 144052 3596
rect 144000 3553 144009 3587
rect 144009 3553 144043 3587
rect 144043 3553 144052 3587
rect 144000 3544 144052 3553
rect 144644 3544 144696 3596
rect 145380 3587 145432 3596
rect 145380 3553 145389 3587
rect 145389 3553 145423 3587
rect 145423 3553 145432 3587
rect 145380 3544 145432 3553
rect 122564 3519 122616 3528
rect 122564 3485 122573 3519
rect 122573 3485 122607 3519
rect 122607 3485 122616 3519
rect 122564 3476 122616 3485
rect 138940 3519 138992 3528
rect 138940 3485 138949 3519
rect 138949 3485 138983 3519
rect 138983 3485 138992 3519
rect 138940 3476 138992 3485
rect 143172 3476 143224 3528
rect 144276 3519 144328 3528
rect 144276 3485 144285 3519
rect 144285 3485 144319 3519
rect 144319 3485 144328 3519
rect 144276 3476 144328 3485
rect 139124 3451 139176 3460
rect 139124 3417 139133 3451
rect 139133 3417 139167 3451
rect 139167 3417 139176 3451
rect 139124 3408 139176 3417
rect 140688 3408 140740 3460
rect 144828 3408 144880 3460
rect 147956 3612 148008 3664
rect 148048 3612 148100 3664
rect 154488 3612 154540 3664
rect 156052 3612 156104 3664
rect 161020 3680 161072 3732
rect 161940 3680 161992 3732
rect 173164 3680 173216 3732
rect 207480 3680 207532 3732
rect 162676 3612 162728 3664
rect 210056 3655 210108 3664
rect 148968 3544 149020 3596
rect 154580 3544 154632 3596
rect 156328 3587 156380 3596
rect 156328 3553 156337 3587
rect 156337 3553 156371 3587
rect 156371 3553 156380 3587
rect 156328 3544 156380 3553
rect 156604 3587 156656 3596
rect 156604 3553 156613 3587
rect 156613 3553 156647 3587
rect 156647 3553 156656 3587
rect 156604 3544 156656 3553
rect 156696 3587 156748 3596
rect 156696 3553 156730 3587
rect 156730 3553 156748 3587
rect 156696 3544 156748 3553
rect 156880 3587 156932 3596
rect 156880 3553 156889 3587
rect 156889 3553 156923 3587
rect 156923 3553 156932 3587
rect 156880 3544 156932 3553
rect 158352 3587 158404 3596
rect 158352 3553 158361 3587
rect 158361 3553 158395 3587
rect 158395 3553 158404 3587
rect 158352 3544 158404 3553
rect 159272 3587 159324 3596
rect 159272 3553 159281 3587
rect 159281 3553 159315 3587
rect 159315 3553 159324 3587
rect 159272 3544 159324 3553
rect 159548 3587 159600 3596
rect 159548 3553 159557 3587
rect 159557 3553 159591 3587
rect 159591 3553 159600 3587
rect 159548 3544 159600 3553
rect 122840 3383 122892 3392
rect 122840 3349 122849 3383
rect 122849 3349 122883 3383
rect 122883 3349 122892 3383
rect 122840 3340 122892 3349
rect 138572 3340 138624 3392
rect 143816 3340 143868 3392
rect 146300 3519 146352 3528
rect 146300 3485 146309 3519
rect 146309 3485 146343 3519
rect 146343 3485 146352 3519
rect 146300 3476 146352 3485
rect 146484 3476 146536 3528
rect 147496 3476 147548 3528
rect 152372 3476 152424 3528
rect 154672 3476 154724 3528
rect 155224 3519 155276 3528
rect 155224 3485 155233 3519
rect 155233 3485 155267 3519
rect 155267 3485 155276 3519
rect 155224 3476 155276 3485
rect 155868 3519 155920 3528
rect 155868 3485 155877 3519
rect 155877 3485 155911 3519
rect 155911 3485 155920 3519
rect 155868 3476 155920 3485
rect 158536 3519 158588 3528
rect 158536 3485 158545 3519
rect 158545 3485 158579 3519
rect 158579 3485 158588 3519
rect 158536 3476 158588 3485
rect 159456 3476 159508 3528
rect 148416 3451 148468 3460
rect 148416 3417 148425 3451
rect 148425 3417 148459 3451
rect 148459 3417 148468 3451
rect 148416 3408 148468 3417
rect 148692 3408 148744 3460
rect 148876 3408 148928 3460
rect 150072 3451 150124 3460
rect 150072 3417 150081 3451
rect 150081 3417 150115 3451
rect 150115 3417 150124 3451
rect 150072 3408 150124 3417
rect 151176 3408 151228 3460
rect 154856 3408 154908 3460
rect 146852 3340 146904 3392
rect 149152 3340 149204 3392
rect 154396 3340 154448 3392
rect 156880 3340 156932 3392
rect 156972 3340 157024 3392
rect 176660 3544 176712 3596
rect 205088 3544 205140 3596
rect 160836 3519 160888 3528
rect 160836 3485 160845 3519
rect 160845 3485 160879 3519
rect 160879 3485 160888 3519
rect 160836 3476 160888 3485
rect 162492 3476 162544 3528
rect 204260 3476 204312 3528
rect 204904 3519 204956 3528
rect 204904 3485 204913 3519
rect 204913 3485 204947 3519
rect 204947 3485 204956 3519
rect 204904 3476 204956 3485
rect 207204 3587 207256 3596
rect 207204 3553 207213 3587
rect 207213 3553 207247 3587
rect 207247 3553 207256 3587
rect 207204 3544 207256 3553
rect 207664 3587 207716 3596
rect 207664 3553 207673 3587
rect 207673 3553 207707 3587
rect 207707 3553 207716 3587
rect 210056 3621 210065 3655
rect 210065 3621 210099 3655
rect 210099 3621 210108 3655
rect 210056 3612 210108 3621
rect 207664 3544 207716 3553
rect 161296 3408 161348 3460
rect 162676 3451 162728 3460
rect 162676 3417 162685 3451
rect 162685 3417 162719 3451
rect 162719 3417 162728 3451
rect 162676 3408 162728 3417
rect 163412 3408 163464 3460
rect 180892 3408 180944 3460
rect 205088 3451 205140 3460
rect 205088 3417 205097 3451
rect 205097 3417 205131 3451
rect 205131 3417 205140 3451
rect 205088 3408 205140 3417
rect 160560 3383 160612 3392
rect 160560 3349 160569 3383
rect 160569 3349 160603 3383
rect 160603 3349 160612 3383
rect 160560 3340 160612 3349
rect 160652 3340 160704 3392
rect 207112 3408 207164 3460
rect 207756 3408 207808 3460
rect 208400 3340 208452 3392
rect 209688 3408 209740 3460
rect 210332 3408 210384 3460
rect 210148 3340 210200 3392
rect 224500 3680 224552 3732
rect 225236 3680 225288 3732
rect 210608 3612 210660 3664
rect 210700 3587 210752 3596
rect 210700 3553 210709 3587
rect 210709 3553 210743 3587
rect 210743 3553 210752 3587
rect 210700 3544 210752 3553
rect 211252 3544 211304 3596
rect 213092 3587 213144 3596
rect 213092 3553 213101 3587
rect 213101 3553 213135 3587
rect 213135 3553 213144 3587
rect 213092 3544 213144 3553
rect 214656 3612 214708 3664
rect 215760 3612 215812 3664
rect 214380 3544 214432 3596
rect 216128 3587 216180 3596
rect 216128 3553 216137 3587
rect 216137 3553 216171 3587
rect 216171 3553 216180 3587
rect 216128 3544 216180 3553
rect 217416 3612 217468 3664
rect 217508 3612 217560 3664
rect 226248 3612 226300 3664
rect 227352 3723 227404 3732
rect 227352 3689 227361 3723
rect 227361 3689 227395 3723
rect 227395 3689 227404 3723
rect 227352 3680 227404 3689
rect 251456 3680 251508 3732
rect 256516 3680 256568 3732
rect 258540 3680 258592 3732
rect 265348 3723 265400 3732
rect 265348 3689 265357 3723
rect 265357 3689 265391 3723
rect 265391 3689 265400 3723
rect 265348 3680 265400 3689
rect 265992 3723 266044 3732
rect 265992 3689 266001 3723
rect 266001 3689 266035 3723
rect 266035 3689 266044 3723
rect 265992 3680 266044 3689
rect 238576 3612 238628 3664
rect 259920 3612 259972 3664
rect 268016 3612 268068 3664
rect 269488 3680 269540 3732
rect 270592 3680 270644 3732
rect 270776 3680 270828 3732
rect 269212 3612 269264 3664
rect 269580 3612 269632 3664
rect 269856 3612 269908 3664
rect 218888 3587 218940 3596
rect 218888 3553 218897 3587
rect 218897 3553 218931 3587
rect 218931 3553 218940 3587
rect 218888 3544 218940 3553
rect 224960 3544 225012 3596
rect 212540 3476 212592 3528
rect 213368 3519 213420 3528
rect 213368 3485 213377 3519
rect 213377 3485 213411 3519
rect 213411 3485 213420 3519
rect 213368 3476 213420 3485
rect 213460 3519 213512 3528
rect 213460 3485 213494 3519
rect 213494 3485 213512 3519
rect 213460 3476 213512 3485
rect 213644 3519 213696 3528
rect 213644 3485 213653 3519
rect 213653 3485 213687 3519
rect 213687 3485 213696 3519
rect 213644 3476 213696 3485
rect 215392 3519 215444 3528
rect 215392 3485 215401 3519
rect 215401 3485 215435 3519
rect 215435 3485 215444 3519
rect 215392 3476 215444 3485
rect 216404 3519 216456 3528
rect 216404 3485 216413 3519
rect 216413 3485 216447 3519
rect 216447 3485 216456 3519
rect 216404 3476 216456 3485
rect 217232 3476 217284 3528
rect 219164 3476 219216 3528
rect 212356 3451 212408 3460
rect 212356 3417 212365 3451
rect 212365 3417 212399 3451
rect 212399 3417 212408 3451
rect 212356 3408 212408 3417
rect 215852 3340 215904 3392
rect 216496 3340 216548 3392
rect 217416 3383 217468 3392
rect 217416 3349 217425 3383
rect 217425 3349 217459 3383
rect 217459 3349 217468 3383
rect 217416 3340 217468 3349
rect 220176 3408 220228 3460
rect 222752 3519 222804 3528
rect 222752 3485 222761 3519
rect 222761 3485 222795 3519
rect 222795 3485 222804 3519
rect 222752 3476 222804 3485
rect 225144 3544 225196 3596
rect 226156 3587 226208 3596
rect 226156 3553 226165 3587
rect 226165 3553 226199 3587
rect 226199 3553 226208 3587
rect 226156 3544 226208 3553
rect 227720 3544 227772 3596
rect 225696 3519 225748 3528
rect 225696 3485 225705 3519
rect 225705 3485 225739 3519
rect 225739 3485 225748 3519
rect 225696 3476 225748 3485
rect 226432 3519 226484 3528
rect 226432 3485 226441 3519
rect 226441 3485 226475 3519
rect 226475 3485 226484 3519
rect 226432 3476 226484 3485
rect 226708 3519 226760 3528
rect 226708 3485 226717 3519
rect 226717 3485 226751 3519
rect 226751 3485 226760 3519
rect 226708 3476 226760 3485
rect 225604 3408 225656 3460
rect 231492 3476 231544 3528
rect 242900 3544 242952 3596
rect 253940 3544 253992 3596
rect 268108 3544 268160 3596
rect 248972 3476 249024 3528
rect 251916 3476 251968 3528
rect 258080 3519 258132 3528
rect 258080 3485 258089 3519
rect 258089 3485 258123 3519
rect 258123 3485 258132 3519
rect 258080 3476 258132 3485
rect 258264 3476 258316 3528
rect 229192 3408 229244 3460
rect 251456 3408 251508 3460
rect 227720 3383 227772 3392
rect 227720 3349 227729 3383
rect 227729 3349 227763 3383
rect 227763 3349 227772 3383
rect 227720 3340 227772 3349
rect 229836 3340 229888 3392
rect 230756 3340 230808 3392
rect 242992 3340 243044 3392
rect 257620 3408 257672 3460
rect 260840 3476 260892 3528
rect 266084 3476 266136 3528
rect 266176 3519 266228 3528
rect 266176 3485 266185 3519
rect 266185 3485 266219 3519
rect 266219 3485 266228 3519
rect 266176 3476 266228 3485
rect 267372 3519 267424 3528
rect 267372 3485 267381 3519
rect 267381 3485 267415 3519
rect 267415 3485 267424 3519
rect 267372 3476 267424 3485
rect 267740 3476 267792 3528
rect 260012 3408 260064 3460
rect 267648 3408 267700 3460
rect 268200 3476 268252 3528
rect 268752 3476 268804 3528
rect 269948 3476 270000 3528
rect 269028 3408 269080 3460
rect 271972 3408 272024 3460
rect 252376 3383 252428 3392
rect 252376 3349 252385 3383
rect 252385 3349 252419 3383
rect 252419 3349 252428 3383
rect 252376 3340 252428 3349
rect 265624 3340 265676 3392
rect 267740 3340 267792 3392
rect 270040 3340 270092 3392
rect 68546 3238 68598 3290
rect 68610 3238 68662 3290
rect 68674 3238 68726 3290
rect 68738 3238 68790 3290
rect 68802 3238 68854 3290
rect 136143 3238 136195 3290
rect 136207 3238 136259 3290
rect 136271 3238 136323 3290
rect 136335 3238 136387 3290
rect 136399 3238 136451 3290
rect 203740 3238 203792 3290
rect 203804 3238 203856 3290
rect 203868 3238 203920 3290
rect 203932 3238 203984 3290
rect 203996 3238 204048 3290
rect 271337 3238 271389 3290
rect 271401 3238 271453 3290
rect 271465 3238 271517 3290
rect 271529 3238 271581 3290
rect 271593 3238 271645 3290
rect 27252 3136 27304 3188
rect 37556 3136 37608 3188
rect 23848 3000 23900 3052
rect 19248 2932 19300 2984
rect 24860 2932 24912 2984
rect 25228 2975 25280 2984
rect 25228 2941 25237 2975
rect 25237 2941 25271 2975
rect 25271 2941 25280 2975
rect 25228 2932 25280 2941
rect 22928 2864 22980 2916
rect 19984 2796 20036 2848
rect 26332 3068 26384 3120
rect 27068 3068 27120 3120
rect 25412 3043 25464 3052
rect 25412 3009 25421 3043
rect 25421 3009 25455 3043
rect 25455 3009 25464 3043
rect 25412 3000 25464 3009
rect 26148 3000 26200 3052
rect 26056 2975 26108 2984
rect 26056 2941 26065 2975
rect 26065 2941 26099 2975
rect 26099 2941 26108 2975
rect 27620 3068 27672 3120
rect 35900 3068 35952 3120
rect 27896 3000 27948 3052
rect 27988 3043 28040 3052
rect 27988 3009 27997 3043
rect 27997 3009 28031 3043
rect 28031 3009 28040 3043
rect 27988 3000 28040 3009
rect 26056 2932 26108 2941
rect 25596 2839 25648 2848
rect 25596 2805 25605 2839
rect 25605 2805 25639 2839
rect 25639 2805 25648 2839
rect 25596 2796 25648 2805
rect 26424 2839 26476 2848
rect 26424 2805 26433 2839
rect 26433 2805 26467 2839
rect 26467 2805 26476 2839
rect 26424 2796 26476 2805
rect 38016 3068 38068 3120
rect 38108 3111 38160 3120
rect 38108 3077 38117 3111
rect 38117 3077 38151 3111
rect 38151 3077 38160 3111
rect 38108 3068 38160 3077
rect 38200 3111 38252 3120
rect 38200 3077 38209 3111
rect 38209 3077 38243 3111
rect 38243 3077 38252 3111
rect 38200 3068 38252 3077
rect 38568 3111 38620 3120
rect 38568 3077 38577 3111
rect 38577 3077 38611 3111
rect 38611 3077 38620 3111
rect 38568 3068 38620 3077
rect 38936 3111 38988 3120
rect 38936 3077 38945 3111
rect 38945 3077 38979 3111
rect 38979 3077 38988 3111
rect 38936 3068 38988 3077
rect 39856 3111 39908 3120
rect 39856 3077 39865 3111
rect 39865 3077 39899 3111
rect 39899 3077 39908 3111
rect 39856 3068 39908 3077
rect 40132 3111 40184 3120
rect 40132 3077 40141 3111
rect 40141 3077 40175 3111
rect 40175 3077 40184 3111
rect 40132 3068 40184 3077
rect 40500 3068 40552 3120
rect 41052 3068 41104 3120
rect 37188 3000 37240 3052
rect 38476 3000 38528 3052
rect 39948 3000 40000 3052
rect 40224 3043 40276 3052
rect 40224 3009 40233 3043
rect 40233 3009 40267 3043
rect 40267 3009 40276 3043
rect 40224 3000 40276 3009
rect 40776 3000 40828 3052
rect 52276 3136 52328 3188
rect 81440 3136 81492 3188
rect 41880 3068 41932 3120
rect 86040 3068 86092 3120
rect 98644 3136 98696 3188
rect 98736 3179 98788 3188
rect 98736 3145 98745 3179
rect 98745 3145 98779 3179
rect 98779 3145 98788 3179
rect 98736 3136 98788 3145
rect 101496 3179 101548 3188
rect 101496 3145 101505 3179
rect 101505 3145 101539 3179
rect 101539 3145 101548 3179
rect 101496 3136 101548 3145
rect 102048 3136 102100 3188
rect 54116 3000 54168 3052
rect 82360 3043 82412 3052
rect 82360 3009 82369 3043
rect 82369 3009 82403 3043
rect 82403 3009 82412 3043
rect 82360 3000 82412 3009
rect 86592 3043 86644 3052
rect 86592 3009 86601 3043
rect 86601 3009 86635 3043
rect 86635 3009 86644 3043
rect 86592 3000 86644 3009
rect 40960 2932 41012 2984
rect 67548 2932 67600 2984
rect 82084 2975 82136 2984
rect 82084 2941 82093 2975
rect 82093 2941 82127 2975
rect 82127 2941 82136 2975
rect 82084 2932 82136 2941
rect 84292 2975 84344 2984
rect 84292 2941 84301 2975
rect 84301 2941 84335 2975
rect 84335 2941 84344 2975
rect 84292 2932 84344 2941
rect 84476 2975 84528 2984
rect 84476 2941 84485 2975
rect 84485 2941 84519 2975
rect 84519 2941 84528 2975
rect 84476 2932 84528 2941
rect 86776 2975 86828 2984
rect 86776 2941 86785 2975
rect 86785 2941 86819 2975
rect 86819 2941 86828 2975
rect 86776 2932 86828 2941
rect 28080 2864 28132 2916
rect 39120 2907 39172 2916
rect 39120 2873 39129 2907
rect 39129 2873 39163 2907
rect 39163 2873 39172 2907
rect 39120 2864 39172 2873
rect 41144 2907 41196 2916
rect 41144 2873 41153 2907
rect 41153 2873 41187 2907
rect 41187 2873 41196 2907
rect 41144 2864 41196 2873
rect 73160 2864 73212 2916
rect 27712 2839 27764 2848
rect 27712 2805 27721 2839
rect 27721 2805 27755 2839
rect 27755 2805 27764 2839
rect 27712 2796 27764 2805
rect 30932 2796 30984 2848
rect 37464 2796 37516 2848
rect 106280 3136 106332 3188
rect 89168 3043 89220 3052
rect 89168 3009 89177 3043
rect 89177 3009 89211 3043
rect 89211 3009 89220 3043
rect 89168 3000 89220 3009
rect 92296 3043 92348 3052
rect 92296 3009 92305 3043
rect 92305 3009 92339 3043
rect 92339 3009 92348 3043
rect 92296 3000 92348 3009
rect 94228 3043 94280 3052
rect 94228 3009 94237 3043
rect 94237 3009 94271 3043
rect 94271 3009 94280 3043
rect 94228 3000 94280 3009
rect 96068 3043 96120 3052
rect 96068 3009 96077 3043
rect 96077 3009 96111 3043
rect 96111 3009 96120 3043
rect 96068 3000 96120 3009
rect 96896 3043 96948 3052
rect 96896 3009 96905 3043
rect 96905 3009 96939 3043
rect 96939 3009 96948 3043
rect 96896 3000 96948 3009
rect 109500 3068 109552 3120
rect 98092 3043 98144 3052
rect 98092 3009 98101 3043
rect 98101 3009 98135 3043
rect 98135 3009 98144 3043
rect 98092 3000 98144 3009
rect 99656 3043 99708 3052
rect 99656 3009 99665 3043
rect 99665 3009 99699 3043
rect 99699 3009 99708 3043
rect 99656 3000 99708 3009
rect 101680 3043 101732 3052
rect 101680 3009 101689 3043
rect 101689 3009 101723 3043
rect 101723 3009 101732 3043
rect 101680 3000 101732 3009
rect 90088 2975 90140 2984
rect 90088 2941 90097 2975
rect 90097 2941 90131 2975
rect 90131 2941 90140 2975
rect 90088 2932 90140 2941
rect 90272 2975 90324 2984
rect 90272 2941 90281 2975
rect 90281 2941 90315 2975
rect 90315 2941 90324 2975
rect 90272 2932 90324 2941
rect 91652 2932 91704 2984
rect 89812 2864 89864 2916
rect 93768 2932 93820 2984
rect 97172 2932 97224 2984
rect 99472 2932 99524 2984
rect 99840 2975 99892 2984
rect 99840 2941 99849 2975
rect 99849 2941 99883 2975
rect 99883 2941 99892 2975
rect 99840 2932 99892 2941
rect 100392 2932 100444 2984
rect 100668 2975 100720 2984
rect 100668 2941 100702 2975
rect 100702 2941 100720 2975
rect 100668 2932 100720 2941
rect 101404 2932 101456 2984
rect 101864 2975 101916 2984
rect 101864 2941 101873 2975
rect 101873 2941 101907 2975
rect 101907 2941 101916 2975
rect 101864 2932 101916 2941
rect 102232 2932 102284 2984
rect 102600 3009 102627 3018
rect 102627 3009 102652 3018
rect 102600 2966 102652 3009
rect 102876 3043 102928 3052
rect 102876 3009 102885 3043
rect 102885 3009 102919 3043
rect 102919 3009 102928 3043
rect 102876 3000 102928 3009
rect 92296 2864 92348 2916
rect 89352 2839 89404 2848
rect 89352 2805 89361 2839
rect 89361 2805 89395 2839
rect 89395 2805 89404 2839
rect 89352 2796 89404 2805
rect 96804 2796 96856 2848
rect 96988 2796 97040 2848
rect 97356 2796 97408 2848
rect 99932 2864 99984 2916
rect 104624 2975 104676 2984
rect 104624 2941 104633 2975
rect 104633 2941 104667 2975
rect 104667 2941 104676 2975
rect 104624 2932 104676 2941
rect 107108 3043 107160 3052
rect 107108 3009 107117 3043
rect 107117 3009 107151 3043
rect 107151 3009 107160 3043
rect 107108 3000 107160 3009
rect 109316 3000 109368 3052
rect 112720 3068 112772 3120
rect 116676 3068 116728 3120
rect 117688 3068 117740 3120
rect 110236 3043 110288 3052
rect 110236 3009 110245 3043
rect 110245 3009 110279 3043
rect 110279 3009 110288 3043
rect 110236 3000 110288 3009
rect 107292 2975 107344 2984
rect 106188 2864 106240 2916
rect 103336 2796 103388 2848
rect 107292 2941 107301 2975
rect 107301 2941 107335 2975
rect 107335 2941 107344 2975
rect 107292 2932 107344 2941
rect 107660 2975 107712 2984
rect 107660 2941 107669 2975
rect 107669 2941 107703 2975
rect 107703 2941 107712 2975
rect 107660 2932 107712 2941
rect 109684 2932 109736 2984
rect 115940 3000 115992 3052
rect 116124 3000 116176 3052
rect 116492 3043 116544 3052
rect 116492 3009 116501 3043
rect 116501 3009 116535 3043
rect 116535 3009 116544 3043
rect 116492 3000 116544 3009
rect 113548 2932 113600 2984
rect 116308 2932 116360 2984
rect 114652 2864 114704 2916
rect 115756 2907 115808 2916
rect 115756 2873 115765 2907
rect 115765 2873 115799 2907
rect 115799 2873 115808 2907
rect 115756 2864 115808 2873
rect 116952 2975 117004 2984
rect 116952 2941 116961 2975
rect 116961 2941 116995 2975
rect 116995 2941 117004 2975
rect 116952 2932 117004 2941
rect 120632 3111 120684 3120
rect 120632 3077 120641 3111
rect 120641 3077 120675 3111
rect 120675 3077 120684 3111
rect 120632 3068 120684 3077
rect 123576 3068 123628 3120
rect 120264 3000 120316 3052
rect 121920 2932 121972 2984
rect 116952 2796 117004 2848
rect 124312 2796 124364 2848
rect 138940 3136 138992 3188
rect 141792 3136 141844 3188
rect 144828 3136 144880 3188
rect 137744 3043 137796 3052
rect 137744 3009 137753 3043
rect 137753 3009 137787 3043
rect 137787 3009 137796 3043
rect 137744 3000 137796 3009
rect 138664 3043 138716 3052
rect 138664 3009 138673 3043
rect 138673 3009 138707 3043
rect 138707 3009 138716 3043
rect 138664 3000 138716 3009
rect 137928 2975 137980 2984
rect 137928 2941 137937 2975
rect 137937 2941 137971 2975
rect 137971 2941 137980 2975
rect 137928 2932 137980 2941
rect 138756 2975 138808 2984
rect 138756 2941 138790 2975
rect 138790 2941 138808 2975
rect 138756 2932 138808 2941
rect 138940 2975 138992 2984
rect 138940 2941 138949 2975
rect 138949 2941 138983 2975
rect 138983 2941 138992 2975
rect 138940 2932 138992 2941
rect 139124 2932 139176 2984
rect 142160 3068 142212 3120
rect 147496 3179 147548 3188
rect 147496 3145 147505 3179
rect 147505 3145 147539 3179
rect 147539 3145 147548 3179
rect 147496 3136 147548 3145
rect 148140 3136 148192 3188
rect 148048 3068 148100 3120
rect 141884 3000 141936 3052
rect 143724 3043 143776 3052
rect 143724 3009 143733 3043
rect 143733 3009 143767 3043
rect 143767 3009 143776 3043
rect 143724 3000 143776 3009
rect 138388 2907 138440 2916
rect 138388 2873 138397 2907
rect 138397 2873 138431 2907
rect 138431 2873 138440 2907
rect 138388 2864 138440 2873
rect 140780 2864 140832 2916
rect 142712 2932 142764 2984
rect 143448 2975 143500 2984
rect 143448 2941 143457 2975
rect 143457 2941 143491 2975
rect 143491 2941 143500 2975
rect 143448 2932 143500 2941
rect 143908 2932 143960 2984
rect 144000 2975 144052 2984
rect 144000 2941 144009 2975
rect 144009 2941 144043 2975
rect 144043 2941 144052 2975
rect 144000 2932 144052 2941
rect 144368 2932 144420 2984
rect 146576 3043 146628 3052
rect 146576 3009 146585 3043
rect 146585 3009 146619 3043
rect 146619 3009 146628 3043
rect 146576 3000 146628 3009
rect 146852 3043 146904 3052
rect 146852 3009 146861 3043
rect 146861 3009 146895 3043
rect 146895 3009 146904 3043
rect 146852 3000 146904 3009
rect 147772 3000 147824 3052
rect 148876 3043 148928 3052
rect 148876 3009 148885 3043
rect 148885 3009 148919 3043
rect 148919 3009 148928 3043
rect 148876 3000 148928 3009
rect 149152 3043 149204 3052
rect 149152 3009 149161 3043
rect 149161 3009 149195 3043
rect 149195 3009 149204 3043
rect 149152 3000 149204 3009
rect 145564 2932 145616 2984
rect 146760 2932 146812 2984
rect 148140 2975 148192 2984
rect 148140 2941 148149 2975
rect 148149 2941 148183 2975
rect 148183 2941 148192 2975
rect 148140 2932 148192 2941
rect 142712 2796 142764 2848
rect 144828 2796 144880 2848
rect 148692 2932 148744 2984
rect 148968 2975 149020 2984
rect 148968 2941 149002 2975
rect 149002 2941 149020 2975
rect 148968 2932 149020 2941
rect 150992 3136 151044 3188
rect 152924 3068 152976 3120
rect 155960 3043 156012 3052
rect 155960 3009 155969 3043
rect 155969 3009 156003 3043
rect 156003 3009 156012 3043
rect 155960 3000 156012 3009
rect 156144 3068 156196 3120
rect 157892 3068 157944 3120
rect 160836 3068 160888 3120
rect 149244 2796 149296 2848
rect 156144 2975 156196 2984
rect 156144 2941 156153 2975
rect 156153 2941 156187 2975
rect 156187 2941 156196 2975
rect 156144 2932 156196 2941
rect 156880 3043 156932 3052
rect 156880 3009 156889 3043
rect 156889 3009 156923 3043
rect 156923 3009 156932 3043
rect 156880 3000 156932 3009
rect 156972 3043 157024 3052
rect 156972 3009 157006 3043
rect 157006 3009 157024 3043
rect 156972 3000 157024 3009
rect 157984 2932 158036 2984
rect 158812 3043 158864 3052
rect 158812 3009 158821 3043
rect 158821 3009 158855 3043
rect 158855 3009 158864 3043
rect 158812 3000 158864 3009
rect 158904 3043 158956 3052
rect 158904 3009 158938 3043
rect 158938 3009 158956 3043
rect 158904 3000 158956 3009
rect 160192 3043 160244 3052
rect 160192 3009 160201 3043
rect 160201 3009 160235 3043
rect 160235 3009 160244 3043
rect 160560 3043 160612 3052
rect 160192 3000 160244 3009
rect 160560 3009 160569 3043
rect 160569 3009 160603 3043
rect 160603 3009 160612 3043
rect 162676 3068 162728 3120
rect 175924 3068 175976 3120
rect 204904 3136 204956 3188
rect 213368 3136 213420 3188
rect 213920 3136 213972 3188
rect 214472 3179 214524 3188
rect 214472 3145 214481 3179
rect 214481 3145 214515 3179
rect 214515 3145 214524 3179
rect 214472 3136 214524 3145
rect 216036 3136 216088 3188
rect 217232 3179 217284 3188
rect 217232 3145 217241 3179
rect 217241 3145 217275 3179
rect 217275 3145 217284 3179
rect 217232 3136 217284 3145
rect 218704 3179 218756 3188
rect 218704 3145 218713 3179
rect 218713 3145 218747 3179
rect 218747 3145 218756 3179
rect 218704 3136 218756 3145
rect 207940 3068 207992 3120
rect 218060 3068 218112 3120
rect 218888 3068 218940 3120
rect 225696 3136 225748 3188
rect 226248 3136 226300 3188
rect 246212 3136 246264 3188
rect 252376 3136 252428 3188
rect 262220 3136 262272 3188
rect 264060 3136 264112 3188
rect 268476 3136 268528 3188
rect 269304 3136 269356 3188
rect 160560 3000 160612 3009
rect 162032 3000 162084 3052
rect 162952 3043 163004 3052
rect 162952 3009 162961 3043
rect 162961 3009 162995 3043
rect 162995 3009 163004 3043
rect 162952 3000 163004 3009
rect 156604 2907 156656 2916
rect 156604 2873 156613 2907
rect 156613 2873 156647 2907
rect 156647 2873 156656 2907
rect 156604 2864 156656 2873
rect 161296 2932 161348 2984
rect 167736 2975 167788 2984
rect 167736 2941 167745 2975
rect 167745 2941 167779 2975
rect 167779 2941 167788 2975
rect 167736 2932 167788 2941
rect 202328 2975 202380 2984
rect 202328 2941 202337 2975
rect 202337 2941 202371 2975
rect 202371 2941 202380 2975
rect 202328 2932 202380 2941
rect 153108 2796 153160 2848
rect 156052 2796 156104 2848
rect 158628 2864 158680 2916
rect 159548 2864 159600 2916
rect 203800 2907 203852 2916
rect 203800 2873 203809 2907
rect 203809 2873 203843 2907
rect 203843 2873 203852 2907
rect 203800 2864 203852 2873
rect 158352 2796 158404 2848
rect 160652 2796 160704 2848
rect 163136 2839 163188 2848
rect 163136 2805 163145 2839
rect 163145 2805 163179 2839
rect 163179 2805 163188 2839
rect 163136 2796 163188 2805
rect 205088 2932 205140 2984
rect 204444 2864 204496 2916
rect 207204 3000 207256 3052
rect 207388 3000 207440 3052
rect 208676 3043 208728 3052
rect 208676 3009 208685 3043
rect 208685 3009 208719 3043
rect 208719 3009 208728 3043
rect 208676 3000 208728 3009
rect 210976 3043 211028 3052
rect 210976 3009 210985 3043
rect 210985 3009 211019 3043
rect 211019 3009 211028 3043
rect 210976 3000 211028 3009
rect 211068 3043 211120 3052
rect 211068 3009 211102 3043
rect 211102 3009 211120 3043
rect 211068 3000 211120 3009
rect 212172 3000 212224 3052
rect 213552 3043 213604 3052
rect 213552 3009 213561 3043
rect 213561 3009 213595 3043
rect 213595 3009 213604 3043
rect 213552 3000 213604 3009
rect 213736 3000 213788 3052
rect 206376 2932 206428 2984
rect 208400 2975 208452 2984
rect 208400 2941 208409 2975
rect 208409 2941 208443 2975
rect 208443 2941 208452 2975
rect 208400 2932 208452 2941
rect 208860 2932 208912 2984
rect 209596 2932 209648 2984
rect 210240 2975 210292 2984
rect 210240 2941 210249 2975
rect 210249 2941 210283 2975
rect 210283 2941 210292 2975
rect 210240 2932 210292 2941
rect 211252 2975 211304 2984
rect 211252 2941 211261 2975
rect 211261 2941 211295 2975
rect 211295 2941 211304 2975
rect 211252 2932 211304 2941
rect 211436 2932 211488 2984
rect 212816 2975 212868 2984
rect 212816 2941 212825 2975
rect 212825 2941 212859 2975
rect 212859 2941 212868 2975
rect 212816 2932 212868 2941
rect 214380 2932 214432 2984
rect 216312 3043 216364 3052
rect 216312 3009 216321 3043
rect 216321 3009 216355 3043
rect 216355 3009 216364 3043
rect 216312 3000 216364 3009
rect 216588 3043 216640 3052
rect 216588 3009 216597 3043
rect 216597 3009 216631 3043
rect 216631 3009 216640 3043
rect 216588 3000 216640 3009
rect 226064 3111 226116 3120
rect 226064 3077 226073 3111
rect 226073 3077 226107 3111
rect 226107 3077 226116 3111
rect 226064 3068 226116 3077
rect 226800 3068 226852 3120
rect 226984 3068 227036 3120
rect 230388 3068 230440 3120
rect 259736 3068 259788 3120
rect 259920 3068 259972 3120
rect 269948 3136 270000 3188
rect 271144 3136 271196 3188
rect 271972 3136 272024 3188
rect 223212 3043 223264 3052
rect 223212 3009 223221 3043
rect 223221 3009 223255 3043
rect 223255 3009 223264 3043
rect 223212 3000 223264 3009
rect 223304 3000 223356 3052
rect 226892 3000 226944 3052
rect 228088 3043 228140 3052
rect 228088 3009 228097 3043
rect 228097 3009 228131 3043
rect 228131 3009 228140 3043
rect 228088 3000 228140 3009
rect 215668 2932 215720 2984
rect 215760 2932 215812 2984
rect 216496 2932 216548 2984
rect 216772 2932 216824 2984
rect 218152 2932 218204 2984
rect 219072 2975 219124 2984
rect 219072 2941 219081 2975
rect 219081 2941 219115 2975
rect 219115 2941 219124 2975
rect 219072 2932 219124 2941
rect 221004 2932 221056 2984
rect 223580 2932 223632 2984
rect 226064 2932 226116 2984
rect 227628 2932 227680 2984
rect 242532 3000 242584 3052
rect 257988 3000 258040 3052
rect 259000 3043 259052 3052
rect 259000 3009 259009 3043
rect 259009 3009 259043 3043
rect 259043 3009 259052 3043
rect 259000 3000 259052 3009
rect 266268 3000 266320 3052
rect 266820 3043 266872 3052
rect 266820 3009 266829 3043
rect 266829 3009 266863 3043
rect 266863 3009 266872 3043
rect 266820 3000 266872 3009
rect 267464 3043 267516 3052
rect 267464 3009 267473 3043
rect 267473 3009 267507 3043
rect 267507 3009 267516 3043
rect 267464 3000 267516 3009
rect 268660 3000 268712 3052
rect 272064 3068 272116 3120
rect 269856 3043 269908 3052
rect 269856 3009 269865 3043
rect 269865 3009 269899 3043
rect 269899 3009 269908 3043
rect 269856 3000 269908 3009
rect 271880 3000 271932 3052
rect 210792 2796 210844 2848
rect 215760 2796 215812 2848
rect 217416 2864 217468 2916
rect 235816 2975 235868 2984
rect 235816 2941 235825 2975
rect 235825 2941 235859 2975
rect 235859 2941 235868 2975
rect 235816 2932 235868 2941
rect 236092 2932 236144 2984
rect 255320 2932 255372 2984
rect 262404 2932 262456 2984
rect 229836 2864 229888 2916
rect 246488 2864 246540 2916
rect 267188 2864 267240 2916
rect 268292 2932 268344 2984
rect 269120 2864 269172 2916
rect 216588 2796 216640 2848
rect 217784 2796 217836 2848
rect 219440 2839 219492 2848
rect 219440 2805 219449 2839
rect 219449 2805 219483 2839
rect 219483 2805 219492 2839
rect 219440 2796 219492 2805
rect 223488 2796 223540 2848
rect 226524 2796 226576 2848
rect 227260 2839 227312 2848
rect 227260 2805 227269 2839
rect 227269 2805 227303 2839
rect 227303 2805 227312 2839
rect 227260 2796 227312 2805
rect 228272 2839 228324 2848
rect 228272 2805 228281 2839
rect 228281 2805 228315 2839
rect 228315 2805 228324 2839
rect 228272 2796 228324 2805
rect 231676 2796 231728 2848
rect 238668 2796 238720 2848
rect 258080 2796 258132 2848
rect 259184 2839 259236 2848
rect 259184 2805 259193 2839
rect 259193 2805 259227 2839
rect 259227 2805 259236 2839
rect 259184 2796 259236 2805
rect 265532 2839 265584 2848
rect 265532 2805 265541 2839
rect 265541 2805 265575 2839
rect 265575 2805 265584 2839
rect 265532 2796 265584 2805
rect 266636 2839 266688 2848
rect 266636 2805 266645 2839
rect 266645 2805 266679 2839
rect 266679 2805 266688 2839
rect 266636 2796 266688 2805
rect 266820 2796 266872 2848
rect 268476 2796 268528 2848
rect 270500 2796 270552 2848
rect 34748 2694 34800 2746
rect 34812 2694 34864 2746
rect 34876 2694 34928 2746
rect 34940 2694 34992 2746
rect 35004 2694 35056 2746
rect 102345 2694 102397 2746
rect 102409 2694 102461 2746
rect 102473 2694 102525 2746
rect 102537 2694 102589 2746
rect 102601 2694 102653 2746
rect 169942 2694 169994 2746
rect 170006 2694 170058 2746
rect 170070 2694 170122 2746
rect 170134 2694 170186 2746
rect 170198 2694 170250 2746
rect 237539 2694 237591 2746
rect 237603 2694 237655 2746
rect 237667 2694 237719 2746
rect 237731 2694 237783 2746
rect 237795 2694 237847 2746
rect 23480 2592 23532 2644
rect 25780 2592 25832 2644
rect 26240 2635 26292 2644
rect 26240 2601 26249 2635
rect 26249 2601 26283 2635
rect 26283 2601 26292 2635
rect 26240 2592 26292 2601
rect 26516 2592 26568 2644
rect 27988 2592 28040 2644
rect 58900 2592 58952 2644
rect 60740 2592 60792 2644
rect 85396 2592 85448 2644
rect 4804 2524 4856 2576
rect 23572 2524 23624 2576
rect 25136 2524 25188 2576
rect 33140 2524 33192 2576
rect 70860 2524 70912 2576
rect 36636 2456 36688 2508
rect 37188 2456 37240 2508
rect 53748 2499 53800 2508
rect 53748 2465 53757 2499
rect 53757 2465 53791 2499
rect 53791 2465 53800 2499
rect 53748 2456 53800 2465
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 23756 2431 23808 2440
rect 23756 2397 23765 2431
rect 23765 2397 23799 2431
rect 23799 2397 23808 2431
rect 23756 2388 23808 2397
rect 24952 2431 25004 2440
rect 24952 2397 24961 2431
rect 24961 2397 24995 2431
rect 24995 2397 25004 2431
rect 24952 2388 25004 2397
rect 25044 2431 25096 2440
rect 25044 2397 25053 2431
rect 25053 2397 25087 2431
rect 25087 2397 25096 2431
rect 25044 2388 25096 2397
rect 25504 2388 25556 2440
rect 25688 2388 25740 2440
rect 2596 2320 2648 2372
rect 26148 2388 26200 2440
rect 26792 2431 26844 2440
rect 26792 2397 26801 2431
rect 26801 2397 26835 2431
rect 26835 2397 26844 2431
rect 26792 2388 26844 2397
rect 27344 2388 27396 2440
rect 27896 2431 27948 2440
rect 27896 2397 27905 2431
rect 27905 2397 27939 2431
rect 27939 2397 27948 2431
rect 27896 2388 27948 2397
rect 28540 2431 28592 2440
rect 28540 2397 28549 2431
rect 28549 2397 28583 2431
rect 28583 2397 28592 2431
rect 28540 2388 28592 2397
rect 31944 2388 31996 2440
rect 32496 2388 32548 2440
rect 38660 2388 38712 2440
rect 53472 2388 53524 2440
rect 54024 2388 54076 2440
rect 54208 2388 54260 2440
rect 55036 2388 55088 2440
rect 57520 2388 57572 2440
rect 59268 2388 59320 2440
rect 60004 2388 60056 2440
rect 62672 2388 62724 2440
rect 65248 2388 65300 2440
rect 71320 2431 71372 2440
rect 71320 2397 71329 2431
rect 71329 2397 71363 2431
rect 71363 2397 71372 2431
rect 71320 2388 71372 2397
rect 73160 2388 73212 2440
rect 73528 2431 73580 2440
rect 73528 2397 73537 2431
rect 73537 2397 73571 2431
rect 73571 2397 73580 2431
rect 73528 2388 73580 2397
rect 73804 2431 73856 2440
rect 73804 2397 73813 2431
rect 73813 2397 73847 2431
rect 73847 2397 73856 2431
rect 73804 2388 73856 2397
rect 76472 2431 76524 2440
rect 76472 2397 76481 2431
rect 76481 2397 76515 2431
rect 76515 2397 76524 2431
rect 76472 2388 76524 2397
rect 76748 2431 76800 2440
rect 76748 2397 76757 2431
rect 76757 2397 76791 2431
rect 76791 2397 76800 2431
rect 76748 2388 76800 2397
rect 77944 2431 77996 2440
rect 77944 2397 77953 2431
rect 77953 2397 77987 2431
rect 77987 2397 77996 2431
rect 77944 2388 77996 2397
rect 78220 2499 78272 2508
rect 78220 2465 78229 2499
rect 78229 2465 78263 2499
rect 78263 2465 78272 2499
rect 78220 2456 78272 2465
rect 79416 2431 79468 2440
rect 79416 2397 79425 2431
rect 79425 2397 79459 2431
rect 79459 2397 79468 2431
rect 79416 2388 79468 2397
rect 79968 2388 80020 2440
rect 27252 2252 27304 2304
rect 35624 2320 35676 2372
rect 36452 2320 36504 2372
rect 27896 2252 27948 2304
rect 28724 2295 28776 2304
rect 28724 2261 28733 2295
rect 28733 2261 28767 2295
rect 28767 2261 28776 2295
rect 28724 2252 28776 2261
rect 32312 2252 32364 2304
rect 33048 2295 33100 2304
rect 33048 2261 33057 2295
rect 33057 2261 33091 2295
rect 33091 2261 33100 2295
rect 33048 2252 33100 2261
rect 36728 2252 36780 2304
rect 37096 2320 37148 2372
rect 37280 2363 37332 2372
rect 37280 2329 37289 2363
rect 37289 2329 37323 2363
rect 37323 2329 37332 2363
rect 37280 2320 37332 2329
rect 40040 2320 40092 2372
rect 82360 2431 82412 2440
rect 82360 2397 82369 2431
rect 82369 2397 82403 2431
rect 82403 2397 82412 2431
rect 82360 2388 82412 2397
rect 37740 2252 37792 2304
rect 38200 2295 38252 2304
rect 38200 2261 38209 2295
rect 38209 2261 38243 2295
rect 38243 2261 38252 2295
rect 38200 2252 38252 2261
rect 53840 2252 53892 2304
rect 54852 2295 54904 2304
rect 54852 2261 54861 2295
rect 54861 2261 54895 2295
rect 54895 2261 54904 2295
rect 54852 2252 54904 2261
rect 55680 2295 55732 2304
rect 55680 2261 55689 2295
rect 55689 2261 55723 2295
rect 55723 2261 55732 2295
rect 55680 2252 55732 2261
rect 57796 2295 57848 2304
rect 57796 2261 57805 2295
rect 57805 2261 57839 2295
rect 57839 2261 57848 2295
rect 57796 2252 57848 2261
rect 59360 2295 59412 2304
rect 59360 2261 59369 2295
rect 59369 2261 59403 2295
rect 59403 2261 59412 2295
rect 59360 2252 59412 2261
rect 62948 2295 63000 2304
rect 62948 2261 62957 2295
rect 62957 2261 62991 2295
rect 62991 2261 63000 2295
rect 62948 2252 63000 2261
rect 65616 2252 65668 2304
rect 66628 2295 66680 2304
rect 66628 2261 66637 2295
rect 66637 2261 66671 2295
rect 66671 2261 66680 2295
rect 66628 2252 66680 2261
rect 83004 2320 83056 2372
rect 87972 2456 88024 2508
rect 96344 2456 96396 2508
rect 83740 2363 83792 2372
rect 83740 2329 83749 2363
rect 83749 2329 83783 2363
rect 83783 2329 83792 2363
rect 83740 2320 83792 2329
rect 84016 2320 84068 2372
rect 85396 2363 85448 2372
rect 85396 2329 85405 2363
rect 85405 2329 85439 2363
rect 85439 2329 85448 2363
rect 85396 2320 85448 2329
rect 88340 2431 88392 2440
rect 88340 2397 88349 2431
rect 88349 2397 88383 2431
rect 88383 2397 88392 2431
rect 88340 2388 88392 2397
rect 89904 2388 89956 2440
rect 91100 2388 91152 2440
rect 92756 2388 92808 2440
rect 93676 2431 93728 2440
rect 93676 2397 93685 2431
rect 93685 2397 93719 2431
rect 93719 2397 93728 2431
rect 93676 2388 93728 2397
rect 94412 2431 94464 2440
rect 94412 2397 94421 2431
rect 94421 2397 94455 2431
rect 94455 2397 94464 2431
rect 94412 2388 94464 2397
rect 95424 2388 95476 2440
rect 96252 2388 96304 2440
rect 96896 2524 96948 2576
rect 97356 2567 97408 2576
rect 97356 2533 97365 2567
rect 97365 2533 97399 2567
rect 97399 2533 97408 2567
rect 97356 2524 97408 2533
rect 97448 2456 97500 2508
rect 97632 2431 97684 2440
rect 97632 2397 97641 2431
rect 97641 2397 97675 2431
rect 97675 2397 97684 2431
rect 97632 2388 97684 2397
rect 97908 2431 97960 2474
rect 97908 2422 97917 2431
rect 97917 2422 97951 2431
rect 97951 2422 97960 2431
rect 98092 2456 98144 2508
rect 98552 2635 98604 2644
rect 98552 2601 98561 2635
rect 98561 2601 98595 2635
rect 98595 2601 98604 2635
rect 98552 2592 98604 2601
rect 98828 2592 98880 2644
rect 98644 2524 98696 2576
rect 103336 2524 103388 2576
rect 104164 2524 104216 2576
rect 105268 2635 105320 2644
rect 105268 2601 105277 2635
rect 105277 2601 105311 2635
rect 105311 2601 105320 2635
rect 105268 2592 105320 2601
rect 107660 2592 107712 2644
rect 149152 2592 149204 2644
rect 143724 2567 143776 2576
rect 98460 2456 98512 2508
rect 99748 2456 99800 2508
rect 103428 2499 103480 2508
rect 103428 2465 103437 2499
rect 103437 2465 103471 2499
rect 103471 2465 103480 2499
rect 103428 2456 103480 2465
rect 104348 2499 104400 2508
rect 104348 2465 104357 2499
rect 104357 2465 104391 2499
rect 104391 2465 104400 2499
rect 104348 2456 104400 2465
rect 107476 2456 107528 2508
rect 107936 2456 107988 2508
rect 109040 2499 109092 2508
rect 109040 2465 109049 2499
rect 109049 2465 109083 2499
rect 109083 2465 109092 2499
rect 109040 2456 109092 2465
rect 139124 2499 139176 2508
rect 139124 2465 139133 2499
rect 139133 2465 139167 2499
rect 139167 2465 139176 2499
rect 139124 2456 139176 2465
rect 141148 2456 141200 2508
rect 143724 2533 143733 2567
rect 143733 2533 143767 2567
rect 143767 2533 143776 2567
rect 143724 2524 143776 2533
rect 145656 2524 145708 2576
rect 148876 2567 148928 2576
rect 148876 2533 148885 2567
rect 148885 2533 148919 2567
rect 148919 2533 148928 2567
rect 148876 2524 148928 2533
rect 143172 2456 143224 2508
rect 144460 2456 144512 2508
rect 146208 2456 146260 2508
rect 149152 2499 149204 2508
rect 149152 2465 149161 2499
rect 149161 2465 149195 2499
rect 149195 2465 149204 2499
rect 149152 2456 149204 2465
rect 150992 2456 151044 2508
rect 152372 2499 152424 2508
rect 152372 2465 152381 2499
rect 152381 2465 152415 2499
rect 152415 2465 152424 2499
rect 152372 2456 152424 2465
rect 156880 2592 156932 2644
rect 156972 2592 157024 2644
rect 157156 2592 157208 2644
rect 157340 2592 157392 2644
rect 160100 2592 160152 2644
rect 160744 2592 160796 2644
rect 161388 2592 161440 2644
rect 176660 2592 176712 2644
rect 155132 2524 155184 2576
rect 159456 2524 159508 2576
rect 156880 2456 156932 2508
rect 87604 2295 87656 2304
rect 87604 2261 87613 2295
rect 87613 2261 87647 2295
rect 87647 2261 87656 2295
rect 87604 2252 87656 2261
rect 89536 2320 89588 2372
rect 89260 2252 89312 2304
rect 91008 2320 91060 2372
rect 90272 2252 90324 2304
rect 90824 2295 90876 2304
rect 90824 2261 90833 2295
rect 90833 2261 90867 2295
rect 90867 2261 90876 2295
rect 90824 2252 90876 2261
rect 91744 2295 91796 2304
rect 91744 2261 91753 2295
rect 91753 2261 91787 2295
rect 91787 2261 91796 2295
rect 91744 2252 91796 2261
rect 93032 2295 93084 2304
rect 93032 2261 93041 2295
rect 93041 2261 93075 2295
rect 93075 2261 93084 2295
rect 93032 2252 93084 2261
rect 93860 2295 93912 2304
rect 93860 2261 93869 2295
rect 93869 2261 93903 2295
rect 93903 2261 93912 2295
rect 93860 2252 93912 2261
rect 94596 2295 94648 2304
rect 94596 2261 94605 2295
rect 94605 2261 94639 2295
rect 94639 2261 94648 2295
rect 94596 2252 94648 2261
rect 95332 2295 95384 2304
rect 95332 2261 95341 2295
rect 95341 2261 95375 2295
rect 95375 2261 95384 2295
rect 95332 2252 95384 2261
rect 96068 2295 96120 2304
rect 96068 2261 96077 2295
rect 96077 2261 96111 2295
rect 96111 2261 96120 2295
rect 96068 2252 96120 2261
rect 99012 2295 99064 2304
rect 99012 2261 99021 2295
rect 99021 2261 99055 2295
rect 99055 2261 99064 2295
rect 99012 2252 99064 2261
rect 99196 2320 99248 2372
rect 104624 2431 104676 2440
rect 104624 2397 104633 2431
rect 104633 2397 104667 2431
rect 104667 2397 104676 2431
rect 104624 2388 104676 2397
rect 122012 2388 122064 2440
rect 124496 2388 124548 2440
rect 126244 2388 126296 2440
rect 127900 2388 127952 2440
rect 128636 2388 128688 2440
rect 129648 2388 129700 2440
rect 131672 2388 131724 2440
rect 133328 2388 133380 2440
rect 133604 2388 133656 2440
rect 134340 2388 134392 2440
rect 101220 2363 101272 2372
rect 101220 2329 101229 2363
rect 101229 2329 101263 2363
rect 101263 2329 101272 2363
rect 101220 2320 101272 2329
rect 107292 2320 107344 2372
rect 109316 2320 109368 2372
rect 133236 2320 133288 2372
rect 142804 2388 142856 2440
rect 144184 2388 144236 2440
rect 144276 2431 144328 2440
rect 144276 2397 144285 2431
rect 144285 2397 144319 2431
rect 144319 2397 144328 2431
rect 144276 2388 144328 2397
rect 147772 2388 147824 2440
rect 149428 2431 149480 2440
rect 149428 2397 149437 2431
rect 149437 2397 149471 2431
rect 149471 2397 149480 2431
rect 149428 2388 149480 2397
rect 155224 2431 155276 2440
rect 155224 2397 155233 2431
rect 155233 2397 155267 2431
rect 155267 2397 155276 2431
rect 155224 2388 155276 2397
rect 156604 2388 156656 2440
rect 157340 2431 157392 2440
rect 157340 2397 157349 2431
rect 157349 2397 157383 2431
rect 157383 2397 157392 2431
rect 157340 2388 157392 2397
rect 157708 2431 157760 2440
rect 157708 2397 157717 2431
rect 157717 2397 157751 2431
rect 157751 2397 157760 2431
rect 157708 2388 157760 2397
rect 157800 2388 157852 2440
rect 158628 2431 158680 2440
rect 158628 2397 158637 2431
rect 158637 2397 158671 2431
rect 158671 2397 158680 2431
rect 158628 2388 158680 2397
rect 159916 2431 159968 2440
rect 159916 2397 159925 2431
rect 159925 2397 159959 2431
rect 159959 2397 159968 2431
rect 159916 2388 159968 2397
rect 160008 2388 160060 2440
rect 160376 2431 160428 2440
rect 160376 2397 160385 2431
rect 160385 2397 160419 2431
rect 160419 2397 160428 2431
rect 160376 2388 160428 2397
rect 103520 2252 103572 2304
rect 104624 2252 104676 2304
rect 108396 2252 108448 2304
rect 122656 2295 122708 2304
rect 122656 2261 122665 2295
rect 122665 2261 122699 2295
rect 122699 2261 122708 2295
rect 122656 2252 122708 2261
rect 124772 2295 124824 2304
rect 124772 2261 124781 2295
rect 124781 2261 124815 2295
rect 124815 2261 124824 2295
rect 124772 2252 124824 2261
rect 126336 2295 126388 2304
rect 126336 2261 126345 2295
rect 126345 2261 126379 2295
rect 126379 2261 126388 2295
rect 126336 2252 126388 2261
rect 127808 2295 127860 2304
rect 127808 2261 127817 2295
rect 127817 2261 127851 2295
rect 127851 2261 127860 2295
rect 127808 2252 127860 2261
rect 128360 2252 128412 2304
rect 130016 2295 130068 2304
rect 130016 2261 130025 2295
rect 130025 2261 130059 2295
rect 130059 2261 130068 2295
rect 130016 2252 130068 2261
rect 131580 2295 131632 2304
rect 131580 2261 131589 2295
rect 131589 2261 131623 2295
rect 131623 2261 131632 2295
rect 131580 2252 131632 2261
rect 132960 2295 133012 2304
rect 132960 2261 132969 2295
rect 132969 2261 133003 2295
rect 133003 2261 133012 2295
rect 132960 2252 133012 2261
rect 133696 2295 133748 2304
rect 133696 2261 133705 2295
rect 133705 2261 133739 2295
rect 133739 2261 133748 2295
rect 133696 2252 133748 2261
rect 134432 2295 134484 2304
rect 134432 2261 134441 2295
rect 134441 2261 134475 2295
rect 134475 2261 134484 2295
rect 134432 2252 134484 2261
rect 134984 2295 135036 2304
rect 134984 2261 134993 2295
rect 134993 2261 135027 2295
rect 135027 2261 135036 2295
rect 134984 2252 135036 2261
rect 139952 2320 140004 2372
rect 155776 2320 155828 2372
rect 156880 2320 156932 2372
rect 141332 2252 141384 2304
rect 148968 2252 149020 2304
rect 156328 2252 156380 2304
rect 156512 2252 156564 2304
rect 158168 2320 158220 2372
rect 158536 2320 158588 2372
rect 162308 2388 162360 2440
rect 163964 2388 164016 2440
rect 164424 2431 164476 2440
rect 164424 2397 164433 2431
rect 164433 2397 164467 2431
rect 164467 2397 164476 2431
rect 164424 2388 164476 2397
rect 165620 2388 165672 2440
rect 165896 2431 165948 2440
rect 165896 2397 165905 2431
rect 165905 2397 165939 2431
rect 165939 2397 165948 2431
rect 165896 2388 165948 2397
rect 167460 2388 167512 2440
rect 167736 2431 167788 2440
rect 167736 2397 167745 2431
rect 167745 2397 167779 2431
rect 167779 2397 167788 2431
rect 167736 2388 167788 2397
rect 167828 2431 167880 2440
rect 167828 2397 167837 2431
rect 167837 2397 167871 2431
rect 167871 2397 167880 2431
rect 167828 2388 167880 2397
rect 176660 2431 176712 2440
rect 176660 2397 176669 2431
rect 176669 2397 176703 2431
rect 176703 2397 176712 2431
rect 176660 2388 176712 2397
rect 176936 2431 176988 2440
rect 176936 2397 176945 2431
rect 176945 2397 176979 2431
rect 176979 2397 176988 2431
rect 176936 2388 176988 2397
rect 179604 2431 179656 2440
rect 179604 2397 179613 2431
rect 179613 2397 179647 2431
rect 179647 2397 179656 2431
rect 179604 2388 179656 2397
rect 186964 2431 187016 2440
rect 186964 2397 186973 2431
rect 186973 2397 187007 2431
rect 187007 2397 187016 2431
rect 186964 2388 187016 2397
rect 190460 2592 190512 2644
rect 191840 2592 191892 2644
rect 202880 2592 202932 2644
rect 202604 2456 202656 2508
rect 213184 2592 213236 2644
rect 221924 2592 221976 2644
rect 224960 2592 225012 2644
rect 226248 2592 226300 2644
rect 227996 2592 228048 2644
rect 231676 2592 231728 2644
rect 236000 2635 236052 2644
rect 236000 2601 236009 2635
rect 236009 2601 236043 2635
rect 236043 2601 236052 2635
rect 236000 2592 236052 2601
rect 236736 2592 236788 2644
rect 242808 2592 242860 2644
rect 258080 2592 258132 2644
rect 266452 2592 266504 2644
rect 268384 2592 268436 2644
rect 210148 2524 210200 2576
rect 210792 2524 210844 2576
rect 213736 2524 213788 2576
rect 205088 2499 205140 2508
rect 205088 2465 205097 2499
rect 205097 2465 205131 2499
rect 205131 2465 205140 2499
rect 205088 2456 205140 2465
rect 205364 2499 205416 2508
rect 205364 2465 205373 2499
rect 205373 2465 205407 2499
rect 205407 2465 205416 2499
rect 205364 2456 205416 2465
rect 208124 2456 208176 2508
rect 189724 2388 189776 2440
rect 190368 2431 190420 2440
rect 190368 2397 190377 2431
rect 190377 2397 190411 2431
rect 190411 2397 190420 2431
rect 190368 2388 190420 2397
rect 191380 2388 191432 2440
rect 192392 2388 192444 2440
rect 195704 2388 195756 2440
rect 196256 2431 196308 2440
rect 196256 2397 196265 2431
rect 196265 2397 196299 2431
rect 196299 2397 196308 2431
rect 196256 2388 196308 2397
rect 197176 2431 197228 2440
rect 197176 2397 197185 2431
rect 197185 2397 197219 2431
rect 197219 2397 197228 2431
rect 197176 2388 197228 2397
rect 197268 2431 197320 2440
rect 197268 2397 197277 2431
rect 197277 2397 197311 2431
rect 197311 2397 197320 2431
rect 197268 2388 197320 2397
rect 199200 2388 199252 2440
rect 200856 2388 200908 2440
rect 201224 2431 201276 2440
rect 201224 2397 201233 2431
rect 201233 2397 201267 2431
rect 201267 2397 201276 2431
rect 201224 2388 201276 2397
rect 201316 2388 201368 2440
rect 209964 2388 210016 2440
rect 211068 2431 211120 2440
rect 211068 2397 211102 2431
rect 211102 2397 211120 2431
rect 211068 2388 211120 2397
rect 211252 2431 211304 2440
rect 211252 2397 211261 2431
rect 211261 2397 211295 2431
rect 211295 2397 211304 2431
rect 211252 2388 211304 2397
rect 216128 2456 216180 2508
rect 214104 2388 214156 2440
rect 218612 2499 218664 2508
rect 218612 2465 218621 2499
rect 218621 2465 218655 2499
rect 218655 2465 218664 2499
rect 218612 2456 218664 2465
rect 221004 2499 221056 2508
rect 221004 2465 221013 2499
rect 221013 2465 221047 2499
rect 221047 2465 221056 2499
rect 221004 2456 221056 2465
rect 255320 2524 255372 2576
rect 269028 2524 269080 2576
rect 221924 2499 221976 2508
rect 221924 2465 221933 2499
rect 221933 2465 221967 2499
rect 221967 2465 221976 2499
rect 221924 2456 221976 2465
rect 161664 2320 161716 2372
rect 167552 2320 167604 2372
rect 168196 2320 168248 2372
rect 174728 2320 174780 2372
rect 157432 2252 157484 2304
rect 160928 2295 160980 2304
rect 160928 2261 160937 2295
rect 160937 2261 160971 2295
rect 160971 2261 160980 2295
rect 160928 2252 160980 2261
rect 161756 2295 161808 2304
rect 161756 2261 161765 2295
rect 161765 2261 161799 2295
rect 161799 2261 161808 2295
rect 161756 2252 161808 2261
rect 162124 2252 162176 2304
rect 162492 2252 162544 2304
rect 163872 2295 163924 2304
rect 163872 2261 163881 2295
rect 163881 2261 163915 2295
rect 163915 2261 163924 2295
rect 163872 2252 163924 2261
rect 164240 2252 164292 2304
rect 165344 2295 165396 2304
rect 165344 2261 165353 2295
rect 165353 2261 165387 2295
rect 165387 2261 165396 2295
rect 165344 2252 165396 2261
rect 166080 2295 166132 2304
rect 166080 2261 166089 2295
rect 166089 2261 166123 2295
rect 166123 2261 166132 2295
rect 166080 2252 166132 2261
rect 166816 2295 166868 2304
rect 166816 2261 166825 2295
rect 166825 2261 166859 2295
rect 166859 2261 166868 2295
rect 166816 2252 166868 2261
rect 168012 2295 168064 2304
rect 168012 2261 168021 2295
rect 168021 2261 168055 2295
rect 168055 2261 168064 2295
rect 168012 2252 168064 2261
rect 173808 2252 173860 2304
rect 183560 2252 183612 2304
rect 191288 2295 191340 2304
rect 191288 2261 191297 2295
rect 191297 2261 191331 2295
rect 191331 2261 191340 2295
rect 191288 2252 191340 2261
rect 194692 2252 194744 2304
rect 195980 2252 196032 2304
rect 197452 2295 197504 2304
rect 197452 2261 197461 2295
rect 197461 2261 197495 2295
rect 197495 2261 197504 2295
rect 197452 2252 197504 2261
rect 198556 2295 198608 2304
rect 198556 2261 198565 2295
rect 198565 2261 198599 2295
rect 198599 2261 198608 2295
rect 198556 2252 198608 2261
rect 199936 2295 199988 2304
rect 199936 2261 199945 2295
rect 199945 2261 199979 2295
rect 199979 2261 199988 2295
rect 199936 2252 199988 2261
rect 201408 2295 201460 2304
rect 201408 2261 201417 2295
rect 201417 2261 201451 2295
rect 201451 2261 201460 2295
rect 201408 2252 201460 2261
rect 204260 2295 204312 2304
rect 204260 2261 204269 2295
rect 204269 2261 204303 2295
rect 204303 2261 204312 2295
rect 204260 2252 204312 2261
rect 205364 2252 205416 2304
rect 207020 2295 207072 2304
rect 207020 2261 207029 2295
rect 207029 2261 207063 2295
rect 207063 2261 207072 2295
rect 207020 2252 207072 2261
rect 207112 2252 207164 2304
rect 213184 2252 213236 2304
rect 213276 2252 213328 2304
rect 218060 2388 218112 2440
rect 219072 2388 219124 2440
rect 220728 2320 220780 2372
rect 216404 2252 216456 2304
rect 218152 2252 218204 2304
rect 219808 2252 219860 2304
rect 221372 2388 221424 2440
rect 223028 2431 223080 2440
rect 223028 2397 223037 2431
rect 223037 2397 223071 2431
rect 223071 2397 223080 2431
rect 223028 2388 223080 2397
rect 223580 2456 223632 2508
rect 223672 2388 223724 2440
rect 258724 2456 258776 2508
rect 221648 2320 221700 2372
rect 225328 2431 225380 2440
rect 225328 2397 225337 2431
rect 225337 2397 225371 2431
rect 225371 2397 225380 2431
rect 225328 2388 225380 2397
rect 226156 2388 226208 2440
rect 226248 2431 226300 2440
rect 226248 2397 226257 2431
rect 226257 2397 226291 2431
rect 226291 2397 226300 2431
rect 226248 2388 226300 2397
rect 226984 2431 227036 2440
rect 226984 2397 226993 2431
rect 226993 2397 227027 2431
rect 227027 2397 227036 2431
rect 226984 2388 227036 2397
rect 227628 2388 227680 2440
rect 228364 2388 228416 2440
rect 228824 2431 228876 2440
rect 228824 2397 228833 2431
rect 228833 2397 228867 2431
rect 228867 2397 228876 2431
rect 228824 2388 228876 2397
rect 231768 2388 231820 2440
rect 231860 2431 231912 2440
rect 231860 2397 231869 2431
rect 231869 2397 231903 2431
rect 231903 2397 231912 2431
rect 231860 2388 231912 2397
rect 232596 2431 232648 2440
rect 232596 2397 232605 2431
rect 232605 2397 232639 2431
rect 232639 2397 232648 2431
rect 232596 2388 232648 2397
rect 236092 2388 236144 2440
rect 236552 2431 236604 2440
rect 236552 2397 236561 2431
rect 236561 2397 236595 2431
rect 236595 2397 236604 2431
rect 236552 2388 236604 2397
rect 243452 2431 243504 2440
rect 243452 2397 243461 2431
rect 243461 2397 243495 2431
rect 243495 2397 243504 2431
rect 243452 2388 243504 2397
rect 246396 2431 246448 2440
rect 246396 2397 246405 2431
rect 246405 2397 246439 2431
rect 246439 2397 246448 2431
rect 246396 2388 246448 2397
rect 256700 2431 256752 2440
rect 256700 2397 256709 2431
rect 256709 2397 256743 2431
rect 256743 2397 256752 2431
rect 256700 2388 256752 2397
rect 256976 2431 257028 2440
rect 256976 2397 256985 2431
rect 256985 2397 257019 2431
rect 257019 2397 257028 2431
rect 256976 2388 257028 2397
rect 259092 2431 259144 2440
rect 259092 2397 259101 2431
rect 259101 2397 259135 2431
rect 259135 2397 259144 2431
rect 259092 2388 259144 2397
rect 261576 2431 261628 2440
rect 261576 2397 261585 2431
rect 261585 2397 261619 2431
rect 261619 2397 261628 2431
rect 261576 2388 261628 2397
rect 263968 2431 264020 2440
rect 263968 2397 263977 2431
rect 263977 2397 264011 2431
rect 264011 2397 264020 2431
rect 263968 2388 264020 2397
rect 264244 2388 264296 2440
rect 267280 2431 267332 2442
rect 267280 2397 267289 2431
rect 267289 2397 267323 2431
rect 267323 2397 267332 2431
rect 267280 2390 267332 2397
rect 224040 2320 224092 2372
rect 221372 2252 221424 2304
rect 222476 2252 222528 2304
rect 222568 2295 222620 2304
rect 222568 2261 222577 2295
rect 222577 2261 222611 2295
rect 222611 2261 222620 2295
rect 222568 2252 222620 2261
rect 223764 2252 223816 2304
rect 224224 2252 224276 2304
rect 227812 2320 227864 2372
rect 237196 2320 237248 2372
rect 258080 2363 258132 2372
rect 258080 2329 258089 2363
rect 258089 2329 258123 2363
rect 258123 2329 258132 2363
rect 258080 2320 258132 2329
rect 264428 2320 264480 2372
rect 268568 2431 268620 2440
rect 268568 2397 268577 2431
rect 268577 2397 268611 2431
rect 268611 2397 268620 2431
rect 268568 2388 268620 2397
rect 270132 2456 270184 2508
rect 269212 2431 269264 2440
rect 269212 2397 269221 2431
rect 269221 2397 269255 2431
rect 269255 2397 269264 2431
rect 269212 2388 269264 2397
rect 269672 2388 269724 2440
rect 270500 2388 270552 2440
rect 225604 2252 225656 2304
rect 226708 2252 226760 2304
rect 227168 2252 227220 2304
rect 228456 2252 228508 2304
rect 231308 2295 231360 2304
rect 231308 2261 231317 2295
rect 231317 2261 231351 2295
rect 231351 2261 231360 2295
rect 231308 2252 231360 2261
rect 232044 2295 232096 2304
rect 232044 2261 232053 2295
rect 232053 2261 232087 2295
rect 232087 2261 232096 2295
rect 232044 2252 232096 2261
rect 232780 2295 232832 2304
rect 232780 2261 232789 2295
rect 232789 2261 232823 2295
rect 232823 2261 232832 2295
rect 232780 2252 232832 2261
rect 236736 2295 236788 2304
rect 236736 2261 236745 2295
rect 236745 2261 236779 2295
rect 236779 2261 236788 2295
rect 236736 2252 236788 2261
rect 244280 2252 244332 2304
rect 255412 2252 255464 2304
rect 257712 2252 257764 2304
rect 257896 2252 257948 2304
rect 259920 2295 259972 2304
rect 259920 2261 259929 2295
rect 259929 2261 259963 2295
rect 259963 2261 259972 2295
rect 259920 2252 259972 2261
rect 261852 2252 261904 2304
rect 264980 2295 265032 2304
rect 264980 2261 264989 2295
rect 264989 2261 265023 2295
rect 265023 2261 265032 2295
rect 264980 2252 265032 2261
rect 267556 2252 267608 2304
rect 268844 2320 268896 2372
rect 268200 2252 268252 2304
rect 269948 2252 270000 2304
rect 270040 2295 270092 2304
rect 270040 2261 270049 2295
rect 270049 2261 270083 2295
rect 270083 2261 270092 2295
rect 270040 2252 270092 2261
rect 270776 2295 270828 2304
rect 270776 2261 270785 2295
rect 270785 2261 270819 2295
rect 270819 2261 270828 2295
rect 270776 2252 270828 2261
rect 68546 2150 68598 2202
rect 68610 2150 68662 2202
rect 68674 2150 68726 2202
rect 68738 2150 68790 2202
rect 68802 2150 68854 2202
rect 136143 2150 136195 2202
rect 136207 2150 136259 2202
rect 136271 2150 136323 2202
rect 136335 2150 136387 2202
rect 136399 2150 136451 2202
rect 203740 2150 203792 2202
rect 203804 2150 203856 2202
rect 203868 2150 203920 2202
rect 203932 2150 203984 2202
rect 203996 2150 204048 2202
rect 271337 2150 271389 2202
rect 271401 2150 271453 2202
rect 271465 2150 271517 2202
rect 271529 2150 271581 2202
rect 271593 2150 271645 2202
rect 9220 2023 9272 2032
rect 9220 1989 9229 2023
rect 9229 1989 9263 2023
rect 9263 1989 9272 2023
rect 9220 1980 9272 1989
rect 17132 2023 17184 2032
rect 17132 1989 17141 2023
rect 17141 1989 17175 2023
rect 17175 1989 17184 2023
rect 17132 1980 17184 1989
rect 23848 2091 23900 2100
rect 23848 2057 23857 2091
rect 23857 2057 23891 2091
rect 23891 2057 23900 2091
rect 23848 2048 23900 2057
rect 26332 2091 26384 2100
rect 26332 2057 26341 2091
rect 26341 2057 26375 2091
rect 26375 2057 26384 2091
rect 26332 2048 26384 2057
rect 25136 1980 25188 2032
rect 25596 1980 25648 2032
rect 26424 1980 26476 2032
rect 2596 1955 2648 1964
rect 2596 1921 2605 1955
rect 2605 1921 2639 1955
rect 2639 1921 2648 1955
rect 2596 1912 2648 1921
rect 4804 1955 4856 1964
rect 4804 1921 4813 1955
rect 4813 1921 4847 1955
rect 4847 1921 4856 1955
rect 4804 1912 4856 1921
rect 6828 1955 6880 1964
rect 6828 1921 6837 1955
rect 6837 1921 6871 1955
rect 6871 1921 6880 1955
rect 6828 1912 6880 1921
rect 7564 1955 7616 1964
rect 7564 1921 7573 1955
rect 7573 1921 7607 1955
rect 7607 1921 7616 1955
rect 7564 1912 7616 1921
rect 9036 1955 9088 1964
rect 9036 1921 9045 1955
rect 9045 1921 9079 1955
rect 9079 1921 9088 1955
rect 9036 1912 9088 1921
rect 14372 1955 14424 1964
rect 14372 1921 14381 1955
rect 14381 1921 14415 1955
rect 14415 1921 14424 1955
rect 14372 1912 14424 1921
rect 15660 1955 15712 1964
rect 15660 1921 15669 1955
rect 15669 1921 15703 1955
rect 15703 1921 15712 1955
rect 15660 1912 15712 1921
rect 15844 1955 15896 1964
rect 15844 1921 15853 1955
rect 15853 1921 15887 1955
rect 15887 1921 15896 1955
rect 15844 1912 15896 1921
rect 16580 1912 16632 1964
rect 23572 1955 23624 1964
rect 23572 1921 23581 1955
rect 23581 1921 23615 1955
rect 23615 1921 23624 1955
rect 23572 1912 23624 1921
rect 2320 1887 2372 1896
rect 2320 1853 2329 1887
rect 2329 1853 2363 1887
rect 2363 1853 2372 1887
rect 2320 1844 2372 1853
rect 4528 1887 4580 1896
rect 4528 1853 4537 1887
rect 4537 1853 4571 1887
rect 4571 1853 4580 1887
rect 4528 1844 4580 1853
rect 14096 1887 14148 1896
rect 14096 1853 14105 1887
rect 14105 1853 14139 1887
rect 14139 1853 14148 1887
rect 14096 1844 14148 1853
rect 23940 1912 23992 1964
rect 24952 1912 25004 1964
rect 25688 1912 25740 1964
rect 27712 1980 27764 2032
rect 27896 1980 27948 2032
rect 28448 1912 28500 1964
rect 29552 1955 29604 1964
rect 29552 1921 29561 1955
rect 29561 1921 29595 1955
rect 29595 1921 29604 1955
rect 29552 1912 29604 1921
rect 30380 1955 30432 1964
rect 30380 1921 30389 1955
rect 30389 1921 30423 1955
rect 30423 1921 30432 1955
rect 30380 1912 30432 1921
rect 31208 1912 31260 1964
rect 33048 1980 33100 2032
rect 35532 2023 35584 2032
rect 35532 1989 35541 2023
rect 35541 1989 35575 2023
rect 35575 1989 35584 2023
rect 35532 1980 35584 1989
rect 35808 2023 35860 2032
rect 35808 1989 35817 2023
rect 35817 1989 35851 2023
rect 35851 1989 35860 2023
rect 35808 1980 35860 1989
rect 36360 1980 36412 2032
rect 36636 2023 36688 2032
rect 36636 1989 36645 2023
rect 36645 1989 36679 2023
rect 36679 1989 36688 2023
rect 36636 1980 36688 1989
rect 37280 1980 37332 2032
rect 25044 1844 25096 1896
rect 25136 1844 25188 1896
rect 31024 1844 31076 1896
rect 32496 1955 32548 1964
rect 32496 1921 32505 1955
rect 32505 1921 32539 1955
rect 32539 1921 32548 1955
rect 32496 1912 32548 1921
rect 38660 1980 38712 2032
rect 39304 2023 39356 2032
rect 39304 1989 39313 2023
rect 39313 1989 39347 2023
rect 39347 1989 39356 2023
rect 39304 1980 39356 1989
rect 39764 2023 39816 2032
rect 39764 1989 39773 2023
rect 39773 1989 39807 2023
rect 39807 1989 39816 2023
rect 39764 1980 39816 1989
rect 38108 1955 38160 1964
rect 38108 1921 38117 1955
rect 38117 1921 38151 1955
rect 38151 1921 38160 1955
rect 38108 1912 38160 1921
rect 38292 1912 38344 1964
rect 40040 1980 40092 2032
rect 40132 2023 40184 2032
rect 40132 1989 40141 2023
rect 40141 1989 40175 2023
rect 40175 1989 40184 2023
rect 40132 1980 40184 1989
rect 54208 2023 54260 2032
rect 54208 1989 54217 2023
rect 54217 1989 54251 2023
rect 54251 1989 54260 2023
rect 54208 1980 54260 1989
rect 55036 2023 55088 2032
rect 55036 1989 55045 2023
rect 55045 1989 55079 2023
rect 55079 1989 55088 2023
rect 55036 1980 55088 1989
rect 57520 2091 57572 2100
rect 57520 2057 57529 2091
rect 57529 2057 57563 2091
rect 57563 2057 57572 2091
rect 57520 2048 57572 2057
rect 58532 2091 58584 2100
rect 58532 2057 58541 2091
rect 58541 2057 58575 2091
rect 58575 2057 58584 2091
rect 58532 2048 58584 2057
rect 59268 2091 59320 2100
rect 59268 2057 59277 2091
rect 59277 2057 59311 2091
rect 59311 2057 59320 2091
rect 59268 2048 59320 2057
rect 62672 2091 62724 2100
rect 62672 2057 62681 2091
rect 62681 2057 62715 2091
rect 62715 2057 62724 2091
rect 62672 2048 62724 2057
rect 65248 2091 65300 2100
rect 65248 2057 65257 2091
rect 65257 2057 65291 2091
rect 65291 2057 65300 2091
rect 65248 2048 65300 2057
rect 39948 1912 40000 1964
rect 45468 1955 45520 1964
rect 45468 1921 45477 1955
rect 45477 1921 45511 1955
rect 45511 1921 45520 1955
rect 45468 1912 45520 1921
rect 50620 1955 50672 1964
rect 50620 1921 50629 1955
rect 50629 1921 50663 1955
rect 50663 1921 50672 1955
rect 50620 1912 50672 1921
rect 52920 1955 52972 1964
rect 52920 1921 52929 1955
rect 52929 1921 52963 1955
rect 52963 1921 52972 1955
rect 52920 1912 52972 1921
rect 54024 1955 54076 1964
rect 54024 1921 54033 1955
rect 54033 1921 54067 1955
rect 54067 1921 54076 1955
rect 54024 1912 54076 1921
rect 55404 1912 55456 1964
rect 56324 1955 56376 1964
rect 56324 1921 56333 1955
rect 56333 1921 56367 1955
rect 56367 1921 56376 1955
rect 56324 1912 56376 1921
rect 57152 1955 57204 1964
rect 57152 1921 57161 1955
rect 57161 1921 57195 1955
rect 57195 1921 57204 1955
rect 57152 1912 57204 1921
rect 37188 1844 37240 1896
rect 53472 1844 53524 1896
rect 54392 1844 54444 1896
rect 58532 1844 58584 1896
rect 58900 1887 58952 1896
rect 58900 1853 58909 1887
rect 58909 1853 58943 1887
rect 58943 1853 58952 1887
rect 58900 1844 58952 1853
rect 59820 1955 59872 1964
rect 59820 1921 59829 1955
rect 59829 1921 59863 1955
rect 59863 1921 59872 1955
rect 59820 1912 59872 1921
rect 59912 1844 59964 1896
rect 60648 1955 60700 1964
rect 60648 1921 60657 1955
rect 60657 1921 60691 1955
rect 60691 1921 60700 1955
rect 60648 1912 60700 1921
rect 61568 1955 61620 1964
rect 61568 1921 61577 1955
rect 61577 1921 61611 1955
rect 61611 1921 61620 1955
rect 61568 1912 61620 1921
rect 62396 1955 62448 1964
rect 62396 1921 62405 1955
rect 62405 1921 62439 1955
rect 62439 1921 62448 1955
rect 62396 1912 62448 1921
rect 63224 1955 63276 1964
rect 63224 1921 63233 1955
rect 63233 1921 63267 1955
rect 63267 1921 63276 1955
rect 63224 1912 63276 1921
rect 64052 1955 64104 1964
rect 64052 1921 64061 1955
rect 64061 1921 64095 1955
rect 64095 1921 64104 1955
rect 64052 1912 64104 1921
rect 64880 1887 64932 1896
rect 64880 1853 64889 1887
rect 64889 1853 64923 1887
rect 64923 1853 64932 1887
rect 64880 1844 64932 1853
rect 65708 1955 65760 1964
rect 65708 1921 65717 1955
rect 65717 1921 65751 1955
rect 65751 1921 65760 1955
rect 65708 1912 65760 1921
rect 66628 1955 66680 1964
rect 66628 1921 66637 1955
rect 66637 1921 66671 1955
rect 66671 1921 66680 1955
rect 66628 1912 66680 1921
rect 66720 1955 66772 1964
rect 66720 1921 66729 1955
rect 66729 1921 66763 1955
rect 66763 1921 66772 1955
rect 66720 1912 66772 1921
rect 70860 1955 70912 1964
rect 70860 1921 70869 1955
rect 70869 1921 70903 1955
rect 70903 1921 70912 1955
rect 70860 1912 70912 1921
rect 72332 1955 72384 1964
rect 72332 1921 72341 1955
rect 72341 1921 72375 1955
rect 72375 1921 72384 1955
rect 72332 1912 72384 1921
rect 91008 2048 91060 2100
rect 91100 2091 91152 2100
rect 91100 2057 91109 2091
rect 91109 2057 91143 2091
rect 91143 2057 91152 2091
rect 91100 2048 91152 2057
rect 92756 2091 92808 2100
rect 92756 2057 92765 2091
rect 92765 2057 92799 2091
rect 92799 2057 92808 2091
rect 92756 2048 92808 2057
rect 93676 2048 93728 2100
rect 95424 2091 95476 2100
rect 95424 2057 95433 2091
rect 95433 2057 95467 2091
rect 95467 2057 95476 2091
rect 95424 2048 95476 2057
rect 96252 2091 96304 2100
rect 96252 2057 96261 2091
rect 96261 2057 96295 2091
rect 96295 2057 96304 2091
rect 96252 2048 96304 2057
rect 96344 2048 96396 2100
rect 98644 2048 98696 2100
rect 100668 2048 100720 2100
rect 100760 2048 100812 2100
rect 106556 2048 106608 2100
rect 116400 2048 116452 2100
rect 122012 2091 122064 2100
rect 122012 2057 122021 2091
rect 122021 2057 122055 2091
rect 122055 2057 122064 2091
rect 122012 2048 122064 2057
rect 124496 2091 124548 2100
rect 124496 2057 124505 2091
rect 124505 2057 124539 2091
rect 124539 2057 124548 2091
rect 124496 2048 124548 2057
rect 126244 2091 126296 2100
rect 126244 2057 126253 2091
rect 126253 2057 126287 2091
rect 126287 2057 126296 2091
rect 126244 2048 126296 2057
rect 127900 2091 127952 2100
rect 127900 2057 127909 2091
rect 127909 2057 127943 2091
rect 127943 2057 127952 2091
rect 127900 2048 127952 2057
rect 129648 2091 129700 2100
rect 129648 2057 129657 2091
rect 129657 2057 129691 2091
rect 129691 2057 129700 2091
rect 129648 2048 129700 2057
rect 131672 2091 131724 2100
rect 131672 2057 131681 2091
rect 131681 2057 131715 2091
rect 131715 2057 131724 2091
rect 131672 2048 131724 2057
rect 99380 1980 99432 2032
rect 100208 1980 100260 2032
rect 80152 1955 80204 1964
rect 80152 1921 80161 1955
rect 80161 1921 80195 1955
rect 80195 1921 80204 1955
rect 80152 1912 80204 1921
rect 83740 1912 83792 1964
rect 86408 1955 86460 1964
rect 86408 1921 86417 1955
rect 86417 1921 86451 1955
rect 86451 1921 86460 1955
rect 86408 1912 86460 1921
rect 88064 1955 88116 1964
rect 88064 1921 88073 1955
rect 88073 1921 88107 1955
rect 88107 1921 88116 1955
rect 88064 1912 88116 1921
rect 70584 1887 70636 1896
rect 70584 1853 70593 1887
rect 70593 1853 70627 1887
rect 70627 1853 70636 1887
rect 70584 1844 70636 1853
rect 72056 1887 72108 1896
rect 72056 1853 72065 1887
rect 72065 1853 72099 1887
rect 72099 1853 72108 1887
rect 72056 1844 72108 1853
rect 74264 1887 74316 1896
rect 74264 1853 74273 1887
rect 74273 1853 74307 1887
rect 74307 1853 74316 1887
rect 74264 1844 74316 1853
rect 22192 1776 22244 1828
rect 37832 1776 37884 1828
rect 40316 1819 40368 1828
rect 40316 1785 40325 1819
rect 40325 1785 40359 1819
rect 40359 1785 40368 1819
rect 40316 1776 40368 1785
rect 44548 1776 44600 1828
rect 50528 1776 50580 1828
rect 53932 1776 53984 1828
rect 75736 1887 75788 1896
rect 75736 1853 75745 1887
rect 75745 1853 75779 1887
rect 75779 1853 75788 1887
rect 75736 1844 75788 1853
rect 77208 1887 77260 1896
rect 77208 1853 77217 1887
rect 77217 1853 77251 1887
rect 77251 1853 77260 1887
rect 77208 1844 77260 1853
rect 80060 1844 80112 1896
rect 81348 1844 81400 1896
rect 81440 1887 81492 1896
rect 81440 1853 81449 1887
rect 81449 1853 81483 1887
rect 81483 1853 81492 1887
rect 81440 1844 81492 1853
rect 82636 1844 82688 1896
rect 83832 1887 83884 1896
rect 83832 1853 83841 1887
rect 83841 1853 83875 1887
rect 83875 1853 83884 1887
rect 83832 1844 83884 1853
rect 84016 1887 84068 1896
rect 84016 1853 84025 1887
rect 84025 1853 84059 1887
rect 84059 1853 84068 1887
rect 84016 1844 84068 1853
rect 86040 1844 86092 1896
rect 86132 1887 86184 1896
rect 86132 1853 86141 1887
rect 86141 1853 86175 1887
rect 86175 1853 86184 1887
rect 86132 1844 86184 1853
rect 89168 1912 89220 1964
rect 88524 1844 88576 1896
rect 89076 1887 89128 1896
rect 89076 1853 89085 1887
rect 89085 1853 89119 1887
rect 89119 1853 89128 1887
rect 89076 1844 89128 1853
rect 89904 1912 89956 1964
rect 89996 1955 90048 1964
rect 89996 1921 90005 1955
rect 90005 1921 90039 1955
rect 90039 1921 90048 1955
rect 89996 1912 90048 1921
rect 89536 1844 89588 1896
rect 90732 1955 90784 1964
rect 90732 1921 90741 1955
rect 90741 1921 90775 1955
rect 90775 1921 90784 1955
rect 90732 1912 90784 1921
rect 92020 1844 92072 1896
rect 92296 1912 92348 1964
rect 93308 1955 93360 1964
rect 93308 1921 93317 1955
rect 93317 1921 93351 1955
rect 93351 1921 93360 1955
rect 93308 1912 93360 1921
rect 94136 1955 94188 1964
rect 94136 1921 94145 1955
rect 94145 1921 94179 1955
rect 94179 1921 94188 1955
rect 94136 1912 94188 1921
rect 95148 1955 95200 1964
rect 95148 1921 95157 1955
rect 95157 1921 95191 1955
rect 95191 1921 95200 1955
rect 95148 1912 95200 1921
rect 98552 1955 98604 1964
rect 94964 1844 95016 1896
rect 98552 1921 98561 1955
rect 98561 1921 98595 1955
rect 98595 1921 98604 1955
rect 98552 1912 98604 1921
rect 95240 1776 95292 1828
rect 95976 1776 96028 1828
rect 97540 1887 97592 1896
rect 97540 1853 97549 1887
rect 97549 1853 97583 1887
rect 97583 1853 97592 1887
rect 97540 1844 97592 1853
rect 98368 1887 98420 1896
rect 98368 1853 98377 1887
rect 98377 1853 98411 1887
rect 98411 1853 98420 1887
rect 98368 1844 98420 1853
rect 100116 1912 100168 1964
rect 99840 1844 99892 1896
rect 96804 1776 96856 1828
rect 107108 1955 107160 1964
rect 107108 1921 107117 1955
rect 107117 1921 107151 1955
rect 107151 1921 107160 1955
rect 107108 1912 107160 1921
rect 112260 1955 112312 1964
rect 112260 1921 112269 1955
rect 112269 1921 112303 1955
rect 112303 1921 112312 1955
rect 112260 1912 112312 1921
rect 117320 1912 117372 1964
rect 121184 1980 121236 2032
rect 122840 1912 122892 1964
rect 124128 1955 124180 1964
rect 124128 1921 124137 1955
rect 124137 1921 124171 1955
rect 124171 1921 124180 1955
rect 124128 1912 124180 1921
rect 125048 1955 125100 1964
rect 125048 1921 125057 1955
rect 125057 1921 125091 1955
rect 125091 1921 125100 1955
rect 125048 1912 125100 1921
rect 125968 1955 126020 1964
rect 125968 1921 125977 1955
rect 125977 1921 126011 1955
rect 126011 1921 126020 1955
rect 125968 1912 126020 1921
rect 126704 1955 126756 1964
rect 126704 1921 126713 1955
rect 126713 1921 126747 1955
rect 126747 1921 126756 1955
rect 126704 1912 126756 1921
rect 127624 1955 127676 1964
rect 127624 1921 127633 1955
rect 127633 1921 127667 1955
rect 127667 1921 127676 1955
rect 127624 1912 127676 1921
rect 129188 1980 129240 2032
rect 129556 1980 129608 2032
rect 121644 1887 121696 1896
rect 121644 1853 121653 1887
rect 121653 1853 121687 1887
rect 121687 1853 121696 1887
rect 121644 1844 121696 1853
rect 122472 1887 122524 1896
rect 122472 1853 122481 1887
rect 122481 1853 122515 1887
rect 122515 1853 122524 1887
rect 122472 1844 122524 1853
rect 123300 1887 123352 1896
rect 123300 1853 123309 1887
rect 123309 1853 123343 1887
rect 123343 1853 123352 1887
rect 123300 1844 123352 1853
rect 128452 1844 128504 1896
rect 129556 1844 129608 1896
rect 133604 2023 133656 2032
rect 133604 1989 133613 2023
rect 133613 1989 133647 2023
rect 133647 1989 133656 2023
rect 133604 1980 133656 1989
rect 130568 1955 130620 1964
rect 130568 1921 130577 1955
rect 130577 1921 130611 1955
rect 130611 1921 130620 1955
rect 130568 1912 130620 1921
rect 129740 1844 129792 1896
rect 131120 1912 131172 1964
rect 131856 1912 131908 1964
rect 133052 1912 133104 1964
rect 134984 1980 135036 2032
rect 139952 2023 140004 2032
rect 139952 1989 139961 2023
rect 139961 1989 139995 2023
rect 139995 1989 140004 2023
rect 139952 1980 140004 1989
rect 150808 2048 150860 2100
rect 157892 2048 157944 2100
rect 157984 2048 158036 2100
rect 162124 2048 162176 2100
rect 162308 2091 162360 2100
rect 162308 2057 162317 2091
rect 162317 2057 162351 2091
rect 162351 2057 162360 2091
rect 162308 2048 162360 2057
rect 163964 2091 164016 2100
rect 163964 2057 163973 2091
rect 163973 2057 164007 2091
rect 164007 2057 164016 2091
rect 163964 2048 164016 2057
rect 165620 2091 165672 2100
rect 165620 2057 165629 2091
rect 165629 2057 165663 2091
rect 165663 2057 165672 2091
rect 165620 2048 165672 2057
rect 165896 2048 165948 2100
rect 167460 2091 167512 2100
rect 167460 2057 167469 2091
rect 167469 2057 167503 2091
rect 167503 2057 167512 2091
rect 167460 2048 167512 2057
rect 167552 2048 167604 2100
rect 157156 1980 157208 2032
rect 133144 1844 133196 1896
rect 134064 1844 134116 1896
rect 138112 1955 138164 1964
rect 138112 1921 138121 1955
rect 138121 1921 138155 1955
rect 138155 1921 138164 1955
rect 138112 1912 138164 1921
rect 139032 1955 139084 1964
rect 139032 1921 139041 1955
rect 139041 1921 139075 1955
rect 139075 1921 139084 1955
rect 139032 1912 139084 1921
rect 139216 1912 139268 1964
rect 140412 1912 140464 1964
rect 141424 1955 141476 1964
rect 141424 1921 141433 1955
rect 141433 1921 141467 1955
rect 141467 1921 141476 1955
rect 141424 1912 141476 1921
rect 141700 1955 141752 1964
rect 141700 1921 141709 1955
rect 141709 1921 141743 1955
rect 141743 1921 141752 1955
rect 141700 1912 141752 1921
rect 142988 1955 143040 1964
rect 142988 1921 142997 1955
rect 142997 1921 143031 1955
rect 143031 1921 143040 1955
rect 142988 1912 143040 1921
rect 144920 1955 144972 1964
rect 144920 1921 144929 1955
rect 144929 1921 144963 1955
rect 144963 1921 144972 1955
rect 144920 1912 144972 1921
rect 150072 1955 150124 1964
rect 150072 1921 150081 1955
rect 150081 1921 150115 1955
rect 150115 1921 150124 1955
rect 150072 1912 150124 1921
rect 138296 1887 138348 1896
rect 138296 1853 138305 1887
rect 138305 1853 138339 1887
rect 138339 1853 138348 1887
rect 138296 1844 138348 1853
rect 138388 1844 138440 1896
rect 23664 1708 23716 1760
rect 23756 1708 23808 1760
rect 24860 1708 24912 1760
rect 28908 1708 28960 1760
rect 29736 1708 29788 1760
rect 30564 1708 30616 1760
rect 31760 1751 31812 1760
rect 31760 1717 31769 1751
rect 31769 1717 31803 1751
rect 31803 1717 31812 1751
rect 31760 1708 31812 1717
rect 33140 1708 33192 1760
rect 36820 1751 36872 1760
rect 36820 1717 36829 1751
rect 36829 1717 36863 1751
rect 36863 1717 36872 1751
rect 36820 1708 36872 1717
rect 53472 1751 53524 1760
rect 53472 1717 53481 1751
rect 53481 1717 53515 1751
rect 53515 1717 53524 1751
rect 53472 1708 53524 1717
rect 56048 1708 56100 1760
rect 56876 1708 56928 1760
rect 58440 1708 58492 1760
rect 60648 1708 60700 1760
rect 61384 1708 61436 1760
rect 61844 1751 61896 1760
rect 61844 1717 61853 1751
rect 61853 1717 61887 1751
rect 61887 1717 61896 1751
rect 61844 1708 61896 1717
rect 63592 1751 63644 1760
rect 63592 1717 63601 1751
rect 63601 1717 63635 1751
rect 63635 1717 63644 1751
rect 63592 1708 63644 1717
rect 64328 1708 64380 1760
rect 65984 1708 66036 1760
rect 67548 1751 67600 1760
rect 67548 1717 67557 1751
rect 67557 1717 67591 1751
rect 67591 1717 67600 1751
rect 67548 1708 67600 1717
rect 86040 1751 86092 1760
rect 86040 1717 86049 1751
rect 86049 1717 86083 1751
rect 86083 1717 86092 1751
rect 86040 1708 86092 1717
rect 90456 1708 90508 1760
rect 92020 1708 92072 1760
rect 93308 1708 93360 1760
rect 96620 1708 96672 1760
rect 97172 1708 97224 1760
rect 98552 1708 98604 1760
rect 100116 1708 100168 1760
rect 101312 1751 101364 1760
rect 101312 1717 101321 1751
rect 101321 1717 101355 1751
rect 101355 1717 101364 1751
rect 101312 1708 101364 1717
rect 121184 1751 121236 1760
rect 121184 1717 121193 1751
rect 121193 1717 121227 1751
rect 121227 1717 121236 1751
rect 121184 1708 121236 1717
rect 122932 1708 122984 1760
rect 123760 1708 123812 1760
rect 125416 1751 125468 1760
rect 125416 1717 125425 1751
rect 125425 1717 125459 1751
rect 125459 1717 125468 1751
rect 125416 1708 125468 1717
rect 127072 1751 127124 1760
rect 127072 1717 127081 1751
rect 127081 1717 127115 1751
rect 127115 1717 127124 1751
rect 127072 1708 127124 1717
rect 129096 1708 129148 1760
rect 130660 1708 130712 1760
rect 132592 1751 132644 1760
rect 132592 1717 132601 1751
rect 132601 1717 132635 1751
rect 132635 1717 132644 1751
rect 132592 1708 132644 1717
rect 135260 1708 135312 1760
rect 138848 1844 138900 1896
rect 140688 1887 140740 1896
rect 140688 1853 140697 1887
rect 140697 1853 140731 1887
rect 140731 1853 140740 1887
rect 140688 1844 140740 1853
rect 141516 1887 141568 1896
rect 141516 1853 141550 1887
rect 141550 1853 141568 1887
rect 141516 1844 141568 1853
rect 143172 1844 143224 1896
rect 155040 1844 155092 1896
rect 156696 1912 156748 1964
rect 156788 1955 156840 1964
rect 156788 1921 156797 1955
rect 156797 1921 156831 1955
rect 156831 1921 156840 1955
rect 156788 1912 156840 1921
rect 141148 1819 141200 1828
rect 141148 1785 141157 1819
rect 141157 1785 141191 1819
rect 141191 1785 141200 1819
rect 141148 1776 141200 1785
rect 142804 1819 142856 1828
rect 142804 1785 142813 1819
rect 142813 1785 142847 1819
rect 142847 1785 142856 1819
rect 142804 1776 142856 1785
rect 148140 1776 148192 1828
rect 140780 1708 140832 1760
rect 146484 1708 146536 1760
rect 155776 1776 155828 1828
rect 155960 1708 156012 1760
rect 156512 1844 156564 1896
rect 157984 1955 158036 1964
rect 157984 1921 157993 1955
rect 157993 1921 158027 1955
rect 158027 1921 158036 1955
rect 157984 1912 158036 1921
rect 159272 1955 159324 1964
rect 159272 1921 159281 1955
rect 159281 1921 159315 1955
rect 159315 1921 159324 1955
rect 159272 1912 159324 1921
rect 157064 1887 157116 1896
rect 157064 1853 157073 1887
rect 157073 1853 157107 1887
rect 157107 1853 157116 1887
rect 157064 1844 157116 1853
rect 158168 1844 158220 1896
rect 158536 1844 158588 1896
rect 159640 1912 159692 1964
rect 160008 1844 160060 1896
rect 161204 1955 161256 1964
rect 161204 1921 161213 1955
rect 161213 1921 161247 1955
rect 161247 1921 161256 1955
rect 161204 1912 161256 1921
rect 161572 1912 161624 1964
rect 162216 1912 162268 1964
rect 163688 1955 163740 1964
rect 163688 1921 163697 1955
rect 163697 1921 163731 1955
rect 163731 1921 163740 1955
rect 163688 1912 163740 1921
rect 163780 1955 163832 1964
rect 163780 1921 163789 1955
rect 163789 1921 163823 1955
rect 163823 1921 163832 1955
rect 163780 1912 163832 1921
rect 163136 1844 163188 1896
rect 164332 1912 164384 1964
rect 165252 1955 165304 1964
rect 165252 1921 165261 1955
rect 165261 1921 165295 1955
rect 165295 1921 165304 1955
rect 165252 1912 165304 1921
rect 166264 1955 166316 1964
rect 166264 1921 166273 1955
rect 166273 1921 166307 1955
rect 166307 1921 166316 1955
rect 166264 1912 166316 1921
rect 167092 1955 167144 1964
rect 167092 1921 167101 1955
rect 167101 1921 167135 1955
rect 167135 1921 167144 1955
rect 167092 1912 167144 1921
rect 167184 1844 167236 1896
rect 167920 1955 167972 1964
rect 167920 1921 167929 1955
rect 167929 1921 167963 1955
rect 167963 1921 167972 1955
rect 167920 1912 167972 1921
rect 167828 1844 167880 1896
rect 173256 1955 173308 1964
rect 173256 1921 173265 1955
rect 173265 1921 173299 1955
rect 173299 1921 173308 1955
rect 173256 1912 173308 1921
rect 174728 1955 174780 1964
rect 174728 1921 174737 1955
rect 174737 1921 174771 1955
rect 174771 1921 174780 1955
rect 174728 1912 174780 1921
rect 176844 1955 176896 1964
rect 176844 1921 176853 1955
rect 176853 1921 176887 1955
rect 176887 1921 176896 1955
rect 176844 1912 176896 1921
rect 181904 1955 181956 1964
rect 181904 1921 181913 1955
rect 181913 1921 181947 1955
rect 181947 1921 181956 1955
rect 181904 1912 181956 1921
rect 183560 1955 183612 1964
rect 183560 1921 183569 1955
rect 183569 1921 183603 1955
rect 183603 1921 183612 1955
rect 183560 1912 183612 1921
rect 185032 1955 185084 1964
rect 185032 1921 185041 1955
rect 185041 1921 185075 1955
rect 185075 1921 185084 1955
rect 185032 1912 185084 1921
rect 190368 2048 190420 2100
rect 192392 2091 192444 2100
rect 192392 2057 192401 2091
rect 192401 2057 192435 2091
rect 192435 2057 192444 2091
rect 192392 2048 192444 2057
rect 195704 2091 195756 2100
rect 195704 2057 195713 2091
rect 195713 2057 195747 2091
rect 195747 2057 195756 2091
rect 195704 2048 195756 2057
rect 196256 2048 196308 2100
rect 199200 2091 199252 2100
rect 199200 2057 199209 2091
rect 199209 2057 199243 2091
rect 199243 2057 199252 2091
rect 199200 2048 199252 2057
rect 200856 2091 200908 2100
rect 200856 2057 200865 2091
rect 200865 2057 200899 2091
rect 200899 2057 200908 2091
rect 200856 2048 200908 2057
rect 201316 2048 201368 2100
rect 207020 2048 207072 2100
rect 211160 2048 211212 2100
rect 215392 2048 215444 2100
rect 216956 2048 217008 2100
rect 217140 2091 217192 2100
rect 217140 2057 217149 2091
rect 217149 2057 217183 2091
rect 217183 2057 217192 2091
rect 217140 2048 217192 2057
rect 221832 2048 221884 2100
rect 223028 2048 223080 2100
rect 224224 2048 224276 2100
rect 225328 2091 225380 2100
rect 225328 2057 225337 2091
rect 225337 2057 225371 2091
rect 225371 2057 225380 2091
rect 225328 2048 225380 2057
rect 226156 2091 226208 2100
rect 226156 2057 226165 2091
rect 226165 2057 226199 2091
rect 226199 2057 226208 2091
rect 226156 2048 226208 2057
rect 226984 2091 227036 2100
rect 226984 2057 226993 2091
rect 226993 2057 227027 2091
rect 227027 2057 227036 2091
rect 226984 2048 227036 2057
rect 228088 2048 228140 2100
rect 229192 2048 229244 2100
rect 236000 2048 236052 2100
rect 236092 2091 236144 2100
rect 236092 2057 236101 2091
rect 236101 2057 236135 2091
rect 236135 2057 236144 2091
rect 236092 2048 236144 2057
rect 189724 1955 189776 1964
rect 189724 1921 189733 1955
rect 189733 1921 189767 1955
rect 189767 1921 189776 1955
rect 189724 1912 189776 1921
rect 190828 1955 190880 1964
rect 190828 1921 190837 1955
rect 190837 1921 190871 1955
rect 190871 1921 190880 1955
rect 190828 1912 190880 1921
rect 190920 1955 190972 1964
rect 190920 1921 190929 1955
rect 190929 1921 190963 1955
rect 190963 1921 190972 1955
rect 190920 1912 190972 1921
rect 192300 1980 192352 2032
rect 193312 1980 193364 2032
rect 172980 1887 173032 1896
rect 172980 1853 172989 1887
rect 172989 1853 173023 1887
rect 173023 1853 173032 1887
rect 172980 1844 173032 1853
rect 174452 1887 174504 1896
rect 174452 1853 174461 1887
rect 174461 1853 174495 1887
rect 174495 1853 174504 1887
rect 174452 1844 174504 1853
rect 176568 1887 176620 1896
rect 176568 1853 176577 1887
rect 176577 1853 176611 1887
rect 176611 1853 176620 1887
rect 176568 1844 176620 1853
rect 177856 1887 177908 1896
rect 177856 1853 177865 1887
rect 177865 1853 177899 1887
rect 177899 1853 177908 1887
rect 177856 1844 177908 1853
rect 156880 1776 156932 1828
rect 179144 1887 179196 1896
rect 179144 1853 179153 1887
rect 179153 1853 179187 1887
rect 179187 1853 179196 1887
rect 179144 1844 179196 1853
rect 183284 1887 183336 1896
rect 183284 1853 183293 1887
rect 183293 1853 183327 1887
rect 183327 1853 183336 1887
rect 183284 1844 183336 1853
rect 184756 1887 184808 1896
rect 184756 1853 184765 1887
rect 184765 1853 184799 1887
rect 184799 1853 184808 1887
rect 184756 1844 184808 1853
rect 186320 1844 186372 1896
rect 188160 1887 188212 1896
rect 188160 1853 188169 1887
rect 188169 1853 188203 1887
rect 188203 1853 188212 1887
rect 188160 1844 188212 1853
rect 179512 1776 179564 1828
rect 189448 1887 189500 1896
rect 189448 1853 189457 1887
rect 189457 1853 189491 1887
rect 189491 1853 189500 1887
rect 189448 1844 189500 1853
rect 193220 1912 193272 1964
rect 194600 1955 194652 1964
rect 194600 1921 194609 1955
rect 194609 1921 194643 1955
rect 194643 1921 194652 1955
rect 194600 1912 194652 1921
rect 195428 1955 195480 1964
rect 195428 1921 195437 1955
rect 195437 1921 195471 1955
rect 195471 1921 195480 1955
rect 195428 1912 195480 1921
rect 196164 1955 196216 1964
rect 196164 1921 196173 1955
rect 196173 1921 196207 1955
rect 196207 1921 196216 1955
rect 196164 1912 196216 1921
rect 196440 1912 196492 1964
rect 197268 1912 197320 1964
rect 198004 1955 198056 1964
rect 198004 1921 198013 1955
rect 198013 1921 198047 1955
rect 198047 1921 198056 1955
rect 198004 1912 198056 1921
rect 198832 1955 198884 1964
rect 198832 1921 198841 1955
rect 198841 1921 198875 1955
rect 198875 1921 198884 1955
rect 198832 1912 198884 1921
rect 199660 1955 199712 1964
rect 199660 1921 199669 1955
rect 199669 1921 199703 1955
rect 199703 1921 199712 1955
rect 199660 1912 199712 1921
rect 200488 1955 200540 1964
rect 200488 1921 200497 1955
rect 200497 1921 200531 1955
rect 200531 1921 200540 1955
rect 200488 1912 200540 1921
rect 201132 1912 201184 1964
rect 202236 1912 202288 1964
rect 216680 2023 216732 2032
rect 216680 1989 216689 2023
rect 216689 1989 216723 2023
rect 216723 1989 216732 2023
rect 216680 1980 216732 1989
rect 211712 1955 211764 1964
rect 211712 1921 211721 1955
rect 211721 1921 211755 1955
rect 211755 1921 211764 1955
rect 211712 1912 211764 1921
rect 216404 1955 216456 1964
rect 216404 1921 216413 1955
rect 216413 1921 216447 1955
rect 216447 1921 216456 1955
rect 216404 1912 216456 1921
rect 219440 1912 219492 1964
rect 222568 1980 222620 2032
rect 220084 1955 220136 1964
rect 220084 1921 220093 1955
rect 220093 1921 220127 1955
rect 220127 1921 220136 1955
rect 220084 1912 220136 1921
rect 220728 1955 220780 1964
rect 220728 1921 220737 1955
rect 220737 1921 220771 1955
rect 220771 1921 220780 1955
rect 220728 1912 220780 1921
rect 220820 1912 220872 1964
rect 222476 1912 222528 1964
rect 223212 1955 223264 1964
rect 223212 1921 223221 1955
rect 223221 1921 223255 1955
rect 223255 1921 223264 1955
rect 223212 1912 223264 1921
rect 223948 1980 224000 2032
rect 225512 1980 225564 2032
rect 224408 1912 224460 1964
rect 224776 1912 224828 1964
rect 218060 1844 218112 1896
rect 216680 1776 216732 1828
rect 221004 1887 221056 1896
rect 221004 1853 221013 1887
rect 221013 1853 221047 1887
rect 221047 1853 221056 1887
rect 221004 1844 221056 1853
rect 222108 1844 222160 1896
rect 223856 1776 223908 1828
rect 224868 1844 224920 1896
rect 225880 1955 225932 1964
rect 225880 1921 225889 1955
rect 225889 1921 225923 1955
rect 225923 1921 225932 1955
rect 225880 1912 225932 1921
rect 226708 1955 226760 1964
rect 226708 1921 226717 1955
rect 226717 1921 226751 1955
rect 226751 1921 226760 1955
rect 226708 1912 226760 1921
rect 226616 1844 226668 1896
rect 227720 1912 227772 1964
rect 228916 1955 228968 1964
rect 228916 1921 228925 1955
rect 228925 1921 228959 1955
rect 228959 1921 228968 1955
rect 228916 1912 228968 1921
rect 228364 1844 228416 1896
rect 229468 1912 229520 1964
rect 229744 1955 229796 1964
rect 229744 1921 229753 1955
rect 229753 1921 229787 1955
rect 229787 1921 229796 1955
rect 229744 1912 229796 1921
rect 229928 1955 229980 1964
rect 229928 1921 229957 1955
rect 229957 1921 229980 1955
rect 231768 2023 231820 2032
rect 231768 1989 231777 2023
rect 231777 1989 231811 2023
rect 231811 1989 231820 2023
rect 231768 1980 231820 1989
rect 231860 1980 231912 2032
rect 229928 1912 229980 1921
rect 230112 1912 230164 1964
rect 230756 1955 230808 1964
rect 230756 1921 230765 1955
rect 230765 1921 230799 1955
rect 230799 1921 230808 1955
rect 230756 1912 230808 1921
rect 231492 1955 231544 1964
rect 231492 1921 231501 1955
rect 231501 1921 231535 1955
rect 231535 1921 231544 1955
rect 231492 1912 231544 1921
rect 231584 1955 231636 1964
rect 231584 1921 231593 1955
rect 231593 1921 231627 1955
rect 231627 1921 231636 1955
rect 231584 1912 231636 1921
rect 232136 1912 232188 1964
rect 232320 1912 232372 1964
rect 233240 1912 233292 1964
rect 233700 1980 233752 2032
rect 233884 1980 233936 2032
rect 251456 2091 251508 2100
rect 251456 2057 251465 2091
rect 251465 2057 251499 2091
rect 251499 2057 251508 2091
rect 251456 2048 251508 2057
rect 257620 2048 257672 2100
rect 258908 2048 258960 2100
rect 259000 2048 259052 2100
rect 233424 1955 233476 1964
rect 233424 1921 233433 1955
rect 233433 1921 233467 1955
rect 233467 1921 233476 1955
rect 233424 1912 233476 1921
rect 229836 1844 229888 1896
rect 234068 1887 234120 1896
rect 234068 1853 234077 1887
rect 234077 1853 234111 1887
rect 234111 1853 234120 1887
rect 234068 1844 234120 1853
rect 234896 1955 234948 1964
rect 234896 1921 234905 1955
rect 234905 1921 234939 1955
rect 234939 1921 234948 1955
rect 234896 1912 234948 1921
rect 236000 1912 236052 1964
rect 237932 1912 237984 1964
rect 240048 1912 240100 1964
rect 243176 1980 243228 2032
rect 257804 1980 257856 2032
rect 251180 1912 251232 1964
rect 252560 1955 252612 1964
rect 252560 1921 252569 1955
rect 252569 1921 252603 1955
rect 252603 1921 252612 1955
rect 252560 1912 252612 1921
rect 255412 1955 255464 1964
rect 255412 1921 255421 1955
rect 255421 1921 255455 1955
rect 255455 1921 255464 1955
rect 255412 1912 255464 1921
rect 256884 1912 256936 1964
rect 257896 1955 257948 1964
rect 257896 1921 257905 1955
rect 257905 1921 257939 1955
rect 257939 1921 257948 1955
rect 257896 1912 257948 1921
rect 259092 1980 259144 2032
rect 258908 1912 258960 1964
rect 259828 1912 259880 1964
rect 261576 2048 261628 2100
rect 269672 2091 269724 2100
rect 269672 2057 269681 2091
rect 269681 2057 269715 2091
rect 269715 2057 269724 2091
rect 269672 2048 269724 2057
rect 269764 2048 269816 2100
rect 260104 1980 260156 2032
rect 264152 1980 264204 2032
rect 267556 1980 267608 2032
rect 235724 1887 235776 1896
rect 235724 1853 235733 1887
rect 235733 1853 235767 1887
rect 235767 1853 235776 1887
rect 235724 1844 235776 1853
rect 235816 1844 235868 1896
rect 241244 1887 241296 1896
rect 241244 1853 241253 1887
rect 241253 1853 241287 1887
rect 241287 1853 241296 1887
rect 241244 1844 241296 1853
rect 242900 1844 242952 1896
rect 243820 1887 243872 1896
rect 243820 1853 243829 1887
rect 243829 1853 243863 1887
rect 243863 1853 243872 1887
rect 243820 1844 243872 1853
rect 244280 1844 244332 1896
rect 246120 1887 246172 1896
rect 246120 1853 246129 1887
rect 246129 1853 246163 1887
rect 246163 1853 246172 1887
rect 246120 1844 246172 1853
rect 160192 1708 160244 1760
rect 161480 1751 161532 1760
rect 161480 1717 161489 1751
rect 161489 1717 161523 1751
rect 161523 1717 161532 1751
rect 161480 1708 161532 1717
rect 163136 1751 163188 1760
rect 163136 1717 163145 1751
rect 163145 1717 163179 1751
rect 163179 1717 163188 1751
rect 163136 1708 163188 1717
rect 164516 1708 164568 1760
rect 168380 1708 168432 1760
rect 181996 1751 182048 1760
rect 181996 1717 182005 1751
rect 182005 1717 182039 1751
rect 182039 1717 182048 1751
rect 181996 1708 182048 1717
rect 193220 1751 193272 1760
rect 193220 1717 193229 1751
rect 193229 1717 193263 1751
rect 193263 1717 193272 1751
rect 193220 1708 193272 1717
rect 193312 1708 193364 1760
rect 194600 1708 194652 1760
rect 196532 1751 196584 1760
rect 196532 1717 196541 1751
rect 196541 1717 196575 1751
rect 196575 1717 196584 1751
rect 196532 1708 196584 1717
rect 197912 1708 197964 1760
rect 199752 1708 199804 1760
rect 201684 1751 201736 1760
rect 201684 1717 201693 1751
rect 201693 1717 201727 1751
rect 201727 1717 201736 1751
rect 201684 1708 201736 1717
rect 202880 1708 202932 1760
rect 216128 1708 216180 1760
rect 224316 1708 224368 1760
rect 225512 1708 225564 1760
rect 229192 1708 229244 1760
rect 229284 1751 229336 1760
rect 229284 1717 229293 1751
rect 229293 1717 229327 1751
rect 229327 1717 229336 1751
rect 229284 1708 229336 1717
rect 229652 1708 229704 1760
rect 230664 1708 230716 1760
rect 231584 1708 231636 1760
rect 232320 1708 232372 1760
rect 233240 1708 233292 1760
rect 239496 1776 239548 1828
rect 242532 1776 242584 1828
rect 248420 1844 248472 1896
rect 248972 1887 249024 1896
rect 248972 1853 248981 1887
rect 248981 1853 249015 1887
rect 249015 1853 249024 1887
rect 248972 1844 249024 1853
rect 249800 1844 249852 1896
rect 252284 1887 252336 1896
rect 252284 1853 252293 1887
rect 252293 1853 252327 1887
rect 252327 1853 252336 1887
rect 252284 1844 252336 1853
rect 253848 1887 253900 1896
rect 253848 1853 253857 1887
rect 253857 1853 253891 1887
rect 253891 1853 253900 1887
rect 253848 1844 253900 1853
rect 254032 1844 254084 1896
rect 255136 1887 255188 1896
rect 255136 1853 255145 1887
rect 255145 1853 255179 1887
rect 255179 1853 255188 1887
rect 255136 1844 255188 1853
rect 256424 1887 256476 1896
rect 256424 1853 256433 1887
rect 256433 1853 256467 1887
rect 256467 1853 256476 1887
rect 256424 1844 256476 1853
rect 260288 1912 260340 1964
rect 261484 1955 261536 1964
rect 261484 1921 261493 1955
rect 261493 1921 261527 1955
rect 261527 1921 261536 1955
rect 261484 1912 261536 1921
rect 262312 1955 262364 1964
rect 262312 1921 262321 1955
rect 262321 1921 262355 1955
rect 262355 1921 262364 1955
rect 262312 1912 262364 1921
rect 262588 1912 262640 1964
rect 264244 1912 264296 1964
rect 269212 1912 269264 1964
rect 269764 1912 269816 1964
rect 270500 2091 270552 2100
rect 270500 2057 270509 2091
rect 270509 2057 270543 2091
rect 270543 2057 270552 2091
rect 270500 2048 270552 2057
rect 271144 1980 271196 2032
rect 272156 1980 272208 2032
rect 263416 1844 263468 1896
rect 265072 1844 265124 1896
rect 265808 1887 265860 1896
rect 265808 1853 265817 1887
rect 265817 1853 265851 1887
rect 265851 1853 265860 1887
rect 265808 1844 265860 1853
rect 266636 1887 266688 1896
rect 266636 1853 266645 1887
rect 266645 1853 266679 1887
rect 266679 1853 266688 1887
rect 266636 1844 266688 1853
rect 266728 1844 266780 1896
rect 268292 1887 268344 1896
rect 268292 1853 268301 1887
rect 268301 1853 268335 1887
rect 268335 1853 268344 1887
rect 268292 1844 268344 1853
rect 270868 1844 270920 1896
rect 259276 1776 259328 1828
rect 269028 1776 269080 1828
rect 233884 1708 233936 1760
rect 233976 1708 234028 1760
rect 234712 1708 234764 1760
rect 237288 1708 237340 1760
rect 257896 1708 257948 1760
rect 260104 1708 260156 1760
rect 260288 1708 260340 1760
rect 261576 1708 261628 1760
rect 262312 1708 262364 1760
rect 263048 1708 263100 1760
rect 264152 1708 264204 1760
rect 265164 1708 265216 1760
rect 265900 1708 265952 1760
rect 266728 1708 266780 1760
rect 267832 1751 267884 1760
rect 267832 1717 267841 1751
rect 267841 1717 267875 1751
rect 267875 1717 267884 1751
rect 267832 1708 267884 1717
rect 268200 1708 268252 1760
rect 34748 1606 34800 1658
rect 34812 1606 34864 1658
rect 34876 1606 34928 1658
rect 34940 1606 34992 1658
rect 35004 1606 35056 1658
rect 102345 1606 102397 1658
rect 102409 1606 102461 1658
rect 102473 1606 102525 1658
rect 102537 1606 102589 1658
rect 102601 1606 102653 1658
rect 169942 1606 169994 1658
rect 170006 1606 170058 1658
rect 170070 1606 170122 1658
rect 170134 1606 170186 1658
rect 170198 1606 170250 1658
rect 237539 1606 237591 1658
rect 237603 1606 237655 1658
rect 237667 1606 237719 1658
rect 237731 1606 237783 1658
rect 237795 1606 237847 1658
rect 22100 1504 22152 1556
rect 28540 1504 28592 1556
rect 35532 1504 35584 1556
rect 35624 1504 35676 1556
rect 58900 1504 58952 1556
rect 60004 1547 60056 1556
rect 60004 1513 60013 1547
rect 60013 1513 60047 1547
rect 60047 1513 60056 1547
rect 60004 1504 60056 1513
rect 94412 1504 94464 1556
rect 95240 1504 95292 1556
rect 99196 1504 99248 1556
rect 99380 1504 99432 1556
rect 107384 1504 107436 1556
rect 113272 1504 113324 1556
rect 121644 1504 121696 1556
rect 156512 1504 156564 1556
rect 156696 1504 156748 1556
rect 157340 1504 157392 1556
rect 175832 1504 175884 1556
rect 23664 1436 23716 1488
rect 30932 1436 30984 1488
rect 31024 1436 31076 1488
rect 848 1368 900 1420
rect 24032 1368 24084 1420
rect 24952 1411 25004 1420
rect 2872 1343 2924 1352
rect 2872 1309 2881 1343
rect 2881 1309 2915 1343
rect 2915 1309 2924 1343
rect 2872 1300 2924 1309
rect 5172 1343 5224 1352
rect 5172 1309 5181 1343
rect 5181 1309 5215 1343
rect 5215 1309 5224 1343
rect 5172 1300 5224 1309
rect 5448 1343 5500 1352
rect 5448 1309 5457 1343
rect 5457 1309 5491 1343
rect 5491 1309 5500 1343
rect 5448 1300 5500 1309
rect 6552 1343 6604 1352
rect 6552 1309 6561 1343
rect 6561 1309 6595 1343
rect 6595 1309 6604 1343
rect 6552 1300 6604 1309
rect 9404 1300 9456 1352
rect 9588 1300 9640 1352
rect 11152 1343 11204 1352
rect 11152 1309 11161 1343
rect 11161 1309 11195 1343
rect 11195 1309 11204 1343
rect 11152 1300 11204 1309
rect 12164 1343 12216 1352
rect 12164 1309 12173 1343
rect 12173 1309 12207 1343
rect 12207 1309 12216 1343
rect 12164 1300 12216 1309
rect 14832 1343 14884 1352
rect 14832 1309 14841 1343
rect 14841 1309 14875 1343
rect 14875 1309 14884 1343
rect 14832 1300 14884 1309
rect 15108 1343 15160 1352
rect 15108 1309 15117 1343
rect 15117 1309 15151 1343
rect 15151 1309 15160 1343
rect 15108 1300 15160 1309
rect 23756 1343 23808 1352
rect 23756 1309 23765 1343
rect 23765 1309 23799 1343
rect 23799 1309 23808 1343
rect 23756 1300 23808 1309
rect 24952 1377 24961 1411
rect 24961 1377 24995 1411
rect 24995 1377 25004 1411
rect 24952 1368 25004 1377
rect 25044 1368 25096 1420
rect 25872 1368 25924 1420
rect 27804 1368 27856 1420
rect 34428 1368 34480 1420
rect 36728 1479 36780 1488
rect 36728 1445 36737 1479
rect 36737 1445 36771 1479
rect 36771 1445 36780 1479
rect 36728 1436 36780 1445
rect 38660 1479 38712 1488
rect 38660 1445 38669 1479
rect 38669 1445 38703 1479
rect 38703 1445 38712 1479
rect 38660 1436 38712 1445
rect 43352 1436 43404 1488
rect 53472 1368 53524 1420
rect 54116 1436 54168 1488
rect 86040 1436 86092 1488
rect 99012 1436 99064 1488
rect 101588 1436 101640 1488
rect 133236 1436 133288 1488
rect 133328 1479 133380 1488
rect 133328 1445 133337 1479
rect 133337 1445 133371 1479
rect 133371 1445 133380 1479
rect 133328 1436 133380 1445
rect 134340 1479 134392 1488
rect 134340 1445 134349 1479
rect 134349 1445 134383 1479
rect 134383 1445 134392 1479
rect 134340 1436 134392 1445
rect 138020 1436 138072 1488
rect 138296 1436 138348 1488
rect 140688 1436 140740 1488
rect 144184 1436 144236 1488
rect 176936 1436 176988 1488
rect 180616 1547 180668 1556
rect 180616 1513 180625 1547
rect 180625 1513 180659 1547
rect 180659 1513 180668 1547
rect 180616 1504 180668 1513
rect 216588 1504 216640 1556
rect 220636 1504 220688 1556
rect 226248 1504 226300 1556
rect 226432 1504 226484 1556
rect 191380 1479 191432 1488
rect 191380 1445 191389 1479
rect 191389 1445 191423 1479
rect 191423 1445 191432 1479
rect 191380 1436 191432 1445
rect 69112 1411 69164 1420
rect 69112 1377 69121 1411
rect 69121 1377 69155 1411
rect 69155 1377 69164 1411
rect 69112 1368 69164 1377
rect 87788 1368 87840 1420
rect 2964 1232 3016 1284
rect 4068 1275 4120 1284
rect 4068 1241 4077 1275
rect 4077 1241 4111 1275
rect 4111 1241 4120 1275
rect 4068 1232 4120 1241
rect 8208 1232 8260 1284
rect 9680 1275 9732 1284
rect 9680 1241 9689 1275
rect 9689 1241 9723 1275
rect 9723 1241 9732 1275
rect 9680 1232 9732 1241
rect 10232 1275 10284 1284
rect 10232 1241 10241 1275
rect 10241 1241 10275 1275
rect 10275 1241 10284 1275
rect 10232 1232 10284 1241
rect 10416 1275 10468 1284
rect 10416 1241 10425 1275
rect 10425 1241 10459 1275
rect 10459 1241 10468 1275
rect 10416 1232 10468 1241
rect 10968 1275 11020 1284
rect 10968 1241 10977 1275
rect 10977 1241 11011 1275
rect 11011 1241 11020 1275
rect 10968 1232 11020 1241
rect 11980 1275 12032 1284
rect 11980 1241 11989 1275
rect 11989 1241 12023 1275
rect 12023 1241 12032 1275
rect 11980 1232 12032 1241
rect 12716 1275 12768 1284
rect 12716 1241 12725 1275
rect 12725 1241 12759 1275
rect 12759 1241 12768 1275
rect 12716 1232 12768 1241
rect 13452 1275 13504 1284
rect 13452 1241 13461 1275
rect 13461 1241 13495 1275
rect 13495 1241 13504 1275
rect 13452 1232 13504 1241
rect 17132 1275 17184 1284
rect 17132 1241 17141 1275
rect 17141 1241 17175 1275
rect 17175 1241 17184 1275
rect 17132 1232 17184 1241
rect 17868 1275 17920 1284
rect 17868 1241 17877 1275
rect 17877 1241 17911 1275
rect 17911 1241 17920 1275
rect 17868 1232 17920 1241
rect 18604 1275 18656 1284
rect 18604 1241 18613 1275
rect 18613 1241 18647 1275
rect 18647 1241 18656 1275
rect 18604 1232 18656 1241
rect 27528 1343 27580 1352
rect 27528 1309 27537 1343
rect 27537 1309 27571 1343
rect 27571 1309 27580 1343
rect 27528 1300 27580 1309
rect 28908 1343 28960 1352
rect 28908 1309 28917 1343
rect 28917 1309 28951 1343
rect 28951 1309 28960 1343
rect 28908 1300 28960 1309
rect 29736 1343 29788 1352
rect 29736 1309 29745 1343
rect 29745 1309 29779 1343
rect 29779 1309 29788 1343
rect 29736 1300 29788 1309
rect 30564 1343 30616 1352
rect 30564 1309 30573 1343
rect 30573 1309 30607 1343
rect 30607 1309 30616 1343
rect 30564 1300 30616 1309
rect 31760 1300 31812 1352
rect 32312 1343 32364 1352
rect 32312 1309 32321 1343
rect 32321 1309 32355 1343
rect 32355 1309 32364 1343
rect 32312 1300 32364 1309
rect 35624 1343 35676 1352
rect 35624 1309 35633 1343
rect 35633 1309 35667 1343
rect 35667 1309 35676 1343
rect 35624 1300 35676 1309
rect 36268 1343 36320 1352
rect 36268 1309 36277 1343
rect 36277 1309 36311 1343
rect 36311 1309 36320 1343
rect 36268 1300 36320 1309
rect 36912 1343 36964 1352
rect 36912 1309 36921 1343
rect 36921 1309 36955 1343
rect 36955 1309 36964 1343
rect 36912 1300 36964 1309
rect 38568 1300 38620 1352
rect 38844 1343 38896 1352
rect 38844 1309 38853 1343
rect 38853 1309 38887 1343
rect 38887 1309 38896 1343
rect 38844 1300 38896 1309
rect 39948 1300 40000 1352
rect 40776 1343 40828 1352
rect 40776 1309 40785 1343
rect 40785 1309 40819 1343
rect 40819 1309 40828 1343
rect 40776 1300 40828 1309
rect 41420 1343 41472 1352
rect 41420 1309 41429 1343
rect 41429 1309 41463 1343
rect 41463 1309 41472 1343
rect 41420 1300 41472 1309
rect 42064 1343 42116 1352
rect 42064 1309 42073 1343
rect 42073 1309 42107 1343
rect 42107 1309 42116 1343
rect 42064 1300 42116 1309
rect 43260 1343 43312 1352
rect 43260 1309 43269 1343
rect 43269 1309 43303 1343
rect 43303 1309 43312 1343
rect 43260 1300 43312 1309
rect 43996 1343 44048 1352
rect 43996 1309 44005 1343
rect 44005 1309 44039 1343
rect 44039 1309 44048 1343
rect 43996 1300 44048 1309
rect 44640 1343 44692 1352
rect 44640 1309 44649 1343
rect 44649 1309 44683 1343
rect 44683 1309 44692 1343
rect 44640 1300 44692 1309
rect 45928 1343 45980 1352
rect 45928 1309 45937 1343
rect 45937 1309 45971 1343
rect 45971 1309 45980 1343
rect 45928 1300 45980 1309
rect 46572 1343 46624 1352
rect 46572 1309 46581 1343
rect 46581 1309 46615 1343
rect 46615 1309 46624 1343
rect 46572 1300 46624 1309
rect 47216 1343 47268 1352
rect 47216 1309 47225 1343
rect 47225 1309 47259 1343
rect 47259 1309 47268 1343
rect 47216 1300 47268 1309
rect 48320 1300 48372 1352
rect 49148 1343 49200 1352
rect 49148 1309 49157 1343
rect 49157 1309 49191 1343
rect 49191 1309 49200 1343
rect 49148 1300 49200 1309
rect 49792 1343 49844 1352
rect 49792 1309 49801 1343
rect 49801 1309 49835 1343
rect 49835 1309 49844 1343
rect 49792 1300 49844 1309
rect 51080 1343 51132 1352
rect 51080 1309 51089 1343
rect 51089 1309 51123 1343
rect 51123 1309 51132 1343
rect 51080 1300 51132 1309
rect 51724 1343 51776 1352
rect 51724 1309 51733 1343
rect 51733 1309 51767 1343
rect 51767 1309 51776 1343
rect 51724 1300 51776 1309
rect 52368 1343 52420 1352
rect 52368 1309 52377 1343
rect 52377 1309 52411 1343
rect 52411 1309 52420 1343
rect 52368 1300 52420 1309
rect 53840 1300 53892 1352
rect 54024 1300 54076 1352
rect 56048 1343 56100 1352
rect 56048 1309 56057 1343
rect 56057 1309 56091 1343
rect 56091 1309 56100 1343
rect 56048 1300 56100 1309
rect 56876 1343 56928 1352
rect 56876 1309 56885 1343
rect 56885 1309 56919 1343
rect 56919 1309 56928 1343
rect 56876 1300 56928 1309
rect 58440 1343 58492 1352
rect 58440 1309 58449 1343
rect 58449 1309 58483 1343
rect 58483 1309 58492 1343
rect 58440 1300 58492 1309
rect 59728 1343 59780 1352
rect 59728 1309 59737 1343
rect 59737 1309 59771 1343
rect 59771 1309 59780 1343
rect 59728 1300 59780 1309
rect 59912 1300 59964 1352
rect 60648 1343 60700 1352
rect 60648 1309 60657 1343
rect 60657 1309 60691 1343
rect 60691 1309 60700 1343
rect 60648 1300 60700 1309
rect 61384 1343 61436 1352
rect 61384 1309 61393 1343
rect 61393 1309 61427 1343
rect 61427 1309 61436 1343
rect 61384 1300 61436 1309
rect 61844 1300 61896 1352
rect 63592 1343 63644 1352
rect 63592 1309 63601 1343
rect 63601 1309 63635 1343
rect 63635 1309 63644 1343
rect 63592 1300 63644 1309
rect 64328 1343 64380 1352
rect 64328 1309 64337 1343
rect 64337 1309 64371 1343
rect 64371 1309 64380 1343
rect 64328 1300 64380 1309
rect 65984 1343 66036 1352
rect 65984 1309 65993 1343
rect 65993 1309 66027 1343
rect 66027 1309 66036 1343
rect 65984 1300 66036 1309
rect 69572 1343 69624 1352
rect 69572 1309 69581 1343
rect 69581 1309 69615 1343
rect 69615 1309 69624 1343
rect 69572 1300 69624 1309
rect 69848 1343 69900 1352
rect 69848 1309 69857 1343
rect 69857 1309 69891 1343
rect 69891 1309 69900 1343
rect 69848 1300 69900 1309
rect 72148 1343 72200 1352
rect 72148 1309 72157 1343
rect 72157 1309 72191 1343
rect 72191 1309 72200 1343
rect 72148 1300 72200 1309
rect 72424 1343 72476 1352
rect 72424 1309 72433 1343
rect 72433 1309 72467 1343
rect 72467 1309 72476 1343
rect 72424 1300 72476 1309
rect 74724 1343 74776 1352
rect 74724 1309 74733 1343
rect 74733 1309 74767 1343
rect 74767 1309 74776 1343
rect 74724 1300 74776 1309
rect 75000 1343 75052 1352
rect 75000 1309 75009 1343
rect 75009 1309 75043 1343
rect 75043 1309 75052 1343
rect 75000 1300 75052 1309
rect 42984 1232 43036 1284
rect 4160 1207 4212 1216
rect 4160 1173 4169 1207
rect 4169 1173 4203 1207
rect 4203 1173 4212 1207
rect 4160 1164 4212 1173
rect 8392 1207 8444 1216
rect 8392 1173 8401 1207
rect 8401 1173 8435 1207
rect 8435 1173 8444 1207
rect 8392 1164 8444 1173
rect 12808 1207 12860 1216
rect 12808 1173 12817 1207
rect 12817 1173 12851 1207
rect 12851 1173 12860 1207
rect 12808 1164 12860 1173
rect 13544 1207 13596 1216
rect 13544 1173 13553 1207
rect 13553 1173 13587 1207
rect 13587 1173 13596 1207
rect 13544 1164 13596 1173
rect 17224 1207 17276 1216
rect 17224 1173 17233 1207
rect 17233 1173 17267 1207
rect 17267 1173 17276 1207
rect 17224 1164 17276 1173
rect 17960 1207 18012 1216
rect 17960 1173 17969 1207
rect 17969 1173 18003 1207
rect 18003 1173 18012 1207
rect 17960 1164 18012 1173
rect 18696 1207 18748 1216
rect 18696 1173 18705 1207
rect 18705 1173 18739 1207
rect 18739 1173 18748 1207
rect 18696 1164 18748 1173
rect 23940 1207 23992 1216
rect 23940 1173 23949 1207
rect 23949 1173 23983 1207
rect 23983 1173 23992 1207
rect 23940 1164 23992 1173
rect 29000 1164 29052 1216
rect 29920 1207 29972 1216
rect 29920 1173 29929 1207
rect 29929 1173 29963 1207
rect 29963 1173 29972 1207
rect 29920 1164 29972 1173
rect 30380 1164 30432 1216
rect 31576 1207 31628 1216
rect 31576 1173 31585 1207
rect 31585 1173 31619 1207
rect 31619 1173 31628 1207
rect 31576 1164 31628 1173
rect 32496 1207 32548 1216
rect 32496 1173 32505 1207
rect 32505 1173 32539 1207
rect 32539 1173 32548 1207
rect 32496 1164 32548 1173
rect 36084 1207 36136 1216
rect 36084 1173 36093 1207
rect 36093 1173 36127 1207
rect 36127 1173 36136 1207
rect 36084 1164 36136 1173
rect 38016 1207 38068 1216
rect 38016 1173 38025 1207
rect 38025 1173 38059 1207
rect 38059 1173 38068 1207
rect 38016 1164 38068 1173
rect 39856 1164 39908 1216
rect 40592 1207 40644 1216
rect 40592 1173 40601 1207
rect 40601 1173 40635 1207
rect 40635 1173 40644 1207
rect 40592 1164 40644 1173
rect 41236 1207 41288 1216
rect 41236 1173 41245 1207
rect 41245 1173 41279 1207
rect 41279 1173 41288 1207
rect 41236 1164 41288 1173
rect 41512 1164 41564 1216
rect 43076 1207 43128 1216
rect 43076 1173 43085 1207
rect 43085 1173 43119 1207
rect 43119 1173 43128 1207
rect 43076 1164 43128 1173
rect 46664 1232 46716 1284
rect 45008 1164 45060 1216
rect 45836 1164 45888 1216
rect 46848 1164 46900 1216
rect 52920 1232 52972 1284
rect 77576 1343 77628 1352
rect 77576 1309 77585 1343
rect 77585 1309 77619 1343
rect 77619 1309 77628 1343
rect 77576 1300 77628 1309
rect 79968 1300 80020 1352
rect 78588 1232 78640 1284
rect 48872 1164 48924 1216
rect 49608 1207 49660 1216
rect 49608 1173 49617 1207
rect 49617 1173 49651 1207
rect 49651 1173 49660 1207
rect 49608 1164 49660 1173
rect 50712 1164 50764 1216
rect 51540 1207 51592 1216
rect 51540 1173 51549 1207
rect 51549 1173 51583 1207
rect 51583 1173 51592 1207
rect 51540 1164 51592 1173
rect 52000 1164 52052 1216
rect 53380 1207 53432 1216
rect 53380 1173 53389 1207
rect 53389 1173 53423 1207
rect 53423 1173 53432 1207
rect 53380 1164 53432 1173
rect 56232 1207 56284 1216
rect 56232 1173 56241 1207
rect 56241 1173 56275 1207
rect 56275 1173 56284 1207
rect 56232 1164 56284 1173
rect 57060 1207 57112 1216
rect 57060 1173 57069 1207
rect 57069 1173 57103 1207
rect 57103 1173 57112 1207
rect 57060 1164 57112 1173
rect 58624 1207 58676 1216
rect 58624 1173 58633 1207
rect 58633 1173 58667 1207
rect 58667 1173 58676 1207
rect 58624 1164 58676 1173
rect 60832 1207 60884 1216
rect 60832 1173 60841 1207
rect 60841 1173 60875 1207
rect 60875 1173 60884 1207
rect 60832 1164 60884 1173
rect 61568 1207 61620 1216
rect 61568 1173 61577 1207
rect 61577 1173 61611 1207
rect 61611 1173 61620 1207
rect 61568 1164 61620 1173
rect 62304 1207 62356 1216
rect 62304 1173 62313 1207
rect 62313 1173 62347 1207
rect 62347 1173 62356 1207
rect 62304 1164 62356 1173
rect 63776 1207 63828 1216
rect 63776 1173 63785 1207
rect 63785 1173 63819 1207
rect 63819 1173 63828 1207
rect 63776 1164 63828 1173
rect 64512 1207 64564 1216
rect 64512 1173 64521 1207
rect 64521 1173 64555 1207
rect 64555 1173 64564 1207
rect 64512 1164 64564 1173
rect 66168 1207 66220 1216
rect 66168 1173 66177 1207
rect 66177 1173 66211 1207
rect 66211 1173 66220 1207
rect 66168 1164 66220 1173
rect 82728 1343 82780 1352
rect 82728 1309 82737 1343
rect 82737 1309 82771 1343
rect 82771 1309 82780 1343
rect 82728 1300 82780 1309
rect 85028 1343 85080 1352
rect 85028 1309 85037 1343
rect 85037 1309 85071 1343
rect 85071 1309 85080 1343
rect 85028 1300 85080 1309
rect 85304 1343 85356 1352
rect 85304 1309 85313 1343
rect 85313 1309 85347 1343
rect 85347 1309 85356 1343
rect 85304 1300 85356 1309
rect 86776 1343 86828 1352
rect 86776 1309 86785 1343
rect 86785 1309 86819 1343
rect 86819 1309 86828 1343
rect 86776 1300 86828 1309
rect 87052 1343 87104 1352
rect 87052 1309 87061 1343
rect 87061 1309 87095 1343
rect 87095 1309 87104 1343
rect 87052 1300 87104 1309
rect 88524 1368 88576 1420
rect 88340 1300 88392 1352
rect 89076 1343 89128 1352
rect 89076 1309 89085 1343
rect 89085 1309 89119 1343
rect 89119 1309 89128 1343
rect 89076 1300 89128 1309
rect 89536 1368 89588 1420
rect 98276 1368 98328 1420
rect 89260 1300 89312 1352
rect 90456 1343 90508 1352
rect 90456 1309 90465 1343
rect 90465 1309 90499 1343
rect 90499 1309 90508 1343
rect 90456 1300 90508 1309
rect 92020 1343 92072 1352
rect 92020 1309 92029 1343
rect 92029 1309 92063 1343
rect 92063 1309 92072 1343
rect 92020 1300 92072 1309
rect 93308 1343 93360 1352
rect 93308 1309 93317 1343
rect 93317 1309 93351 1343
rect 93351 1309 93360 1343
rect 93308 1300 93360 1309
rect 94872 1343 94924 1352
rect 94872 1309 94881 1343
rect 94881 1309 94915 1343
rect 94915 1309 94924 1343
rect 94872 1300 94924 1309
rect 94964 1343 95016 1352
rect 94964 1309 94973 1343
rect 94973 1309 95007 1343
rect 95007 1309 95016 1343
rect 94964 1300 95016 1309
rect 96620 1300 96672 1352
rect 97172 1300 97224 1352
rect 98552 1343 98604 1352
rect 98552 1309 98561 1343
rect 98561 1309 98595 1343
rect 98595 1309 98604 1343
rect 98552 1300 98604 1309
rect 99564 1368 99616 1420
rect 99840 1300 99892 1352
rect 100116 1343 100168 1352
rect 100116 1309 100125 1343
rect 100125 1309 100159 1343
rect 100159 1309 100168 1343
rect 100116 1300 100168 1309
rect 84476 1232 84528 1284
rect 103244 1411 103296 1420
rect 103244 1377 103253 1411
rect 103253 1377 103287 1411
rect 103287 1377 103296 1411
rect 103244 1368 103296 1377
rect 100576 1232 100628 1284
rect 103888 1343 103940 1352
rect 103888 1309 103897 1343
rect 103897 1309 103931 1343
rect 103931 1309 103940 1343
rect 103888 1300 103940 1309
rect 104716 1300 104768 1352
rect 105636 1343 105688 1352
rect 105636 1309 105645 1343
rect 105645 1309 105679 1343
rect 105679 1309 105688 1343
rect 105636 1300 105688 1309
rect 106188 1300 106240 1352
rect 107752 1343 107804 1352
rect 107752 1309 107761 1343
rect 107761 1309 107795 1343
rect 107795 1309 107804 1343
rect 107752 1300 107804 1309
rect 108396 1343 108448 1352
rect 108396 1309 108405 1343
rect 108405 1309 108439 1343
rect 108439 1309 108448 1343
rect 108396 1300 108448 1309
rect 109040 1343 109092 1352
rect 109040 1309 109049 1343
rect 109049 1309 109083 1343
rect 109083 1309 109092 1343
rect 109040 1300 109092 1309
rect 109224 1300 109276 1352
rect 110052 1343 110104 1352
rect 110052 1309 110061 1343
rect 110061 1309 110095 1343
rect 110095 1309 110104 1343
rect 110052 1300 110104 1309
rect 110972 1368 111024 1420
rect 149244 1368 149296 1420
rect 90640 1207 90692 1216
rect 90640 1173 90649 1207
rect 90649 1173 90683 1207
rect 90683 1173 90692 1207
rect 90640 1164 90692 1173
rect 92204 1207 92256 1216
rect 92204 1173 92213 1207
rect 92213 1173 92247 1207
rect 92247 1173 92256 1207
rect 92204 1164 92256 1173
rect 93492 1207 93544 1216
rect 93492 1173 93501 1207
rect 93501 1173 93535 1207
rect 93535 1173 93544 1207
rect 93492 1164 93544 1173
rect 96528 1164 96580 1216
rect 97080 1207 97132 1216
rect 97080 1173 97089 1207
rect 97089 1173 97123 1207
rect 97123 1173 97132 1207
rect 97080 1164 97132 1173
rect 98460 1164 98512 1216
rect 100024 1164 100076 1216
rect 104256 1232 104308 1284
rect 104808 1232 104860 1284
rect 104624 1164 104676 1216
rect 105452 1207 105504 1216
rect 105452 1173 105461 1207
rect 105461 1173 105495 1207
rect 105495 1173 105504 1207
rect 105452 1164 105504 1173
rect 107476 1232 107528 1284
rect 106280 1164 106332 1216
rect 108120 1232 108172 1284
rect 110788 1343 110840 1352
rect 110788 1309 110797 1343
rect 110797 1309 110831 1343
rect 110831 1309 110840 1343
rect 110788 1300 110840 1309
rect 111524 1343 111576 1352
rect 111524 1309 111533 1343
rect 111533 1309 111567 1343
rect 111567 1309 111576 1343
rect 111524 1300 111576 1309
rect 112904 1343 112956 1352
rect 112904 1309 112913 1343
rect 112913 1309 112947 1343
rect 112947 1309 112956 1343
rect 112904 1300 112956 1309
rect 113088 1300 113140 1352
rect 108856 1207 108908 1216
rect 108856 1173 108865 1207
rect 108865 1173 108899 1207
rect 108899 1173 108908 1207
rect 108856 1164 108908 1173
rect 109868 1207 109920 1216
rect 109868 1173 109877 1207
rect 109877 1173 109911 1207
rect 109911 1173 109920 1207
rect 109868 1164 109920 1173
rect 111340 1207 111392 1216
rect 111340 1173 111349 1207
rect 111349 1173 111383 1207
rect 111383 1173 111392 1207
rect 111340 1164 111392 1173
rect 112720 1207 112772 1216
rect 112720 1173 112729 1207
rect 112729 1173 112763 1207
rect 112763 1173 112772 1207
rect 112720 1164 112772 1173
rect 112996 1232 113048 1284
rect 113364 1232 113416 1284
rect 113548 1343 113600 1352
rect 113548 1309 113557 1343
rect 113557 1309 113591 1343
rect 113591 1309 113600 1343
rect 113548 1300 113600 1309
rect 113640 1300 113692 1352
rect 114192 1343 114244 1352
rect 114192 1309 114201 1343
rect 114201 1309 114235 1343
rect 114235 1309 114244 1343
rect 114192 1300 114244 1309
rect 115204 1343 115256 1352
rect 115204 1309 115213 1343
rect 115213 1309 115247 1343
rect 115247 1309 115256 1343
rect 115204 1300 115256 1309
rect 115756 1300 115808 1352
rect 116676 1343 116728 1352
rect 116676 1309 116685 1343
rect 116685 1309 116719 1343
rect 116719 1309 116728 1343
rect 116676 1300 116728 1309
rect 118056 1343 118108 1352
rect 118056 1309 118065 1343
rect 118065 1309 118099 1343
rect 118099 1309 118108 1343
rect 118056 1300 118108 1309
rect 118700 1343 118752 1352
rect 118700 1309 118709 1343
rect 118709 1309 118743 1343
rect 118743 1309 118752 1343
rect 118700 1300 118752 1309
rect 119344 1343 119396 1352
rect 119344 1309 119353 1343
rect 119353 1309 119387 1343
rect 119387 1309 119396 1343
rect 119344 1300 119396 1309
rect 120356 1343 120408 1352
rect 120356 1309 120365 1343
rect 120365 1309 120399 1343
rect 120399 1309 120408 1343
rect 120356 1300 120408 1309
rect 121092 1343 121144 1352
rect 121092 1309 121101 1343
rect 121101 1309 121135 1343
rect 121135 1309 121144 1343
rect 121092 1300 121144 1309
rect 121184 1300 121236 1352
rect 122932 1343 122984 1352
rect 122932 1309 122941 1343
rect 122941 1309 122975 1343
rect 122975 1309 122984 1343
rect 122932 1300 122984 1309
rect 123760 1343 123812 1352
rect 123760 1309 123769 1343
rect 123769 1309 123803 1343
rect 123803 1309 123812 1343
rect 123760 1300 123812 1309
rect 125416 1343 125468 1352
rect 125416 1309 125425 1343
rect 125425 1309 125459 1343
rect 125459 1309 125468 1343
rect 125416 1300 125468 1309
rect 127072 1300 127124 1352
rect 128268 1343 128320 1352
rect 128268 1309 128277 1343
rect 128277 1309 128311 1343
rect 128311 1309 128320 1343
rect 128268 1300 128320 1309
rect 128452 1343 128504 1352
rect 128452 1309 128461 1343
rect 128461 1309 128495 1343
rect 128495 1309 128504 1343
rect 128452 1300 128504 1309
rect 128636 1343 128688 1352
rect 128636 1309 128645 1343
rect 128645 1309 128679 1343
rect 128679 1309 128688 1343
rect 128636 1300 128688 1309
rect 129096 1343 129148 1352
rect 129096 1309 129105 1343
rect 129105 1309 129139 1343
rect 129139 1309 129148 1343
rect 129096 1300 129148 1309
rect 130660 1343 130712 1352
rect 130660 1309 130669 1343
rect 130669 1309 130703 1343
rect 130703 1309 130712 1343
rect 130660 1300 130712 1309
rect 132592 1300 132644 1352
rect 132776 1300 132828 1352
rect 133144 1343 133196 1352
rect 133144 1309 133153 1343
rect 133153 1309 133187 1343
rect 133187 1309 133196 1343
rect 133144 1300 133196 1309
rect 133880 1300 133932 1352
rect 134064 1300 134116 1352
rect 138756 1343 138808 1352
rect 138756 1309 138765 1343
rect 138765 1309 138799 1343
rect 138799 1309 138808 1343
rect 138756 1300 138808 1309
rect 138848 1300 138900 1352
rect 140688 1343 140740 1352
rect 140688 1309 140697 1343
rect 140697 1309 140731 1343
rect 140731 1309 140740 1343
rect 140688 1300 140740 1309
rect 140780 1300 140832 1352
rect 141976 1343 142028 1352
rect 141976 1309 141985 1343
rect 141985 1309 142019 1343
rect 142019 1309 142028 1343
rect 141976 1300 142028 1309
rect 142068 1300 142120 1352
rect 143540 1300 143592 1352
rect 144552 1343 144604 1352
rect 144552 1309 144561 1343
rect 144561 1309 144595 1343
rect 144595 1309 144604 1343
rect 144552 1300 144604 1309
rect 145840 1343 145892 1352
rect 145840 1309 145849 1343
rect 145849 1309 145883 1343
rect 145883 1309 145892 1343
rect 145840 1300 145892 1309
rect 146208 1300 146260 1352
rect 147128 1343 147180 1352
rect 147128 1309 147137 1343
rect 147137 1309 147171 1343
rect 147171 1309 147180 1343
rect 147128 1300 147180 1309
rect 148416 1343 148468 1352
rect 148416 1309 148425 1343
rect 148425 1309 148459 1343
rect 148459 1309 148468 1343
rect 148416 1300 148468 1309
rect 148508 1300 148560 1352
rect 149704 1343 149756 1352
rect 149704 1309 149713 1343
rect 149713 1309 149747 1343
rect 149747 1309 149756 1343
rect 149704 1300 149756 1309
rect 150992 1343 151044 1352
rect 150992 1309 151001 1343
rect 151001 1309 151035 1343
rect 151035 1309 151044 1343
rect 150992 1300 151044 1309
rect 151636 1343 151688 1352
rect 151636 1309 151645 1343
rect 151645 1309 151679 1343
rect 151679 1309 151688 1343
rect 151636 1300 151688 1309
rect 152280 1343 152332 1352
rect 152280 1309 152289 1343
rect 152289 1309 152323 1343
rect 152323 1309 152332 1343
rect 152280 1300 152332 1309
rect 153200 1300 153252 1352
rect 113272 1164 113324 1216
rect 115020 1207 115072 1216
rect 115020 1173 115029 1207
rect 115029 1173 115063 1207
rect 115063 1173 115072 1207
rect 115020 1164 115072 1173
rect 123576 1232 123628 1284
rect 148784 1232 148836 1284
rect 115848 1164 115900 1216
rect 117228 1164 117280 1216
rect 118516 1207 118568 1216
rect 118516 1173 118525 1207
rect 118525 1173 118559 1207
rect 118559 1173 118568 1207
rect 118516 1164 118568 1173
rect 119252 1164 119304 1216
rect 120172 1207 120224 1216
rect 120172 1173 120181 1207
rect 120181 1173 120215 1207
rect 120215 1173 120224 1207
rect 120172 1164 120224 1173
rect 120816 1164 120868 1216
rect 121828 1207 121880 1216
rect 121828 1173 121837 1207
rect 121837 1173 121871 1207
rect 121871 1173 121880 1207
rect 121828 1164 121880 1173
rect 123116 1207 123168 1216
rect 123116 1173 123125 1207
rect 123125 1173 123159 1207
rect 123159 1173 123168 1207
rect 123116 1164 123168 1173
rect 123944 1207 123996 1216
rect 123944 1173 123953 1207
rect 123953 1173 123987 1207
rect 123987 1173 123996 1207
rect 123944 1164 123996 1173
rect 125324 1164 125376 1216
rect 126796 1164 126848 1216
rect 129280 1207 129332 1216
rect 129280 1173 129289 1207
rect 129289 1173 129323 1207
rect 129323 1173 129332 1207
rect 129280 1164 129332 1173
rect 130844 1207 130896 1216
rect 130844 1173 130853 1207
rect 130853 1173 130887 1207
rect 130887 1173 130896 1207
rect 130844 1164 130896 1173
rect 132132 1207 132184 1216
rect 132132 1173 132141 1207
rect 132141 1173 132175 1207
rect 132175 1173 132184 1207
rect 132132 1164 132184 1173
rect 137928 1164 137980 1216
rect 140872 1164 140924 1216
rect 141884 1164 141936 1216
rect 143080 1207 143132 1216
rect 143080 1173 143089 1207
rect 143089 1173 143123 1207
rect 143123 1173 143132 1207
rect 143080 1164 143132 1173
rect 143816 1164 143868 1216
rect 144368 1207 144420 1216
rect 144368 1173 144377 1207
rect 144377 1173 144411 1207
rect 144411 1173 144420 1207
rect 144368 1164 144420 1173
rect 145656 1207 145708 1216
rect 145656 1173 145665 1207
rect 145665 1173 145699 1207
rect 145699 1173 145708 1207
rect 145656 1164 145708 1173
rect 146116 1164 146168 1216
rect 146392 1164 146444 1216
rect 148232 1207 148284 1216
rect 148232 1173 148241 1207
rect 148241 1173 148275 1207
rect 148275 1173 148284 1207
rect 148232 1164 148284 1173
rect 150624 1232 150676 1284
rect 150716 1164 150768 1216
rect 150900 1164 150952 1216
rect 153292 1232 153344 1284
rect 152096 1207 152148 1216
rect 152096 1173 152105 1207
rect 152105 1173 152139 1207
rect 152139 1173 152148 1207
rect 152096 1164 152148 1173
rect 154212 1343 154264 1352
rect 154212 1309 154221 1343
rect 154221 1309 154255 1343
rect 154255 1309 154264 1343
rect 154212 1300 154264 1309
rect 154580 1300 154632 1352
rect 156512 1368 156564 1420
rect 157064 1368 157116 1420
rect 158168 1368 158220 1420
rect 159088 1368 159140 1420
rect 156144 1300 156196 1352
rect 156236 1232 156288 1284
rect 156052 1164 156104 1216
rect 159272 1300 159324 1352
rect 160376 1368 160428 1420
rect 164148 1368 164200 1420
rect 168104 1368 168156 1420
rect 171692 1411 171744 1420
rect 171692 1377 171701 1411
rect 171701 1377 171735 1411
rect 171735 1377 171744 1411
rect 171692 1368 171744 1377
rect 190920 1368 190972 1420
rect 160192 1343 160244 1352
rect 160192 1309 160201 1343
rect 160201 1309 160235 1343
rect 160235 1309 160244 1343
rect 160192 1300 160244 1309
rect 161480 1300 161532 1352
rect 163136 1300 163188 1352
rect 163780 1300 163832 1352
rect 164424 1300 164476 1352
rect 164516 1343 164568 1352
rect 164516 1309 164525 1343
rect 164525 1309 164559 1343
rect 164559 1309 164568 1343
rect 164516 1300 164568 1309
rect 167184 1343 167236 1352
rect 167184 1309 167193 1343
rect 167193 1309 167227 1343
rect 167227 1309 167236 1343
rect 167184 1300 167236 1309
rect 168012 1300 168064 1352
rect 172244 1343 172296 1352
rect 172244 1309 172253 1343
rect 172253 1309 172287 1343
rect 172287 1309 172296 1343
rect 172244 1300 172296 1309
rect 172520 1343 172572 1352
rect 172520 1309 172529 1343
rect 172529 1309 172563 1343
rect 172563 1309 172572 1343
rect 172520 1300 172572 1309
rect 173808 1300 173860 1352
rect 174268 1343 174320 1352
rect 174268 1309 174277 1343
rect 174277 1309 174311 1343
rect 174311 1309 174320 1343
rect 174268 1300 174320 1309
rect 175188 1300 175240 1352
rect 176844 1343 176896 1352
rect 176844 1309 176853 1343
rect 176853 1309 176887 1343
rect 176887 1309 176896 1343
rect 176844 1300 176896 1309
rect 178408 1300 178460 1352
rect 179420 1343 179472 1352
rect 179420 1309 179429 1343
rect 179429 1309 179463 1343
rect 179463 1309 179472 1343
rect 179420 1300 179472 1309
rect 182548 1343 182600 1352
rect 182548 1309 182557 1343
rect 182557 1309 182591 1343
rect 182591 1309 182600 1343
rect 182548 1300 182600 1309
rect 182824 1343 182876 1352
rect 182824 1309 182833 1343
rect 182833 1309 182867 1343
rect 182867 1309 182876 1343
rect 182824 1300 182876 1309
rect 184296 1343 184348 1352
rect 184296 1309 184305 1343
rect 184305 1309 184339 1343
rect 184339 1309 184348 1343
rect 184296 1300 184348 1309
rect 184572 1343 184624 1352
rect 184572 1309 184581 1343
rect 184581 1309 184615 1343
rect 184615 1309 184624 1343
rect 184572 1300 184624 1309
rect 185584 1300 185636 1352
rect 187148 1343 187200 1352
rect 187148 1309 187157 1343
rect 187157 1309 187191 1343
rect 187191 1309 187200 1343
rect 187148 1300 187200 1309
rect 188528 1300 188580 1352
rect 189724 1343 189776 1352
rect 189724 1309 189733 1343
rect 189733 1309 189767 1343
rect 189767 1309 189776 1343
rect 189724 1300 189776 1309
rect 191104 1343 191156 1352
rect 191104 1309 191113 1343
rect 191113 1309 191147 1343
rect 191147 1309 191156 1343
rect 191104 1300 191156 1309
rect 202052 1368 202104 1420
rect 202328 1411 202380 1420
rect 202328 1377 202337 1411
rect 202337 1377 202371 1411
rect 202371 1377 202380 1411
rect 202328 1368 202380 1377
rect 205824 1411 205876 1420
rect 205824 1377 205833 1411
rect 205833 1377 205867 1411
rect 205867 1377 205876 1411
rect 205824 1368 205876 1377
rect 193220 1300 193272 1352
rect 193312 1343 193364 1352
rect 193312 1309 193321 1343
rect 193321 1309 193355 1343
rect 193355 1309 193364 1343
rect 193312 1300 193364 1309
rect 194600 1343 194652 1352
rect 194600 1309 194609 1343
rect 194609 1309 194643 1343
rect 194643 1309 194652 1343
rect 194600 1300 194652 1309
rect 196532 1300 196584 1352
rect 197452 1300 197504 1352
rect 197912 1343 197964 1352
rect 197912 1309 197921 1343
rect 197921 1309 197955 1343
rect 197955 1309 197964 1343
rect 197912 1300 197964 1309
rect 199752 1343 199804 1352
rect 199752 1309 199761 1343
rect 199761 1309 199795 1343
rect 199795 1309 199804 1343
rect 199752 1300 199804 1309
rect 158812 1232 158864 1284
rect 156972 1164 157024 1216
rect 157708 1164 157760 1216
rect 161388 1232 161440 1284
rect 179512 1232 179564 1284
rect 180524 1275 180576 1284
rect 180524 1241 180533 1275
rect 180533 1241 180567 1275
rect 180567 1241 180576 1275
rect 180524 1232 180576 1241
rect 181812 1275 181864 1284
rect 181812 1241 181821 1275
rect 181821 1241 181855 1275
rect 181855 1241 181864 1275
rect 181812 1232 181864 1241
rect 197268 1232 197320 1284
rect 201316 1300 201368 1352
rect 206560 1343 206612 1352
rect 206560 1309 206569 1343
rect 206569 1309 206603 1343
rect 206603 1309 206612 1343
rect 206560 1300 206612 1309
rect 207664 1343 207716 1352
rect 207664 1309 207673 1343
rect 207673 1309 207707 1343
rect 207707 1309 207716 1343
rect 207664 1300 207716 1309
rect 208308 1343 208360 1352
rect 208308 1309 208317 1343
rect 208317 1309 208351 1343
rect 208351 1309 208360 1343
rect 208308 1300 208360 1309
rect 208952 1343 209004 1352
rect 208952 1309 208961 1343
rect 208961 1309 208995 1343
rect 208995 1309 209004 1343
rect 208952 1300 209004 1309
rect 209780 1300 209832 1352
rect 210884 1343 210936 1352
rect 210884 1309 210893 1343
rect 210893 1309 210927 1343
rect 210927 1309 210936 1343
rect 210884 1300 210936 1309
rect 211528 1343 211580 1352
rect 211528 1309 211537 1343
rect 211537 1309 211571 1343
rect 211571 1309 211580 1343
rect 211528 1300 211580 1309
rect 212264 1300 212316 1352
rect 161296 1207 161348 1216
rect 161296 1173 161305 1207
rect 161305 1173 161339 1207
rect 161339 1173 161348 1207
rect 161296 1164 161348 1173
rect 162492 1207 162544 1216
rect 162492 1173 162501 1207
rect 162501 1173 162535 1207
rect 162535 1173 162544 1207
rect 162492 1164 162544 1173
rect 164700 1207 164752 1216
rect 164700 1173 164709 1207
rect 164709 1173 164743 1207
rect 164743 1173 164752 1207
rect 164700 1164 164752 1173
rect 168012 1207 168064 1216
rect 168012 1173 168021 1207
rect 168021 1173 168055 1207
rect 168055 1173 168064 1207
rect 168012 1164 168064 1173
rect 169024 1207 169076 1216
rect 169024 1173 169033 1207
rect 169033 1173 169067 1207
rect 169067 1173 169076 1207
rect 169024 1164 169076 1173
rect 181904 1207 181956 1216
rect 181904 1173 181913 1207
rect 181913 1173 181947 1207
rect 181947 1173 181956 1207
rect 181904 1164 181956 1173
rect 192668 1207 192720 1216
rect 192668 1173 192677 1207
rect 192677 1173 192711 1207
rect 192711 1173 192720 1207
rect 192668 1164 192720 1173
rect 192944 1164 192996 1216
rect 193680 1164 193732 1216
rect 195796 1207 195848 1216
rect 195796 1173 195805 1207
rect 195805 1173 195839 1207
rect 195839 1173 195848 1207
rect 195796 1164 195848 1173
rect 196624 1164 196676 1216
rect 201684 1232 201736 1284
rect 199936 1207 199988 1216
rect 199936 1173 199945 1207
rect 199945 1173 199979 1207
rect 199979 1173 199988 1207
rect 199936 1164 199988 1173
rect 200672 1207 200724 1216
rect 200672 1173 200681 1207
rect 200681 1173 200715 1207
rect 200715 1173 200724 1207
rect 200672 1164 200724 1173
rect 201224 1164 201276 1216
rect 203340 1207 203392 1216
rect 203340 1173 203349 1207
rect 203349 1173 203383 1207
rect 203383 1173 203392 1207
rect 203340 1164 203392 1173
rect 206376 1207 206428 1216
rect 206376 1173 206385 1207
rect 206385 1173 206419 1207
rect 206419 1173 206428 1207
rect 206376 1164 206428 1173
rect 207480 1207 207532 1216
rect 207480 1173 207489 1207
rect 207489 1173 207523 1207
rect 207523 1173 207532 1207
rect 207480 1164 207532 1173
rect 209964 1232 210016 1284
rect 209872 1164 209924 1216
rect 210332 1164 210384 1216
rect 212540 1232 212592 1284
rect 224776 1436 224828 1488
rect 227812 1436 227864 1488
rect 228824 1504 228876 1556
rect 232596 1504 232648 1556
rect 236552 1504 236604 1556
rect 257068 1504 257120 1556
rect 239496 1436 239548 1488
rect 256976 1436 257028 1488
rect 225420 1368 225472 1420
rect 227076 1368 227128 1420
rect 228180 1368 228232 1420
rect 232504 1368 232556 1420
rect 235448 1368 235500 1420
rect 237196 1368 237248 1420
rect 213460 1343 213512 1352
rect 213460 1309 213469 1343
rect 213469 1309 213503 1343
rect 213503 1309 213512 1343
rect 213460 1300 213512 1309
rect 213736 1300 213788 1352
rect 214472 1300 214524 1352
rect 214564 1232 214616 1284
rect 215116 1232 215168 1284
rect 216680 1343 216732 1352
rect 216680 1309 216689 1343
rect 216689 1309 216723 1343
rect 216723 1309 216732 1343
rect 216680 1300 216732 1309
rect 217784 1343 217836 1352
rect 217784 1309 217793 1343
rect 217793 1309 217827 1343
rect 217827 1309 217836 1343
rect 217784 1300 217836 1309
rect 218152 1300 218204 1352
rect 211804 1164 211856 1216
rect 213828 1164 213880 1216
rect 214380 1164 214432 1216
rect 215208 1207 215260 1216
rect 215208 1173 215217 1207
rect 215217 1173 215251 1207
rect 215251 1173 215260 1207
rect 215208 1164 215260 1173
rect 215576 1164 215628 1216
rect 217600 1232 217652 1284
rect 218060 1275 218112 1284
rect 218060 1241 218069 1275
rect 218069 1241 218103 1275
rect 218103 1241 218112 1275
rect 218060 1232 218112 1241
rect 217416 1164 217468 1216
rect 218980 1275 219032 1284
rect 218980 1241 218989 1275
rect 218989 1241 219023 1275
rect 219023 1241 219032 1275
rect 218980 1232 219032 1241
rect 219440 1232 219492 1284
rect 221188 1343 221240 1352
rect 221188 1309 221197 1343
rect 221197 1309 221231 1343
rect 221231 1309 221240 1343
rect 221188 1300 221240 1309
rect 220728 1232 220780 1284
rect 222200 1300 222252 1352
rect 223764 1343 223816 1352
rect 223764 1309 223773 1343
rect 223773 1309 223807 1343
rect 223807 1309 223816 1343
rect 223764 1300 223816 1309
rect 222292 1232 222344 1284
rect 226616 1300 226668 1352
rect 226892 1343 226944 1352
rect 226892 1309 226901 1343
rect 226901 1309 226935 1343
rect 226935 1309 226944 1343
rect 226892 1300 226944 1309
rect 228364 1300 228416 1352
rect 229284 1300 229336 1352
rect 229652 1343 229704 1352
rect 229652 1309 229661 1343
rect 229661 1309 229695 1343
rect 229695 1309 229704 1343
rect 229652 1300 229704 1309
rect 230664 1343 230716 1352
rect 230664 1309 230673 1343
rect 230673 1309 230707 1343
rect 230707 1309 230716 1343
rect 230664 1300 230716 1309
rect 232320 1343 232372 1352
rect 232320 1309 232329 1343
rect 232329 1309 232363 1343
rect 232363 1309 232372 1343
rect 232320 1300 232372 1309
rect 233240 1343 233292 1352
rect 233240 1309 233249 1343
rect 233249 1309 233283 1343
rect 233283 1309 233292 1343
rect 233240 1300 233292 1309
rect 233976 1343 234028 1352
rect 233976 1309 233985 1343
rect 233985 1309 234019 1343
rect 234019 1309 234028 1343
rect 233976 1300 234028 1309
rect 234712 1343 234764 1352
rect 234712 1309 234721 1343
rect 234721 1309 234755 1343
rect 234755 1309 234764 1343
rect 234712 1300 234764 1309
rect 236000 1343 236052 1352
rect 236000 1309 236009 1343
rect 236009 1309 236043 1343
rect 236043 1309 236052 1343
rect 236000 1300 236052 1309
rect 239956 1411 240008 1420
rect 239956 1377 239965 1411
rect 239965 1377 239999 1411
rect 239999 1377 240008 1411
rect 239956 1368 240008 1377
rect 257712 1411 257764 1420
rect 257712 1377 257721 1411
rect 257721 1377 257755 1411
rect 257755 1377 257764 1411
rect 257712 1368 257764 1377
rect 267740 1368 267792 1420
rect 240968 1343 241020 1352
rect 240968 1309 240977 1343
rect 240977 1309 241011 1343
rect 241011 1309 241020 1343
rect 240968 1300 241020 1309
rect 241060 1300 241112 1352
rect 241980 1300 242032 1352
rect 243820 1343 243872 1352
rect 243820 1309 243829 1343
rect 243829 1309 243863 1343
rect 243863 1309 243872 1343
rect 243820 1300 243872 1309
rect 244924 1300 244976 1352
rect 246212 1300 246264 1352
rect 246488 1300 246540 1352
rect 224040 1275 224092 1284
rect 224040 1241 224049 1275
rect 224049 1241 224083 1275
rect 224083 1241 224092 1275
rect 224040 1232 224092 1241
rect 226248 1232 226300 1284
rect 230204 1232 230256 1284
rect 230388 1232 230440 1284
rect 237380 1232 237432 1284
rect 248328 1232 248380 1284
rect 248512 1300 248564 1352
rect 248972 1343 249024 1352
rect 248972 1309 248981 1343
rect 248981 1309 249015 1343
rect 249015 1309 249024 1343
rect 248972 1300 249024 1309
rect 250168 1275 250220 1284
rect 250168 1241 250177 1275
rect 250177 1241 250211 1275
rect 250211 1241 250220 1275
rect 250168 1232 250220 1241
rect 219624 1207 219676 1216
rect 219624 1173 219633 1207
rect 219633 1173 219667 1207
rect 219667 1173 219676 1207
rect 219624 1164 219676 1173
rect 220360 1207 220412 1216
rect 220360 1173 220369 1207
rect 220369 1173 220403 1207
rect 220403 1173 220412 1207
rect 220360 1164 220412 1173
rect 220912 1164 220964 1216
rect 223120 1164 223172 1216
rect 225052 1164 225104 1216
rect 229100 1207 229152 1216
rect 229100 1173 229109 1207
rect 229109 1173 229143 1207
rect 229143 1173 229152 1207
rect 229100 1164 229152 1173
rect 229836 1207 229888 1216
rect 229836 1173 229845 1207
rect 229845 1173 229879 1207
rect 229879 1173 229888 1207
rect 229836 1164 229888 1173
rect 230848 1207 230900 1216
rect 230848 1173 230857 1207
rect 230857 1173 230891 1207
rect 230891 1173 230900 1207
rect 230848 1164 230900 1173
rect 233424 1207 233476 1216
rect 233424 1173 233433 1207
rect 233433 1173 233467 1207
rect 233467 1173 233476 1207
rect 233424 1164 233476 1173
rect 234160 1207 234212 1216
rect 234160 1173 234169 1207
rect 234169 1173 234203 1207
rect 234203 1173 234212 1207
rect 234160 1164 234212 1173
rect 234896 1207 234948 1216
rect 234896 1173 234905 1207
rect 234905 1173 234939 1207
rect 234939 1173 234948 1207
rect 234896 1164 234948 1173
rect 248052 1207 248104 1216
rect 248052 1173 248061 1207
rect 248061 1173 248095 1207
rect 248095 1173 248104 1207
rect 248052 1164 248104 1173
rect 250260 1207 250312 1216
rect 250260 1173 250269 1207
rect 250269 1173 250303 1207
rect 250303 1173 250312 1207
rect 250260 1164 250312 1173
rect 251548 1343 251600 1352
rect 251548 1309 251557 1343
rect 251557 1309 251591 1343
rect 251591 1309 251600 1343
rect 251548 1300 251600 1309
rect 251824 1343 251876 1352
rect 251824 1309 251833 1343
rect 251833 1309 251867 1343
rect 251867 1309 251876 1343
rect 251824 1300 251876 1309
rect 253480 1300 253532 1352
rect 254124 1343 254176 1352
rect 254124 1309 254133 1343
rect 254133 1309 254167 1343
rect 254167 1309 254176 1343
rect 254124 1300 254176 1309
rect 255228 1300 255280 1352
rect 256516 1300 256568 1352
rect 257804 1300 257856 1352
rect 257988 1300 258040 1352
rect 257436 1232 257488 1284
rect 260288 1343 260340 1352
rect 260288 1309 260297 1343
rect 260297 1309 260331 1343
rect 260331 1309 260340 1343
rect 260288 1300 260340 1309
rect 261576 1343 261628 1352
rect 261576 1309 261585 1343
rect 261585 1309 261619 1343
rect 261619 1309 261628 1343
rect 261576 1300 261628 1309
rect 262312 1343 262364 1352
rect 262312 1309 262321 1343
rect 262321 1309 262355 1343
rect 262355 1309 262364 1343
rect 262312 1300 262364 1309
rect 263048 1343 263100 1352
rect 263048 1309 263057 1343
rect 263057 1309 263091 1343
rect 263091 1309 263100 1343
rect 263048 1300 263100 1309
rect 264152 1343 264204 1352
rect 264152 1309 264161 1343
rect 264161 1309 264195 1343
rect 264195 1309 264204 1343
rect 264152 1300 264204 1309
rect 265164 1343 265216 1352
rect 265164 1309 265173 1343
rect 265173 1309 265207 1343
rect 265207 1309 265216 1343
rect 265164 1300 265216 1309
rect 265900 1343 265952 1352
rect 265900 1309 265909 1343
rect 265909 1309 265943 1343
rect 265943 1309 265952 1343
rect 265900 1300 265952 1309
rect 266728 1343 266780 1352
rect 266728 1309 266737 1343
rect 266737 1309 266771 1343
rect 266771 1309 266780 1343
rect 266728 1300 266780 1309
rect 267832 1300 267884 1352
rect 268200 1343 268252 1352
rect 268200 1309 268209 1343
rect 268209 1309 268243 1343
rect 268243 1309 268252 1343
rect 268200 1300 268252 1309
rect 269212 1300 269264 1352
rect 269856 1300 269908 1352
rect 269948 1300 270000 1352
rect 268936 1232 268988 1284
rect 271788 1232 271840 1284
rect 260472 1207 260524 1216
rect 260472 1173 260481 1207
rect 260481 1173 260515 1207
rect 260515 1173 260524 1207
rect 260472 1164 260524 1173
rect 261760 1207 261812 1216
rect 261760 1173 261769 1207
rect 261769 1173 261803 1207
rect 261803 1173 261812 1207
rect 261760 1164 261812 1173
rect 262496 1207 262548 1216
rect 262496 1173 262505 1207
rect 262505 1173 262539 1207
rect 262539 1173 262548 1207
rect 262496 1164 262548 1173
rect 263232 1207 263284 1216
rect 263232 1173 263241 1207
rect 263241 1173 263275 1207
rect 263275 1173 263284 1207
rect 263232 1164 263284 1173
rect 264336 1207 264388 1216
rect 264336 1173 264345 1207
rect 264345 1173 264379 1207
rect 264379 1173 264388 1207
rect 264336 1164 264388 1173
rect 265348 1207 265400 1216
rect 265348 1173 265357 1207
rect 265357 1173 265391 1207
rect 265391 1173 265400 1207
rect 265348 1164 265400 1173
rect 266084 1207 266136 1216
rect 266084 1173 266093 1207
rect 266093 1173 266127 1207
rect 266127 1173 266136 1207
rect 266084 1164 266136 1173
rect 266912 1207 266964 1216
rect 266912 1173 266921 1207
rect 266921 1173 266955 1207
rect 266955 1173 266964 1207
rect 266912 1164 266964 1173
rect 267648 1207 267700 1216
rect 267648 1173 267657 1207
rect 267657 1173 267691 1207
rect 267691 1173 267700 1207
rect 267648 1164 267700 1173
rect 268384 1207 268436 1216
rect 268384 1173 268393 1207
rect 268393 1173 268427 1207
rect 268427 1173 268436 1207
rect 268384 1164 268436 1173
rect 270316 1207 270368 1216
rect 270316 1173 270325 1207
rect 270325 1173 270359 1207
rect 270359 1173 270368 1207
rect 270316 1164 270368 1173
rect 68546 1062 68598 1114
rect 68610 1062 68662 1114
rect 68674 1062 68726 1114
rect 68738 1062 68790 1114
rect 68802 1062 68854 1114
rect 136143 1062 136195 1114
rect 136207 1062 136259 1114
rect 136271 1062 136323 1114
rect 136335 1062 136387 1114
rect 136399 1062 136451 1114
rect 203740 1062 203792 1114
rect 203804 1062 203856 1114
rect 203868 1062 203920 1114
rect 203932 1062 203984 1114
rect 203996 1062 204048 1114
rect 271337 1062 271389 1114
rect 271401 1062 271453 1114
rect 271465 1062 271517 1114
rect 271529 1062 271581 1114
rect 271593 1062 271645 1114
rect 13544 960 13596 1012
rect 47676 960 47728 1012
rect 69848 960 69900 1012
rect 96712 960 96764 1012
rect 106004 960 106056 1012
rect 108856 960 108908 1012
rect 108948 960 109000 1012
rect 109868 960 109920 1012
rect 141516 960 141568 1012
rect 174268 960 174320 1012
rect 207480 960 207532 1012
rect 210240 960 210292 1012
rect 210332 960 210384 1012
rect 212816 960 212868 1012
rect 217968 960 218020 1012
rect 219624 960 219676 1012
rect 18696 892 18748 944
rect 53196 892 53248 944
rect 82360 892 82412 944
rect 114836 892 114888 944
rect 145656 892 145708 944
rect 147772 892 147824 944
rect 152096 892 152148 944
rect 155868 892 155920 944
rect 17224 824 17276 876
rect 51448 824 51500 876
rect 82636 824 82688 876
rect 115112 824 115164 876
rect 141332 824 141384 876
rect 152464 824 152516 876
rect 152556 824 152608 876
rect 182824 892 182876 944
rect 210976 892 211028 944
rect 216864 892 216916 944
rect 218060 892 218112 944
rect 220084 892 220136 944
rect 158904 824 158956 876
rect 189724 824 189776 876
rect 211160 824 211212 876
rect 219808 824 219860 876
rect 4160 756 4212 808
rect 38752 756 38804 808
rect 81440 756 81492 808
rect 12808 688 12860 740
rect 46296 688 46348 740
rect 76748 688 76800 740
rect 100392 688 100444 740
rect 9680 620 9732 672
rect 43904 620 43956 672
rect 73804 620 73856 672
rect 104256 756 104308 808
rect 109960 756 110012 808
rect 142712 756 142764 808
rect 204260 756 204312 808
rect 213644 756 213696 808
rect 246212 960 246264 1012
rect 265532 960 265584 1012
rect 269028 960 269080 1012
rect 220268 892 220320 944
rect 223580 892 223632 944
rect 224868 892 224920 944
rect 226248 892 226300 944
rect 229744 892 229796 944
rect 254124 892 254176 944
rect 222016 824 222068 876
rect 250260 824 250312 876
rect 221556 756 221608 808
rect 254032 756 254084 808
rect 107200 688 107252 740
rect 108856 688 108908 740
rect 8392 552 8444 604
rect 40224 552 40276 604
rect 75000 552 75052 604
rect 17960 484 18012 536
rect 51816 484 51868 536
rect 101864 552 101916 604
rect 105084 484 105136 536
rect 107568 620 107620 672
rect 112720 688 112772 740
rect 146760 688 146812 740
rect 179420 688 179472 740
rect 207204 688 207256 740
rect 217324 688 217376 740
rect 218888 688 218940 740
rect 221188 688 221240 740
rect 224776 688 224828 740
rect 258356 688 258408 740
rect 143908 620 143960 672
rect 176844 620 176896 672
rect 208860 620 208912 672
rect 241060 620 241112 672
rect 111984 552 112036 604
rect 138664 552 138716 604
rect 172520 552 172572 604
rect 217324 552 217376 604
rect 223028 552 223080 604
rect 223120 552 223172 604
rect 248972 552 249024 604
rect 152464 484 152516 536
rect 158352 484 158404 536
rect 5448 416 5500 468
rect 40132 416 40184 468
rect 72424 416 72476 468
rect 99748 416 99800 468
rect 100392 416 100444 468
rect 106372 416 106424 468
rect 148784 416 148836 468
rect 160468 416 160520 468
rect 2872 348 2924 400
rect 37740 348 37792 400
rect 151544 348 151596 400
rect 152556 348 152608 400
rect 154304 348 154356 400
rect 187148 484 187200 536
rect 211068 484 211120 536
rect 243820 484 243872 536
rect 211344 416 211396 468
rect 216588 416 216640 468
rect 227996 416 228048 468
rect 217876 348 217928 400
rect 219624 348 219676 400
rect 220728 348 220780 400
rect 224132 348 224184 400
rect 256516 416 256568 468
rect 235724 348 235776 400
rect 268936 348 268988 400
rect 9404 280 9456 332
rect 41052 280 41104 332
rect 216220 280 216272 332
rect 223120 280 223172 332
rect 227904 280 227956 332
rect 251824 280 251876 332
rect 222844 212 222896 264
rect 229744 212 229796 264
<< metal2 >>
rect 97632 10872 97684 10878
rect 97632 10814 97684 10820
rect 98460 10872 98512 10878
rect 98460 10814 98512 10820
rect 152372 10872 152424 10878
rect 152372 10814 152424 10820
rect 163964 10872 164016 10878
rect 163964 10814 164016 10820
rect 214288 10872 214340 10878
rect 227444 10872 227496 10878
rect 214288 10814 214340 10820
rect 227442 10840 227444 10849
rect 229100 10872 229152 10878
rect 227496 10840 227498 10849
rect 90824 10804 90876 10810
rect 90824 10746 90876 10752
rect 95056 10804 95108 10810
rect 95056 10746 95108 10752
rect 96988 10804 97040 10810
rect 96988 10746 97040 10752
rect 28448 10736 28500 10742
rect 28448 10678 28500 10684
rect 33784 10736 33836 10742
rect 33784 10678 33836 10684
rect 65984 10736 66036 10742
rect 65984 10678 66036 10684
rect 23940 10600 23992 10606
rect 9678 10568 9734 10577
rect 9678 10503 9734 10512
rect 20718 10568 20774 10577
rect 23940 10542 23992 10548
rect 20718 10503 20774 10512
rect 23756 10532 23808 10538
rect 1674 10160 1730 10169
rect 1674 10095 1730 10104
rect 2410 10160 2466 10169
rect 2410 10095 2466 10104
rect 3238 10160 3294 10169
rect 3238 10095 3294 10104
rect 4342 10160 4398 10169
rect 4342 10095 4398 10104
rect 5078 10160 5134 10169
rect 5078 10095 5134 10104
rect 5814 10160 5870 10169
rect 5814 10095 5870 10104
rect 6826 10160 6882 10169
rect 6826 10095 6882 10104
rect 7562 10160 7618 10169
rect 8390 10160 8446 10169
rect 7562 10095 7618 10104
rect 7656 10124 7708 10130
rect 1688 9654 1716 10095
rect 2424 9654 2452 10095
rect 3146 9888 3202 9897
rect 3146 9823 3202 9832
rect 1676 9648 1728 9654
rect 1676 9590 1728 9596
rect 2412 9648 2464 9654
rect 2412 9590 2464 9596
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 1398 9208 1454 9217
rect 2424 9178 2452 9318
rect 1398 9143 1400 9152
rect 1452 9143 1454 9152
rect 2412 9172 2464 9178
rect 1400 9114 1452 9120
rect 2412 9114 2464 9120
rect 2516 9042 2544 9318
rect 2504 9036 2556 9042
rect 2504 8978 2556 8984
rect 3160 8974 3188 9823
rect 3252 9654 3280 10095
rect 4356 9654 4384 10095
rect 5092 9654 5120 10095
rect 5828 9654 5856 10095
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 5920 9722 5948 9998
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 6840 9654 6868 10095
rect 7576 9654 7604 10095
rect 8390 10095 8446 10104
rect 7656 10066 7708 10072
rect 7668 9722 7696 10066
rect 8206 9888 8262 9897
rect 8206 9823 8262 9832
rect 7656 9716 7708 9722
rect 7656 9658 7708 9664
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 7564 9648 7616 9654
rect 7564 9590 7616 9596
rect 3424 9444 3476 9450
rect 3424 9386 3476 9392
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3332 8900 3384 8906
rect 3332 8842 3384 8848
rect 3344 3738 3372 8842
rect 3436 8294 3464 9386
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6932 8634 6960 9318
rect 8220 8974 8248 9823
rect 8404 9654 8432 10095
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8496 9722 8524 9862
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 9692 9586 9720 10503
rect 20732 10402 20760 10503
rect 23756 10474 23808 10480
rect 20720 10396 20772 10402
rect 20720 10338 20772 10344
rect 22836 10328 22888 10334
rect 22836 10270 22888 10276
rect 11978 10160 12034 10169
rect 11978 10095 12034 10104
rect 12714 10160 12770 10169
rect 12714 10095 12770 10104
rect 13726 10160 13782 10169
rect 13726 10095 13782 10104
rect 14646 10160 14702 10169
rect 14646 10095 14702 10104
rect 15382 10160 15438 10169
rect 15382 10095 15438 10104
rect 16118 10160 16174 10169
rect 16118 10095 16174 10104
rect 17130 10160 17186 10169
rect 17130 10095 17186 10104
rect 17866 10160 17922 10169
rect 17866 10095 17922 10104
rect 18602 10160 18658 10169
rect 18602 10095 18658 10104
rect 22374 10160 22430 10169
rect 22374 10095 22430 10104
rect 10506 9888 10562 9897
rect 10506 9823 10562 9832
rect 11242 9888 11298 9897
rect 11242 9823 11298 9832
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8484 8900 8536 8906
rect 8484 8842 8536 8848
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 8496 4486 8524 8842
rect 9968 6322 9996 9454
rect 10520 8974 10548 9823
rect 11256 8974 11284 9823
rect 11992 9654 12020 10095
rect 12728 9654 12756 10095
rect 13450 9888 13506 9897
rect 13450 9823 13506 9832
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 12716 9648 12768 9654
rect 12716 9590 12768 9596
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12820 9110 12848 9318
rect 12808 9104 12860 9110
rect 12808 9046 12860 9052
rect 13464 8974 13492 9823
rect 13740 9654 13768 10095
rect 14660 9654 14688 10095
rect 15396 9654 15424 10095
rect 16132 9654 16160 10095
rect 17144 9654 17172 10095
rect 17316 9988 17368 9994
rect 17316 9930 17368 9936
rect 17328 9654 17356 9930
rect 17880 9654 17908 10095
rect 18616 9654 18644 10095
rect 21454 9888 21510 9897
rect 21454 9823 21510 9832
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 14648 9648 14700 9654
rect 14648 9590 14700 9596
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 16120 9648 16172 9654
rect 16120 9590 16172 9596
rect 17132 9648 17184 9654
rect 17132 9590 17184 9596
rect 17316 9648 17368 9654
rect 17316 9590 17368 9596
rect 17868 9648 17920 9654
rect 17868 9590 17920 9596
rect 18604 9648 18656 9654
rect 18604 9590 18656 9596
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 11348 5642 11376 8774
rect 13556 8362 13584 8774
rect 13544 8356 13596 8362
rect 13544 8298 13596 8304
rect 13740 6390 13768 9386
rect 14752 7954 14780 9454
rect 15568 9444 15620 9450
rect 15568 9386 15620 9392
rect 20352 9444 20404 9450
rect 20352 9386 20404 9392
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 13728 6384 13780 6390
rect 13728 6326 13780 6332
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 15304 5370 15332 9318
rect 15580 6458 15608 9386
rect 17224 8900 17276 8906
rect 17224 8842 17276 8848
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 17236 6186 17264 8842
rect 20364 7478 20392 9386
rect 21468 8906 21496 9823
rect 22388 9654 22416 10095
rect 22376 9648 22428 9654
rect 22376 9590 22428 9596
rect 22848 9042 22876 10270
rect 23664 10056 23716 10062
rect 23664 9998 23716 10004
rect 23572 9580 23624 9586
rect 23572 9522 23624 9528
rect 23388 9376 23440 9382
rect 23388 9318 23440 9324
rect 23112 9172 23164 9178
rect 23112 9114 23164 9120
rect 22744 9036 22796 9042
rect 22744 8978 22796 8984
rect 22836 9036 22888 9042
rect 22836 8978 22888 8984
rect 21456 8900 21508 8906
rect 21456 8842 21508 8848
rect 20352 7472 20404 7478
rect 20352 7414 20404 7420
rect 19246 6896 19302 6905
rect 19246 6831 19302 6840
rect 19982 6896 20038 6905
rect 19982 6831 20038 6840
rect 19260 6662 19288 6831
rect 19996 6798 20024 6831
rect 19984 6792 20036 6798
rect 19984 6734 20036 6740
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 17224 6180 17276 6186
rect 17224 6122 17276 6128
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 20718 5128 20774 5137
rect 20718 5063 20774 5072
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 8484 4480 8536 4486
rect 8484 4422 8536 4428
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 4804 2576 4856 2582
rect 4804 2518 4856 2524
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 846 1456 902 1465
rect 846 1391 848 1400
rect 900 1391 902 1400
rect 848 1362 900 1368
rect 1596 1329 1624 2382
rect 2596 2372 2648 2378
rect 2596 2314 2648 2320
rect 2608 1970 2636 2314
rect 4816 1970 4844 2518
rect 9232 2038 9260 3946
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 9220 2032 9272 2038
rect 9220 1974 9272 1980
rect 2596 1964 2648 1970
rect 2596 1906 2648 1912
rect 4804 1964 4856 1970
rect 4804 1906 4856 1912
rect 6828 1964 6880 1970
rect 6828 1906 6880 1912
rect 7564 1964 7616 1970
rect 7564 1906 7616 1912
rect 9036 1964 9088 1970
rect 9036 1906 9088 1912
rect 2320 1896 2372 1902
rect 2320 1838 2372 1844
rect 4528 1896 4580 1902
rect 4528 1838 4580 1844
rect 1582 1320 1638 1329
rect 1582 1255 1638 1264
rect 2332 1057 2360 1838
rect 2872 1352 2924 1358
rect 2872 1294 2924 1300
rect 2318 1048 2374 1057
rect 2318 983 2374 992
rect 2884 406 2912 1294
rect 2964 1284 3016 1290
rect 2964 1226 3016 1232
rect 4068 1284 4120 1290
rect 4068 1226 4120 1232
rect 2976 785 3004 1226
rect 2962 776 3018 785
rect 2962 711 3018 720
rect 4080 649 4108 1226
rect 4160 1216 4212 1222
rect 4160 1158 4212 1164
rect 4172 814 4200 1158
rect 4540 1057 4568 1838
rect 5172 1352 5224 1358
rect 5172 1294 5224 1300
rect 5448 1352 5500 1358
rect 5448 1294 5500 1300
rect 6552 1352 6604 1358
rect 6552 1294 6604 1300
rect 4526 1048 4582 1057
rect 4526 983 4582 992
rect 4160 808 4212 814
rect 5184 785 5212 1294
rect 4160 750 4212 756
rect 5170 776 5226 785
rect 5170 711 5226 720
rect 4066 640 4122 649
rect 4066 575 4122 584
rect 5460 474 5488 1294
rect 6564 785 6592 1294
rect 6840 1057 6868 1906
rect 6826 1048 6882 1057
rect 6826 983 6882 992
rect 7576 785 7604 1906
rect 8208 1284 8260 1290
rect 8208 1226 8260 1232
rect 6550 776 6606 785
rect 6550 711 6606 720
rect 7562 776 7618 785
rect 7562 711 7618 720
rect 8220 649 8248 1226
rect 8392 1216 8444 1222
rect 8392 1158 8444 1164
rect 8206 640 8262 649
rect 8404 610 8432 1158
rect 9048 785 9076 1906
rect 11164 1358 11192 3402
rect 12176 1358 12204 4762
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14384 1970 14412 4014
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 14372 1964 14424 1970
rect 14372 1906 14424 1912
rect 14096 1896 14148 1902
rect 14096 1838 14148 1844
rect 9404 1352 9456 1358
rect 9404 1294 9456 1300
rect 9588 1352 9640 1358
rect 9588 1294 9640 1300
rect 11152 1352 11204 1358
rect 11152 1294 11204 1300
rect 12164 1352 12216 1358
rect 12164 1294 12216 1300
rect 9034 776 9090 785
rect 9034 711 9090 720
rect 8206 575 8262 584
rect 8392 604 8444 610
rect 8392 546 8444 552
rect 5448 468 5500 474
rect 5448 410 5500 416
rect 2872 400 2924 406
rect 2872 342 2924 348
rect 9416 338 9444 1294
rect 9600 649 9628 1294
rect 9680 1284 9732 1290
rect 9680 1226 9732 1232
rect 10232 1284 10284 1290
rect 10232 1226 10284 1232
rect 10416 1284 10468 1290
rect 10416 1226 10468 1232
rect 10968 1284 11020 1290
rect 10968 1226 11020 1232
rect 11980 1284 12032 1290
rect 11980 1226 12032 1232
rect 12716 1284 12768 1290
rect 12716 1226 12768 1232
rect 13452 1284 13504 1290
rect 13452 1226 13504 1232
rect 9692 678 9720 1226
rect 9680 672 9732 678
rect 9586 640 9642 649
rect 10244 649 10272 1226
rect 10428 1193 10456 1226
rect 10414 1184 10470 1193
rect 10414 1119 10470 1128
rect 10980 649 11008 1226
rect 11992 649 12020 1226
rect 12728 649 12756 1226
rect 12808 1216 12860 1222
rect 12808 1158 12860 1164
rect 12820 746 12848 1158
rect 12808 740 12860 746
rect 12808 682 12860 688
rect 13464 649 13492 1226
rect 13544 1216 13596 1222
rect 13544 1158 13596 1164
rect 13556 1018 13584 1158
rect 14108 1057 14136 1838
rect 15120 1358 15148 3538
rect 17144 2038 17172 4966
rect 19338 4448 19394 4457
rect 19338 4383 19394 4392
rect 19352 3602 19380 4383
rect 19340 3596 19392 3602
rect 19340 3538 19392 3544
rect 20732 3466 20760 5063
rect 22756 3466 22784 8978
rect 23124 8566 23152 9114
rect 23296 8628 23348 8634
rect 23296 8570 23348 8576
rect 23112 8560 23164 8566
rect 23112 8502 23164 8508
rect 23204 8356 23256 8362
rect 23204 8298 23256 8304
rect 23216 8022 23244 8298
rect 23204 8016 23256 8022
rect 23204 7958 23256 7964
rect 23308 4282 23336 8570
rect 23400 7274 23428 9318
rect 23478 8664 23534 8673
rect 23478 8599 23480 8608
rect 23532 8599 23534 8608
rect 23480 8570 23532 8576
rect 23388 7268 23440 7274
rect 23388 7210 23440 7216
rect 23480 7200 23532 7206
rect 23480 7142 23532 7148
rect 23492 6905 23520 7142
rect 23478 6896 23534 6905
rect 23478 6831 23534 6840
rect 23584 6066 23612 9522
rect 23676 6254 23704 9998
rect 23768 9586 23796 10474
rect 23756 9580 23808 9586
rect 23756 9522 23808 9528
rect 23848 9580 23900 9586
rect 23848 9522 23900 9528
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23768 8498 23796 9318
rect 23860 8974 23888 9522
rect 23952 9382 23980 10542
rect 25780 10464 25832 10470
rect 25780 10406 25832 10412
rect 24952 10328 25004 10334
rect 24952 10270 25004 10276
rect 24400 9444 24452 9450
rect 24400 9386 24452 9392
rect 23940 9376 23992 9382
rect 23940 9318 23992 9324
rect 23940 9036 23992 9042
rect 23940 8978 23992 8984
rect 23848 8968 23900 8974
rect 23848 8910 23900 8916
rect 23756 8492 23808 8498
rect 23756 8434 23808 8440
rect 23664 6248 23716 6254
rect 23664 6190 23716 6196
rect 23584 6038 23704 6066
rect 23296 4276 23348 4282
rect 23296 4218 23348 4224
rect 23572 4140 23624 4146
rect 23572 4082 23624 4088
rect 20720 3460 20772 3466
rect 20720 3402 20772 3408
rect 22744 3460 22796 3466
rect 22744 3402 22796 3408
rect 19248 2984 19300 2990
rect 19246 2952 19248 2961
rect 19300 2952 19302 2961
rect 19246 2887 19302 2896
rect 22926 2952 22982 2961
rect 22926 2887 22928 2896
rect 22980 2887 22982 2896
rect 22928 2858 22980 2864
rect 19984 2848 20036 2854
rect 19982 2816 19984 2825
rect 20036 2816 20038 2825
rect 19982 2751 20038 2760
rect 23386 2816 23442 2825
rect 23442 2774 23520 2802
rect 23386 2751 23442 2760
rect 23492 2650 23520 2774
rect 23480 2644 23532 2650
rect 23480 2586 23532 2592
rect 23584 2582 23612 4082
rect 23572 2576 23624 2582
rect 23572 2518 23624 2524
rect 23676 2394 23704 6038
rect 23768 5794 23796 8434
rect 23952 5930 23980 8978
rect 24124 8968 24176 8974
rect 24124 8910 24176 8916
rect 24032 8832 24084 8838
rect 24030 8800 24032 8809
rect 24084 8800 24086 8809
rect 24030 8735 24086 8744
rect 24136 8514 24164 8910
rect 24044 8498 24164 8514
rect 24032 8492 24164 8498
rect 24084 8486 24164 8492
rect 24032 8434 24084 8440
rect 24216 8424 24268 8430
rect 24216 8366 24268 8372
rect 24228 6798 24256 8366
rect 24216 6792 24268 6798
rect 24216 6734 24268 6740
rect 24412 6730 24440 9386
rect 24492 9376 24544 9382
rect 24492 9318 24544 9324
rect 24504 7410 24532 9318
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 24872 8430 24900 8978
rect 24860 8424 24912 8430
rect 24860 8366 24912 8372
rect 24492 7404 24544 7410
rect 24492 7346 24544 7352
rect 24766 6896 24822 6905
rect 24766 6831 24822 6840
rect 24400 6724 24452 6730
rect 24400 6666 24452 6672
rect 24780 6662 24808 6831
rect 24768 6656 24820 6662
rect 24768 6598 24820 6604
rect 23952 5902 24072 5930
rect 23768 5766 23980 5794
rect 23756 3392 23808 3398
rect 23756 3334 23808 3340
rect 23768 2446 23796 3334
rect 23848 3052 23900 3058
rect 23848 2994 23900 3000
rect 23584 2366 23704 2394
rect 23756 2440 23808 2446
rect 23756 2382 23808 2388
rect 17132 2032 17184 2038
rect 15842 2000 15898 2009
rect 15660 1964 15712 1970
rect 17132 1974 17184 1980
rect 23584 1970 23612 2366
rect 23860 2106 23888 2994
rect 23848 2100 23900 2106
rect 23848 2042 23900 2048
rect 23952 1970 23980 5766
rect 15842 1935 15844 1944
rect 15660 1906 15712 1912
rect 15896 1935 15898 1944
rect 16580 1964 16632 1970
rect 15844 1906 15896 1912
rect 16580 1906 16632 1912
rect 23572 1964 23624 1970
rect 23572 1906 23624 1912
rect 23940 1964 23992 1970
rect 23940 1906 23992 1912
rect 14832 1352 14884 1358
rect 14832 1294 14884 1300
rect 15108 1352 15160 1358
rect 15108 1294 15160 1300
rect 14094 1048 14150 1057
rect 13544 1012 13596 1018
rect 14094 983 14150 992
rect 13544 954 13596 960
rect 14844 785 14872 1294
rect 15672 785 15700 1906
rect 16592 1465 16620 1906
rect 22192 1828 22244 1834
rect 22192 1770 22244 1776
rect 22204 1737 22232 1770
rect 23664 1760 23716 1766
rect 22190 1728 22246 1737
rect 23664 1702 23716 1708
rect 23756 1760 23808 1766
rect 23756 1702 23808 1708
rect 22190 1663 22246 1672
rect 22100 1556 22152 1562
rect 22100 1498 22152 1504
rect 22112 1465 22140 1498
rect 23676 1494 23704 1702
rect 23664 1488 23716 1494
rect 16578 1456 16634 1465
rect 16578 1391 16634 1400
rect 22098 1456 22154 1465
rect 23664 1430 23716 1436
rect 22098 1391 22154 1400
rect 23768 1358 23796 1702
rect 24044 1426 24072 5902
rect 24492 3936 24544 3942
rect 24492 3878 24544 3884
rect 24504 3369 24532 3878
rect 24964 3602 24992 10270
rect 25136 9580 25188 9586
rect 25136 9522 25188 9528
rect 25148 9178 25176 9522
rect 25136 9172 25188 9178
rect 25136 9114 25188 9120
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 25056 8498 25084 8910
rect 25136 8900 25188 8906
rect 25136 8842 25188 8848
rect 25044 8492 25096 8498
rect 25044 8434 25096 8440
rect 25056 7886 25084 8434
rect 25044 7880 25096 7886
rect 25044 7822 25096 7828
rect 25056 7410 25084 7822
rect 25148 7546 25176 8842
rect 25686 8800 25742 8809
rect 25686 8735 25742 8744
rect 25700 8566 25728 8735
rect 25688 8560 25740 8566
rect 25688 8502 25740 8508
rect 25792 8430 25820 10406
rect 25964 10396 26016 10402
rect 25964 10338 26016 10344
rect 25870 9616 25926 9625
rect 25870 9551 25926 9560
rect 25884 9450 25912 9551
rect 25872 9444 25924 9450
rect 25872 9386 25924 9392
rect 25976 8566 26004 10338
rect 26056 10260 26108 10266
rect 26056 10202 26108 10208
rect 26068 9518 26096 10202
rect 27620 10192 27672 10198
rect 27620 10134 27672 10140
rect 26700 10124 26752 10130
rect 26700 10066 26752 10072
rect 26712 9908 26740 10066
rect 27068 9988 27120 9994
rect 27068 9930 27120 9936
rect 26976 9920 27028 9926
rect 26712 9880 26976 9908
rect 26976 9862 27028 9868
rect 26056 9512 26108 9518
rect 26056 9454 26108 9460
rect 25964 8560 26016 8566
rect 25964 8502 26016 8508
rect 25504 8424 25556 8430
rect 25504 8366 25556 8372
rect 25780 8424 25832 8430
rect 26068 8378 26096 9454
rect 26884 9376 26936 9382
rect 26884 9318 26936 9324
rect 26240 9036 26292 9042
rect 26240 8978 26292 8984
rect 26148 8832 26200 8838
rect 26148 8774 26200 8780
rect 25780 8366 25832 8372
rect 25228 8356 25280 8362
rect 25228 8298 25280 8304
rect 25240 8090 25268 8298
rect 25228 8084 25280 8090
rect 25228 8026 25280 8032
rect 25136 7540 25188 7546
rect 25136 7482 25188 7488
rect 25044 7404 25096 7410
rect 25044 7346 25096 7352
rect 25228 7336 25280 7342
rect 25228 7278 25280 7284
rect 24952 3596 25004 3602
rect 24952 3538 25004 3544
rect 25044 3528 25096 3534
rect 25044 3470 25096 3476
rect 24490 3360 24546 3369
rect 24490 3295 24546 3304
rect 24860 2984 24912 2990
rect 24860 2926 24912 2932
rect 24872 1766 24900 2926
rect 25056 2446 25084 3470
rect 25240 3097 25268 7278
rect 25412 3528 25464 3534
rect 25412 3470 25464 3476
rect 25226 3088 25282 3097
rect 25424 3058 25452 3470
rect 25226 3023 25282 3032
rect 25412 3052 25464 3058
rect 25240 2990 25268 3023
rect 25412 2994 25464 3000
rect 25228 2984 25280 2990
rect 25228 2926 25280 2932
rect 25136 2576 25188 2582
rect 25136 2518 25188 2524
rect 24952 2440 25004 2446
rect 24952 2382 25004 2388
rect 25044 2440 25096 2446
rect 25044 2382 25096 2388
rect 24964 1970 24992 2382
rect 24952 1964 25004 1970
rect 24952 1906 25004 1912
rect 25056 1902 25084 2382
rect 25148 2038 25176 2518
rect 25516 2446 25544 8366
rect 25884 8350 26096 8378
rect 25688 7744 25740 7750
rect 25688 7686 25740 7692
rect 25596 2848 25648 2854
rect 25596 2790 25648 2796
rect 25504 2440 25556 2446
rect 25504 2382 25556 2388
rect 25608 2038 25636 2790
rect 25700 2446 25728 7686
rect 25780 4140 25832 4146
rect 25780 4082 25832 4088
rect 25792 2650 25820 4082
rect 25780 2644 25832 2650
rect 25780 2586 25832 2592
rect 25688 2440 25740 2446
rect 25688 2382 25740 2388
rect 25136 2032 25188 2038
rect 25136 1974 25188 1980
rect 25596 2032 25648 2038
rect 25596 1974 25648 1980
rect 25700 1970 25728 2382
rect 25688 1964 25740 1970
rect 25688 1906 25740 1912
rect 25044 1896 25096 1902
rect 25044 1838 25096 1844
rect 25136 1896 25188 1902
rect 25136 1838 25188 1844
rect 24860 1760 24912 1766
rect 24860 1702 24912 1708
rect 25056 1426 25084 1838
rect 24032 1420 24084 1426
rect 24032 1362 24084 1368
rect 24952 1420 25004 1426
rect 24952 1362 25004 1368
rect 25044 1420 25096 1426
rect 25044 1362 25096 1368
rect 23756 1352 23808 1358
rect 23756 1294 23808 1300
rect 24964 1306 24992 1362
rect 25148 1306 25176 1838
rect 25884 1426 25912 8350
rect 26056 7336 26108 7342
rect 26056 7278 26108 7284
rect 25964 3392 26016 3398
rect 25964 3334 26016 3340
rect 25872 1420 25924 1426
rect 25872 1362 25924 1368
rect 25976 1329 26004 3334
rect 26068 2990 26096 7278
rect 26160 6866 26188 8774
rect 26252 8566 26280 8978
rect 26424 8900 26476 8906
rect 26424 8842 26476 8848
rect 26240 8560 26292 8566
rect 26240 8502 26292 8508
rect 26252 7818 26280 8502
rect 26240 7812 26292 7818
rect 26240 7754 26292 7760
rect 26252 7410 26280 7754
rect 26436 7546 26464 8842
rect 26896 8838 26924 9318
rect 27080 8906 27108 9930
rect 27528 9580 27580 9586
rect 27528 9522 27580 9528
rect 27540 8974 27568 9522
rect 27528 8968 27580 8974
rect 27528 8910 27580 8916
rect 27068 8900 27120 8906
rect 27068 8842 27120 8848
rect 26884 8832 26936 8838
rect 26884 8774 26936 8780
rect 26698 8392 26754 8401
rect 26698 8327 26754 8336
rect 26608 7880 26660 7886
rect 26608 7822 26660 7828
rect 26516 7744 26568 7750
rect 26516 7686 26568 7692
rect 26424 7540 26476 7546
rect 26424 7482 26476 7488
rect 26240 7404 26292 7410
rect 26240 7346 26292 7352
rect 26240 7200 26292 7206
rect 26240 7142 26292 7148
rect 26252 6905 26280 7142
rect 26238 6896 26294 6905
rect 26148 6860 26200 6866
rect 26238 6831 26294 6840
rect 26148 6802 26200 6808
rect 26528 6798 26556 7686
rect 26620 7546 26648 7822
rect 26608 7540 26660 7546
rect 26608 7482 26660 7488
rect 26516 6792 26568 6798
rect 26516 6734 26568 6740
rect 26620 6474 26648 7482
rect 26712 6662 26740 8327
rect 26884 8288 26936 8294
rect 26884 8230 26936 8236
rect 26976 8288 27028 8294
rect 26976 8230 27028 8236
rect 26792 7812 26844 7818
rect 26792 7754 26844 7760
rect 26804 7478 26832 7754
rect 26792 7472 26844 7478
rect 26792 7414 26844 7420
rect 26700 6656 26752 6662
rect 26700 6598 26752 6604
rect 26620 6446 26832 6474
rect 26240 3528 26292 3534
rect 26240 3470 26292 3476
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 26148 3052 26200 3058
rect 26148 2994 26200 3000
rect 26056 2984 26108 2990
rect 26056 2926 26108 2932
rect 26160 2446 26188 2994
rect 26252 2650 26280 3470
rect 26332 3120 26384 3126
rect 26332 3062 26384 3068
rect 26240 2644 26292 2650
rect 26240 2586 26292 2592
rect 26148 2440 26200 2446
rect 26148 2382 26200 2388
rect 26344 2106 26372 3062
rect 26424 2848 26476 2854
rect 26424 2790 26476 2796
rect 26332 2100 26384 2106
rect 26332 2042 26384 2048
rect 26436 2038 26464 2790
rect 26528 2650 26556 3470
rect 26700 3392 26752 3398
rect 26700 3334 26752 3340
rect 26516 2644 26568 2650
rect 26516 2586 26568 2592
rect 26424 2032 26476 2038
rect 26424 1974 26476 1980
rect 26712 1329 26740 3334
rect 26804 2446 26832 6446
rect 26896 5302 26924 8230
rect 26988 6934 27016 8230
rect 26976 6928 27028 6934
rect 26976 6870 27028 6876
rect 26884 5296 26936 5302
rect 26884 5238 26936 5244
rect 27080 3126 27108 8842
rect 27540 7886 27568 8910
rect 27632 8294 27660 10134
rect 27712 9512 27764 9518
rect 27712 9454 27764 9460
rect 27724 9178 27752 9454
rect 28172 9376 28224 9382
rect 28172 9318 28224 9324
rect 27712 9172 27764 9178
rect 27712 9114 27764 9120
rect 27620 8288 27672 8294
rect 27620 8230 27672 8236
rect 27344 7880 27396 7886
rect 27344 7822 27396 7828
rect 27528 7880 27580 7886
rect 27528 7822 27580 7828
rect 27252 3188 27304 3194
rect 27252 3130 27304 3136
rect 27068 3120 27120 3126
rect 27068 3062 27120 3068
rect 26792 2440 26844 2446
rect 26792 2382 26844 2388
rect 27264 2310 27292 3130
rect 27356 2446 27384 7822
rect 27724 7290 27752 9114
rect 28184 7886 28212 9318
rect 28460 8498 28488 10678
rect 29920 10668 29972 10674
rect 29920 10610 29972 10616
rect 29092 10260 29144 10266
rect 29092 10202 29144 10208
rect 29000 9988 29052 9994
rect 29000 9930 29052 9936
rect 29012 9654 29040 9930
rect 28908 9648 28960 9654
rect 28908 9590 28960 9596
rect 29000 9648 29052 9654
rect 29000 9590 29052 9596
rect 28724 9580 28776 9586
rect 28724 9522 28776 9528
rect 28736 8634 28764 9522
rect 28814 9480 28870 9489
rect 28814 9415 28816 9424
rect 28868 9415 28870 9424
rect 28816 9386 28868 9392
rect 28724 8628 28776 8634
rect 28724 8570 28776 8576
rect 28448 8492 28500 8498
rect 28448 8434 28500 8440
rect 28354 8392 28410 8401
rect 28354 8327 28410 8336
rect 28368 8090 28396 8327
rect 28356 8084 28408 8090
rect 28356 8026 28408 8032
rect 28172 7880 28224 7886
rect 27894 7848 27950 7857
rect 28172 7822 28224 7828
rect 27894 7783 27950 7792
rect 27908 7750 27936 7783
rect 27804 7744 27856 7750
rect 27804 7686 27856 7692
rect 27896 7744 27948 7750
rect 27896 7686 27948 7692
rect 27816 7410 27844 7686
rect 27804 7404 27856 7410
rect 27804 7346 27856 7352
rect 27724 7262 27844 7290
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 27436 3392 27488 3398
rect 27436 3334 27488 3340
rect 27344 2440 27396 2446
rect 27344 2382 27396 2388
rect 27252 2304 27304 2310
rect 27252 2246 27304 2252
rect 27448 1329 27476 3334
rect 27540 1358 27568 3470
rect 27620 3460 27672 3466
rect 27620 3402 27672 3408
rect 27632 3126 27660 3402
rect 27620 3120 27672 3126
rect 27620 3062 27672 3068
rect 27712 2848 27764 2854
rect 27712 2790 27764 2796
rect 27724 2038 27752 2790
rect 27712 2032 27764 2038
rect 27712 1974 27764 1980
rect 27816 1426 27844 7262
rect 27896 3052 27948 3058
rect 27896 2994 27948 3000
rect 27988 3052 28040 3058
rect 27988 2994 28040 3000
rect 27908 2446 27936 2994
rect 28000 2650 28028 2994
rect 28080 2916 28132 2922
rect 28080 2858 28132 2864
rect 28092 2825 28120 2858
rect 28078 2816 28134 2825
rect 28078 2751 28134 2760
rect 27988 2644 28040 2650
rect 27988 2586 28040 2592
rect 27896 2440 27948 2446
rect 27896 2382 27948 2388
rect 27908 2310 27936 2382
rect 27896 2304 27948 2310
rect 27896 2246 27948 2252
rect 27908 2038 27936 2246
rect 27896 2032 27948 2038
rect 27896 1974 27948 1980
rect 28460 1970 28488 8434
rect 28540 8016 28592 8022
rect 28540 7958 28592 7964
rect 28552 7274 28580 7958
rect 28920 7886 28948 9590
rect 29104 9518 29132 10202
rect 29736 9580 29788 9586
rect 29736 9522 29788 9528
rect 29000 9512 29052 9518
rect 29000 9454 29052 9460
rect 29092 9512 29144 9518
rect 29092 9454 29144 9460
rect 29012 8974 29040 9454
rect 29000 8968 29052 8974
rect 29000 8910 29052 8916
rect 29012 8498 29040 8910
rect 29552 8900 29604 8906
rect 29552 8842 29604 8848
rect 29092 8832 29144 8838
rect 29092 8774 29144 8780
rect 29460 8832 29512 8838
rect 29460 8774 29512 8780
rect 29000 8492 29052 8498
rect 29000 8434 29052 8440
rect 29104 7886 29132 8774
rect 29472 8498 29500 8774
rect 29460 8492 29512 8498
rect 29460 8434 29512 8440
rect 28908 7880 28960 7886
rect 28908 7822 28960 7828
rect 29092 7880 29144 7886
rect 29092 7822 29144 7828
rect 28540 7268 28592 7274
rect 28540 7210 28592 7216
rect 28540 2440 28592 2446
rect 28540 2382 28592 2388
rect 28448 1964 28500 1970
rect 28448 1906 28500 1912
rect 28552 1562 28580 2382
rect 28724 2304 28776 2310
rect 28724 2246 28776 2252
rect 28540 1556 28592 1562
rect 28540 1498 28592 1504
rect 27804 1420 27856 1426
rect 27804 1362 27856 1368
rect 27528 1352 27580 1358
rect 17132 1284 17184 1290
rect 17132 1226 17184 1232
rect 17868 1284 17920 1290
rect 17868 1226 17920 1232
rect 18604 1284 18656 1290
rect 24964 1278 25176 1306
rect 25962 1320 26018 1329
rect 25962 1255 26018 1264
rect 26698 1320 26754 1329
rect 26698 1255 26754 1264
rect 27434 1320 27490 1329
rect 27528 1294 27580 1300
rect 27434 1255 27490 1264
rect 18604 1226 18656 1232
rect 14830 776 14886 785
rect 14830 711 14886 720
rect 15658 776 15714 785
rect 15658 711 15714 720
rect 17144 649 17172 1226
rect 17224 1216 17276 1222
rect 17224 1158 17276 1164
rect 17236 882 17264 1158
rect 17224 876 17276 882
rect 17224 818 17276 824
rect 17880 649 17908 1226
rect 17960 1216 18012 1222
rect 17960 1158 18012 1164
rect 9680 614 9732 620
rect 10230 640 10286 649
rect 9586 575 9642 584
rect 10230 575 10286 584
rect 10966 640 11022 649
rect 10966 575 11022 584
rect 11978 640 12034 649
rect 11978 575 12034 584
rect 12714 640 12770 649
rect 12714 575 12770 584
rect 13450 640 13506 649
rect 13450 575 13506 584
rect 17130 640 17186 649
rect 17130 575 17186 584
rect 17866 640 17922 649
rect 17866 575 17922 584
rect 17972 542 18000 1158
rect 18616 649 18644 1226
rect 18696 1216 18748 1222
rect 18696 1158 18748 1164
rect 23940 1216 23992 1222
rect 23940 1158 23992 1164
rect 18708 950 18736 1158
rect 18696 944 18748 950
rect 18696 886 18748 892
rect 23952 649 23980 1158
rect 18602 640 18658 649
rect 18602 575 18658 584
rect 23938 640 23994 649
rect 23938 575 23994 584
rect 17960 536 18012 542
rect 28736 513 28764 2246
rect 29564 1970 29592 8842
rect 29642 8664 29698 8673
rect 29642 8599 29644 8608
rect 29696 8599 29698 8608
rect 29644 8570 29696 8576
rect 29748 8566 29776 9522
rect 29932 8906 29960 10610
rect 30012 10532 30064 10538
rect 30012 10474 30064 10480
rect 30024 9382 30052 10474
rect 33796 10402 33824 10678
rect 63224 10668 63276 10674
rect 63224 10610 63276 10616
rect 60372 10600 60424 10606
rect 60372 10542 60424 10548
rect 60096 10532 60148 10538
rect 60096 10474 60148 10480
rect 57152 10464 57204 10470
rect 54666 10432 54722 10441
rect 33784 10396 33836 10402
rect 57152 10406 57204 10412
rect 54666 10367 54722 10376
rect 33784 10338 33836 10344
rect 31758 10296 31814 10305
rect 31758 10231 31814 10240
rect 35162 10296 35218 10305
rect 35162 10231 35218 10240
rect 35622 10296 35678 10305
rect 35622 10231 35678 10240
rect 36266 10296 36322 10305
rect 36266 10231 36322 10240
rect 36910 10296 36966 10305
rect 36910 10231 36966 10240
rect 38106 10296 38162 10305
rect 38106 10231 38162 10240
rect 38842 10296 38898 10305
rect 38842 10231 38898 10240
rect 39486 10296 39542 10305
rect 39486 10231 39542 10240
rect 40314 10296 40370 10305
rect 40314 10231 40370 10240
rect 40774 10296 40830 10305
rect 40774 10231 40830 10240
rect 41418 10296 41474 10305
rect 41418 10231 41474 10240
rect 42062 10296 42118 10305
rect 42062 10231 42118 10240
rect 43258 10296 43314 10305
rect 43258 10231 43314 10240
rect 43994 10296 44050 10305
rect 43994 10231 44050 10240
rect 44638 10296 44694 10305
rect 44638 10231 44694 10240
rect 45466 10296 45522 10305
rect 45466 10231 45522 10240
rect 45926 10296 45982 10305
rect 45926 10231 45982 10240
rect 46570 10296 46626 10305
rect 46570 10231 46626 10240
rect 47214 10296 47270 10305
rect 47214 10231 47270 10240
rect 48226 10296 48282 10305
rect 48226 10231 48282 10240
rect 49146 10296 49202 10305
rect 49146 10231 49202 10240
rect 49790 10296 49846 10305
rect 49790 10231 49846 10240
rect 50618 10296 50674 10305
rect 50618 10231 50674 10240
rect 51354 10296 51410 10305
rect 51354 10231 51410 10240
rect 52090 10296 52146 10305
rect 52090 10231 52146 10240
rect 53010 10296 53066 10305
rect 53010 10231 53066 10240
rect 53194 10296 53250 10305
rect 53194 10231 53250 10240
rect 30380 10192 30432 10198
rect 30380 10134 30432 10140
rect 30012 9376 30064 9382
rect 30012 9318 30064 9324
rect 30392 8974 30420 10134
rect 31208 9988 31260 9994
rect 31208 9930 31260 9936
rect 30380 8968 30432 8974
rect 30380 8910 30432 8916
rect 31116 8968 31168 8974
rect 31220 8956 31248 9930
rect 31772 9178 31800 10231
rect 33048 10056 33100 10062
rect 33048 9998 33100 10004
rect 31852 9920 31904 9926
rect 31852 9862 31904 9868
rect 31760 9172 31812 9178
rect 31760 9114 31812 9120
rect 31300 9104 31352 9110
rect 31484 9104 31536 9110
rect 31352 9052 31484 9058
rect 31300 9046 31536 9052
rect 31312 9030 31524 9046
rect 31168 8928 31248 8956
rect 31116 8910 31168 8916
rect 29920 8900 29972 8906
rect 29920 8842 29972 8848
rect 30288 8832 30340 8838
rect 30288 8774 30340 8780
rect 30194 8664 30250 8673
rect 30194 8599 30196 8608
rect 30248 8599 30250 8608
rect 30196 8570 30248 8576
rect 29736 8560 29788 8566
rect 29736 8502 29788 8508
rect 30300 8498 30328 8774
rect 30288 8492 30340 8498
rect 30288 8434 30340 8440
rect 30392 1970 30420 8910
rect 31116 8832 31168 8838
rect 31116 8774 31168 8780
rect 31128 8498 31156 8774
rect 31116 8492 31168 8498
rect 31116 8434 31168 8440
rect 30932 2848 30984 2854
rect 30932 2790 30984 2796
rect 29552 1964 29604 1970
rect 29552 1906 29604 1912
rect 30380 1964 30432 1970
rect 30380 1906 30432 1912
rect 28908 1760 28960 1766
rect 28908 1702 28960 1708
rect 29736 1760 29788 1766
rect 29736 1702 29788 1708
rect 30564 1760 30616 1766
rect 30564 1702 30616 1708
rect 28920 1358 28948 1702
rect 29748 1358 29776 1702
rect 30576 1358 30604 1702
rect 30944 1494 30972 2790
rect 31220 1970 31248 8928
rect 31298 8664 31354 8673
rect 31298 8599 31300 8608
rect 31352 8599 31354 8608
rect 31300 8570 31352 8576
rect 31864 7546 31892 9862
rect 32586 9616 32642 9625
rect 32586 9551 32642 9560
rect 32680 9580 32732 9586
rect 32600 9450 32628 9551
rect 32680 9522 32732 9528
rect 32588 9444 32640 9450
rect 32588 9386 32640 9392
rect 31944 8968 31996 8974
rect 31944 8910 31996 8916
rect 31956 8634 31984 8910
rect 32496 8832 32548 8838
rect 32496 8774 32548 8780
rect 31944 8628 31996 8634
rect 31944 8570 31996 8576
rect 31852 7540 31904 7546
rect 31852 7482 31904 7488
rect 31956 2446 31984 8570
rect 32508 8498 32536 8774
rect 32692 8634 32720 9522
rect 32588 8628 32640 8634
rect 32588 8570 32640 8576
rect 32680 8628 32732 8634
rect 32680 8570 32732 8576
rect 32600 8498 32628 8570
rect 32496 8492 32548 8498
rect 32496 8434 32548 8440
rect 32588 8492 32640 8498
rect 32588 8434 32640 8440
rect 33060 6798 33088 9998
rect 34748 9276 35056 9285
rect 34748 9274 34754 9276
rect 34810 9274 34834 9276
rect 34890 9274 34914 9276
rect 34970 9274 34994 9276
rect 35050 9274 35056 9276
rect 34810 9222 34812 9274
rect 34992 9222 34994 9274
rect 34748 9220 34754 9222
rect 34810 9220 34834 9222
rect 34890 9220 34914 9222
rect 34970 9220 34994 9222
rect 35050 9220 35056 9222
rect 34748 9211 35056 9220
rect 35176 9178 35204 10231
rect 35636 9586 35664 10231
rect 36280 9586 36308 10231
rect 36924 9586 36952 10231
rect 38120 9586 38148 10231
rect 38856 9586 38884 10231
rect 39500 9586 39528 10231
rect 35624 9580 35676 9586
rect 35624 9522 35676 9528
rect 36268 9580 36320 9586
rect 36268 9522 36320 9528
rect 36912 9580 36964 9586
rect 36912 9522 36964 9528
rect 38108 9580 38160 9586
rect 38108 9522 38160 9528
rect 38844 9580 38896 9586
rect 38844 9522 38896 9528
rect 39488 9580 39540 9586
rect 39488 9522 39540 9528
rect 35808 9376 35860 9382
rect 35808 9318 35860 9324
rect 36636 9376 36688 9382
rect 36636 9318 36688 9324
rect 37096 9376 37148 9382
rect 37096 9318 37148 9324
rect 37924 9376 37976 9382
rect 37924 9318 37976 9324
rect 38108 9376 38160 9382
rect 38108 9318 38160 9324
rect 39304 9376 39356 9382
rect 39304 9318 39356 9324
rect 35164 9172 35216 9178
rect 35164 9114 35216 9120
rect 34748 8188 35056 8197
rect 34748 8186 34754 8188
rect 34810 8186 34834 8188
rect 34890 8186 34914 8188
rect 34970 8186 34994 8188
rect 35050 8186 35056 8188
rect 34810 8134 34812 8186
rect 34992 8134 34994 8186
rect 34748 8132 34754 8134
rect 34810 8132 34834 8134
rect 34890 8132 34914 8134
rect 34970 8132 34994 8134
rect 35050 8132 35056 8134
rect 34748 8123 35056 8132
rect 34748 7100 35056 7109
rect 34748 7098 34754 7100
rect 34810 7098 34834 7100
rect 34890 7098 34914 7100
rect 34970 7098 34994 7100
rect 35050 7098 35056 7100
rect 34810 7046 34812 7098
rect 34992 7046 34994 7098
rect 34748 7044 34754 7046
rect 34810 7044 34834 7046
rect 34890 7044 34914 7046
rect 34970 7044 34994 7046
rect 35050 7044 35056 7046
rect 34748 7035 35056 7044
rect 33048 6792 33100 6798
rect 33048 6734 33100 6740
rect 34748 6012 35056 6021
rect 34748 6010 34754 6012
rect 34810 6010 34834 6012
rect 34890 6010 34914 6012
rect 34970 6010 34994 6012
rect 35050 6010 35056 6012
rect 34810 5958 34812 6010
rect 34992 5958 34994 6010
rect 34748 5956 34754 5958
rect 34810 5956 34834 5958
rect 34890 5956 34914 5958
rect 34970 5956 34994 5958
rect 35050 5956 35056 5958
rect 34748 5947 35056 5956
rect 33232 5772 33284 5778
rect 33232 5714 33284 5720
rect 33244 5030 33272 5714
rect 34612 5364 34664 5370
rect 34612 5306 34664 5312
rect 33232 5024 33284 5030
rect 33232 4966 33284 4972
rect 34624 4758 34652 5306
rect 34748 4924 35056 4933
rect 34748 4922 34754 4924
rect 34810 4922 34834 4924
rect 34890 4922 34914 4924
rect 34970 4922 34994 4924
rect 35050 4922 35056 4924
rect 34810 4870 34812 4922
rect 34992 4870 34994 4922
rect 34748 4868 34754 4870
rect 34810 4868 34834 4870
rect 34890 4868 34914 4870
rect 34970 4868 34994 4870
rect 35050 4868 35056 4870
rect 34748 4859 35056 4868
rect 34612 4752 34664 4758
rect 34612 4694 34664 4700
rect 33140 4684 33192 4690
rect 33140 4626 33192 4632
rect 33152 2582 33180 4626
rect 34748 3836 35056 3845
rect 34748 3834 34754 3836
rect 34810 3834 34834 3836
rect 34890 3834 34914 3836
rect 34970 3834 34994 3836
rect 35050 3834 35056 3836
rect 34810 3782 34812 3834
rect 34992 3782 34994 3834
rect 34748 3780 34754 3782
rect 34810 3780 34834 3782
rect 34890 3780 34914 3782
rect 34970 3780 34994 3782
rect 35050 3780 35056 3782
rect 34748 3771 35056 3780
rect 34748 2748 35056 2757
rect 34748 2746 34754 2748
rect 34810 2746 34834 2748
rect 34890 2746 34914 2748
rect 34970 2746 34994 2748
rect 35050 2746 35056 2748
rect 34810 2694 34812 2746
rect 34992 2694 34994 2746
rect 34748 2692 34754 2694
rect 34810 2692 34834 2694
rect 34890 2692 34914 2694
rect 34970 2692 34994 2694
rect 35050 2692 35056 2694
rect 34748 2683 35056 2692
rect 33140 2576 33192 2582
rect 33140 2518 33192 2524
rect 31944 2440 31996 2446
rect 31944 2382 31996 2388
rect 32496 2440 32548 2446
rect 32496 2382 32548 2388
rect 32312 2304 32364 2310
rect 32312 2246 32364 2252
rect 31208 1964 31260 1970
rect 31208 1906 31260 1912
rect 31024 1896 31076 1902
rect 31024 1838 31076 1844
rect 31036 1494 31064 1838
rect 31760 1760 31812 1766
rect 31760 1702 31812 1708
rect 30932 1488 30984 1494
rect 30932 1430 30984 1436
rect 31024 1488 31076 1494
rect 31024 1430 31076 1436
rect 31772 1358 31800 1702
rect 32324 1358 32352 2246
rect 32508 1970 32536 2382
rect 35624 2372 35676 2378
rect 35624 2314 35676 2320
rect 33048 2304 33100 2310
rect 33048 2246 33100 2252
rect 33060 2038 33088 2246
rect 33048 2032 33100 2038
rect 33048 1974 33100 1980
rect 35532 2032 35584 2038
rect 35532 1974 35584 1980
rect 32496 1964 32548 1970
rect 32496 1906 32548 1912
rect 33140 1760 33192 1766
rect 33140 1702 33192 1708
rect 33152 1465 33180 1702
rect 34748 1660 35056 1669
rect 34748 1658 34754 1660
rect 34810 1658 34834 1660
rect 34890 1658 34914 1660
rect 34970 1658 34994 1660
rect 35050 1658 35056 1660
rect 34810 1606 34812 1658
rect 34992 1606 34994 1658
rect 34748 1604 34754 1606
rect 34810 1604 34834 1606
rect 34890 1604 34914 1606
rect 34970 1604 34994 1606
rect 35050 1604 35056 1606
rect 34748 1595 35056 1604
rect 35544 1562 35572 1974
rect 35636 1562 35664 2314
rect 35820 2038 35848 9318
rect 36360 8560 36412 8566
rect 36360 8502 36412 8508
rect 35898 6488 35954 6497
rect 35898 6423 35954 6432
rect 35912 4826 35940 6423
rect 35900 4820 35952 4826
rect 35900 4762 35952 4768
rect 35900 3392 35952 3398
rect 35900 3334 35952 3340
rect 36084 3392 36136 3398
rect 36084 3334 36136 3340
rect 35912 3126 35940 3334
rect 35900 3120 35952 3126
rect 35900 3062 35952 3068
rect 35808 2032 35860 2038
rect 35808 1974 35860 1980
rect 35532 1556 35584 1562
rect 35532 1498 35584 1504
rect 35624 1556 35676 1562
rect 35624 1498 35676 1504
rect 33138 1456 33194 1465
rect 33138 1391 33194 1400
rect 34428 1420 34480 1426
rect 34428 1362 34480 1368
rect 28908 1352 28960 1358
rect 28908 1294 28960 1300
rect 29736 1352 29788 1358
rect 29736 1294 29788 1300
rect 30564 1352 30616 1358
rect 30564 1294 30616 1300
rect 31760 1352 31812 1358
rect 31760 1294 31812 1300
rect 32312 1352 32364 1358
rect 32312 1294 32364 1300
rect 29000 1216 29052 1222
rect 29000 1158 29052 1164
rect 29920 1216 29972 1222
rect 29920 1158 29972 1164
rect 30380 1216 30432 1222
rect 30380 1158 30432 1164
rect 31576 1216 31628 1222
rect 31576 1158 31628 1164
rect 32496 1216 32548 1222
rect 32496 1158 32548 1164
rect 29012 649 29040 1158
rect 28998 640 29054 649
rect 28998 575 29054 584
rect 29932 513 29960 1158
rect 30392 649 30420 1158
rect 30378 640 30434 649
rect 30378 575 30434 584
rect 17960 478 18012 484
rect 28722 504 28778 513
rect 28722 439 28778 448
rect 29918 504 29974 513
rect 29918 439 29974 448
rect 31588 377 31616 1158
rect 32508 513 32536 1158
rect 32494 504 32550 513
rect 32494 439 32550 448
rect 34440 377 34468 1362
rect 35624 1352 35676 1358
rect 35624 1294 35676 1300
rect 35636 649 35664 1294
rect 36096 1222 36124 3334
rect 36372 2038 36400 8502
rect 36544 6384 36596 6390
rect 36544 6326 36596 6332
rect 36556 5914 36584 6326
rect 36544 5908 36596 5914
rect 36544 5850 36596 5856
rect 36544 4616 36596 4622
rect 36544 4558 36596 4564
rect 36556 4010 36584 4558
rect 36544 4004 36596 4010
rect 36544 3946 36596 3952
rect 36452 3732 36504 3738
rect 36452 3674 36504 3680
rect 36464 2378 36492 3674
rect 36648 3534 36676 9318
rect 37004 8900 37056 8906
rect 37004 8842 37056 8848
rect 37016 7274 37044 8842
rect 37004 7268 37056 7274
rect 37004 7210 37056 7216
rect 36636 3528 36688 3534
rect 36636 3470 36688 3476
rect 36636 2508 36688 2514
rect 36636 2450 36688 2456
rect 36452 2372 36504 2378
rect 36452 2314 36504 2320
rect 36648 2038 36676 2450
rect 37108 2378 37136 9318
rect 37936 5302 37964 9318
rect 37832 5296 37884 5302
rect 37832 5238 37884 5244
rect 37924 5296 37976 5302
rect 37924 5238 37976 5244
rect 37556 3596 37608 3602
rect 37556 3538 37608 3544
rect 37280 3528 37332 3534
rect 37568 3482 37596 3538
rect 37280 3470 37332 3476
rect 37188 3052 37240 3058
rect 37188 2994 37240 3000
rect 37200 2514 37228 2994
rect 37188 2508 37240 2514
rect 37188 2450 37240 2456
rect 37096 2372 37148 2378
rect 37096 2314 37148 2320
rect 36728 2304 36780 2310
rect 36728 2246 36780 2252
rect 36360 2032 36412 2038
rect 36360 1974 36412 1980
rect 36636 2032 36688 2038
rect 36636 1974 36688 1980
rect 36740 1494 36768 2246
rect 37200 1902 37228 2450
rect 37292 2378 37320 3470
rect 37476 3454 37596 3482
rect 37476 2854 37504 3454
rect 37556 3392 37608 3398
rect 37556 3334 37608 3340
rect 37568 3194 37596 3334
rect 37556 3188 37608 3194
rect 37556 3130 37608 3136
rect 37464 2848 37516 2854
rect 37464 2790 37516 2796
rect 37280 2372 37332 2378
rect 37280 2314 37332 2320
rect 37292 2038 37320 2314
rect 37740 2304 37792 2310
rect 37740 2246 37792 2252
rect 37280 2032 37332 2038
rect 37280 1974 37332 1980
rect 37188 1896 37240 1902
rect 37188 1838 37240 1844
rect 36820 1760 36872 1766
rect 36818 1728 36820 1737
rect 36872 1728 36874 1737
rect 36818 1663 36874 1672
rect 36728 1488 36780 1494
rect 36728 1430 36780 1436
rect 36268 1352 36320 1358
rect 36268 1294 36320 1300
rect 36912 1352 36964 1358
rect 36912 1294 36964 1300
rect 36084 1216 36136 1222
rect 36084 1158 36136 1164
rect 36280 649 36308 1294
rect 36924 649 36952 1294
rect 35622 640 35678 649
rect 35622 575 35678 584
rect 36266 640 36322 649
rect 36266 575 36322 584
rect 36910 640 36966 649
rect 36910 575 36966 584
rect 37752 406 37780 2246
rect 37844 1834 37872 5238
rect 38120 3126 38148 9318
rect 38568 6724 38620 6730
rect 38568 6666 38620 6672
rect 38200 5228 38252 5234
rect 38200 5170 38252 5176
rect 38212 3126 38240 5170
rect 38476 5160 38528 5166
rect 38476 5102 38528 5108
rect 38488 3466 38516 5102
rect 38476 3460 38528 3466
rect 38476 3402 38528 3408
rect 38016 3120 38068 3126
rect 38016 3062 38068 3068
rect 38108 3120 38160 3126
rect 38108 3062 38160 3068
rect 38200 3120 38252 3126
rect 38200 3062 38252 3068
rect 37832 1828 37884 1834
rect 37832 1770 37884 1776
rect 38028 1222 38056 3062
rect 38212 2774 38240 3062
rect 38488 3058 38516 3402
rect 38580 3126 38608 6666
rect 38752 5296 38804 5302
rect 38752 5238 38804 5244
rect 38660 3392 38712 3398
rect 38660 3334 38712 3340
rect 38568 3120 38620 3126
rect 38568 3062 38620 3068
rect 38476 3052 38528 3058
rect 38476 2994 38528 3000
rect 38212 2746 38332 2774
rect 38198 2408 38254 2417
rect 38198 2343 38254 2352
rect 38212 2310 38240 2343
rect 38200 2304 38252 2310
rect 38200 2246 38252 2252
rect 38304 1970 38332 2746
rect 38672 2446 38700 3334
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 38660 2032 38712 2038
rect 38660 1974 38712 1980
rect 38108 1964 38160 1970
rect 38108 1906 38160 1912
rect 38292 1964 38344 1970
rect 38292 1906 38344 1912
rect 38016 1216 38068 1222
rect 38016 1158 38068 1164
rect 38120 649 38148 1906
rect 38672 1494 38700 1974
rect 38660 1488 38712 1494
rect 38660 1430 38712 1436
rect 38568 1352 38620 1358
rect 38568 1294 38620 1300
rect 38580 649 38608 1294
rect 38764 814 38792 5238
rect 38936 4140 38988 4146
rect 38936 4082 38988 4088
rect 38948 3126 38976 4082
rect 39118 3496 39174 3505
rect 39118 3431 39174 3440
rect 38936 3120 38988 3126
rect 38936 3062 38988 3068
rect 39132 2922 39160 3431
rect 39120 2916 39172 2922
rect 39120 2858 39172 2864
rect 39316 2038 39344 9318
rect 40328 8974 40356 10231
rect 40788 9586 40816 10231
rect 41432 9586 41460 10231
rect 42076 9586 42104 10231
rect 43272 9586 43300 10231
rect 44008 9586 44036 10231
rect 44652 9586 44680 10231
rect 40776 9580 40828 9586
rect 40776 9522 40828 9528
rect 41420 9580 41472 9586
rect 41420 9522 41472 9528
rect 42064 9580 42116 9586
rect 42064 9522 42116 9528
rect 43260 9580 43312 9586
rect 43260 9522 43312 9528
rect 43996 9580 44048 9586
rect 43996 9522 44048 9528
rect 44640 9580 44692 9586
rect 44640 9522 44692 9528
rect 40868 9376 40920 9382
rect 40868 9318 40920 9324
rect 41696 9376 41748 9382
rect 41696 9318 41748 9324
rect 41880 9376 41932 9382
rect 41880 9318 41932 9324
rect 43260 9376 43312 9382
rect 43260 9318 43312 9324
rect 43352 9376 43404 9382
rect 43904 9376 43956 9382
rect 43352 9318 43404 9324
rect 43548 9336 43904 9364
rect 40316 8968 40368 8974
rect 40316 8910 40368 8916
rect 40132 8832 40184 8838
rect 40132 8774 40184 8780
rect 39764 4752 39816 4758
rect 39764 4694 39816 4700
rect 39776 2038 39804 4694
rect 39948 3732 40000 3738
rect 39948 3674 40000 3680
rect 39856 3120 39908 3126
rect 39856 3062 39908 3068
rect 39304 2032 39356 2038
rect 39304 1974 39356 1980
rect 39764 2032 39816 2038
rect 39764 1974 39816 1980
rect 38844 1352 38896 1358
rect 38844 1294 38896 1300
rect 38752 808 38804 814
rect 38752 750 38804 756
rect 38106 640 38162 649
rect 38106 575 38162 584
rect 38566 640 38622 649
rect 38566 575 38622 584
rect 37740 400 37792 406
rect 31574 368 31630 377
rect 9404 332 9456 338
rect 31574 303 31630 312
rect 34426 368 34482 377
rect 38856 377 38884 1294
rect 39868 1222 39896 3062
rect 39960 3058 39988 3674
rect 40040 3664 40092 3670
rect 40040 3606 40092 3612
rect 39948 3052 40000 3058
rect 39948 2994 40000 3000
rect 39960 1970 39988 2994
rect 40052 2378 40080 3606
rect 40144 3126 40172 8774
rect 40500 6248 40552 6254
rect 40500 6190 40552 6196
rect 40316 5024 40368 5030
rect 40316 4966 40368 4972
rect 40328 4486 40356 4966
rect 40316 4480 40368 4486
rect 40316 4422 40368 4428
rect 40224 4208 40276 4214
rect 40224 4150 40276 4156
rect 40132 3120 40184 3126
rect 40132 3062 40184 3068
rect 40236 3058 40264 4150
rect 40224 3052 40276 3058
rect 40224 2994 40276 3000
rect 40236 2774 40264 2994
rect 40144 2746 40264 2774
rect 40040 2372 40092 2378
rect 40040 2314 40092 2320
rect 40144 2258 40172 2746
rect 40328 2666 40356 4422
rect 40408 3936 40460 3942
rect 40408 3878 40460 3884
rect 40420 3398 40448 3878
rect 40408 3392 40460 3398
rect 40408 3334 40460 3340
rect 40512 3126 40540 6190
rect 40776 5160 40828 5166
rect 40776 5102 40828 5108
rect 40592 4208 40644 4214
rect 40592 4150 40644 4156
rect 40500 3120 40552 3126
rect 40500 3062 40552 3068
rect 40052 2230 40172 2258
rect 40236 2638 40356 2666
rect 40052 2038 40080 2230
rect 40040 2032 40092 2038
rect 40040 1974 40092 1980
rect 40132 2032 40184 2038
rect 40132 1974 40184 1980
rect 39948 1964 40000 1970
rect 39948 1906 40000 1912
rect 39948 1352 40000 1358
rect 39948 1294 40000 1300
rect 39856 1216 39908 1222
rect 39856 1158 39908 1164
rect 39960 649 39988 1294
rect 39946 640 40002 649
rect 39946 575 40002 584
rect 40144 474 40172 1974
rect 40236 610 40264 2638
rect 40314 1864 40370 1873
rect 40314 1799 40316 1808
rect 40368 1799 40370 1808
rect 40316 1770 40368 1776
rect 40604 1222 40632 4150
rect 40788 4078 40816 5102
rect 40880 4146 40908 9318
rect 41236 9172 41288 9178
rect 41236 9114 41288 9120
rect 41144 5160 41196 5166
rect 41144 5102 41196 5108
rect 40960 4820 41012 4826
rect 40960 4762 41012 4768
rect 40972 4706 41000 4762
rect 40972 4678 41092 4706
rect 41156 4690 41184 5102
rect 40960 4480 41012 4486
rect 40960 4422 41012 4428
rect 40972 4321 41000 4422
rect 40958 4312 41014 4321
rect 40958 4247 41014 4256
rect 41064 4146 41092 4678
rect 41144 4684 41196 4690
rect 41144 4626 41196 4632
rect 41248 4554 41276 9114
rect 41328 5568 41380 5574
rect 41328 5510 41380 5516
rect 41340 5250 41368 5510
rect 41340 5222 41644 5250
rect 41236 4548 41288 4554
rect 41236 4490 41288 4496
rect 41340 4434 41368 5222
rect 41616 4554 41644 5222
rect 41604 4548 41656 4554
rect 41604 4490 41656 4496
rect 41248 4406 41368 4434
rect 41248 4214 41276 4406
rect 41418 4312 41474 4321
rect 41418 4247 41474 4256
rect 41236 4208 41288 4214
rect 41236 4150 41288 4156
rect 40868 4140 40920 4146
rect 40868 4082 40920 4088
rect 41052 4140 41104 4146
rect 41052 4082 41104 4088
rect 40776 4072 40828 4078
rect 40776 4014 40828 4020
rect 40788 3670 40816 4014
rect 40776 3664 40828 3670
rect 40776 3606 40828 3612
rect 40788 3058 40816 3606
rect 40960 3460 41012 3466
rect 40960 3402 41012 3408
rect 40776 3052 40828 3058
rect 40776 2994 40828 3000
rect 40972 2990 41000 3402
rect 41236 3392 41288 3398
rect 41236 3334 41288 3340
rect 41052 3120 41104 3126
rect 41052 3062 41104 3068
rect 40960 2984 41012 2990
rect 40960 2926 41012 2932
rect 40776 1352 40828 1358
rect 40776 1294 40828 1300
rect 40592 1216 40644 1222
rect 40592 1158 40644 1164
rect 40788 649 40816 1294
rect 40774 640 40830 649
rect 40224 604 40276 610
rect 40774 575 40830 584
rect 40224 546 40276 552
rect 40132 468 40184 474
rect 40132 410 40184 416
rect 37740 342 37792 348
rect 38842 368 38898 377
rect 34426 303 34482 312
rect 41064 338 41092 3062
rect 41142 2952 41198 2961
rect 41142 2887 41144 2896
rect 41196 2887 41198 2896
rect 41144 2858 41196 2864
rect 41248 1222 41276 3334
rect 41432 1476 41460 4247
rect 41616 3466 41644 4490
rect 41512 3460 41564 3466
rect 41512 3402 41564 3408
rect 41604 3460 41656 3466
rect 41604 3402 41656 3408
rect 41524 3346 41552 3402
rect 41708 3346 41736 9318
rect 41892 9178 41920 9318
rect 41880 9172 41932 9178
rect 41880 9114 41932 9120
rect 41972 7540 42024 7546
rect 41972 7482 42024 7488
rect 41880 3936 41932 3942
rect 41880 3878 41932 3884
rect 41524 3318 41736 3346
rect 41892 3126 41920 3878
rect 41984 3466 42012 7482
rect 42616 6724 42668 6730
rect 42616 6666 42668 6672
rect 42628 6458 42656 6666
rect 42616 6452 42668 6458
rect 42616 6394 42668 6400
rect 42984 6384 43036 6390
rect 42984 6326 43036 6332
rect 42524 6180 42576 6186
rect 42524 6122 42576 6128
rect 42064 5636 42116 5642
rect 42064 5578 42116 5584
rect 42076 5409 42104 5578
rect 42062 5400 42118 5409
rect 42062 5335 42118 5344
rect 42432 5160 42484 5166
rect 42430 5128 42432 5137
rect 42484 5128 42486 5137
rect 42430 5063 42486 5072
rect 42064 5024 42116 5030
rect 42536 5001 42564 6122
rect 42800 5908 42852 5914
rect 42800 5850 42852 5856
rect 42708 5704 42760 5710
rect 42706 5672 42708 5681
rect 42760 5672 42762 5681
rect 42706 5607 42762 5616
rect 42812 5386 42840 5850
rect 42720 5358 42840 5386
rect 42616 5228 42668 5234
rect 42616 5170 42668 5176
rect 42064 4966 42116 4972
rect 42522 4992 42578 5001
rect 42076 4554 42104 4966
rect 42522 4927 42578 4936
rect 42536 4826 42564 4927
rect 42524 4820 42576 4826
rect 42524 4762 42576 4768
rect 42246 4584 42302 4593
rect 42064 4548 42116 4554
rect 42246 4519 42302 4528
rect 42064 4490 42116 4496
rect 42260 4486 42288 4519
rect 42248 4480 42300 4486
rect 42248 4422 42300 4428
rect 42628 4214 42656 5170
rect 42720 5114 42748 5358
rect 42720 5086 42840 5114
rect 42616 4208 42668 4214
rect 42616 4150 42668 4156
rect 42812 3942 42840 5086
rect 42892 5092 42944 5098
rect 42892 5034 42944 5040
rect 42904 4282 42932 5034
rect 42892 4276 42944 4282
rect 42892 4218 42944 4224
rect 42800 3936 42852 3942
rect 42800 3878 42852 3884
rect 41972 3460 42024 3466
rect 41972 3402 42024 3408
rect 41880 3120 41932 3126
rect 41880 3062 41932 3068
rect 41432 1448 41552 1476
rect 41420 1352 41472 1358
rect 41420 1294 41472 1300
rect 41236 1216 41288 1222
rect 41236 1158 41288 1164
rect 41432 649 41460 1294
rect 41524 1222 41552 1448
rect 42064 1352 42116 1358
rect 42064 1294 42116 1300
rect 41512 1216 41564 1222
rect 41512 1158 41564 1164
rect 42076 649 42104 1294
rect 42996 1290 43024 6326
rect 43168 6316 43220 6322
rect 43168 6258 43220 6264
rect 43180 5817 43208 6258
rect 43166 5808 43222 5817
rect 43166 5743 43222 5752
rect 43272 4622 43300 9318
rect 43364 6390 43392 9318
rect 43444 8832 43496 8838
rect 43444 8774 43496 8780
rect 43352 6384 43404 6390
rect 43352 6326 43404 6332
rect 43456 5710 43484 8774
rect 43444 5704 43496 5710
rect 43444 5646 43496 5652
rect 43548 5370 43576 9336
rect 43904 9318 43956 9324
rect 45480 8974 45508 10231
rect 45940 9586 45968 10231
rect 46204 9648 46256 9654
rect 46256 9596 46336 9602
rect 46204 9590 46336 9596
rect 45928 9580 45980 9586
rect 46216 9574 46336 9590
rect 46584 9586 46612 10231
rect 47228 9586 47256 10231
rect 48240 9586 48268 10231
rect 49160 9586 49188 10231
rect 49804 9586 49832 10231
rect 50632 9586 50660 10231
rect 51080 9716 51132 9722
rect 51080 9658 51132 9664
rect 45928 9522 45980 9528
rect 46308 9518 46336 9574
rect 46572 9580 46624 9586
rect 46572 9522 46624 9528
rect 47216 9580 47268 9586
rect 47216 9522 47268 9528
rect 48228 9580 48280 9586
rect 48228 9522 48280 9528
rect 49148 9580 49200 9586
rect 49148 9522 49200 9528
rect 49792 9580 49844 9586
rect 49792 9522 49844 9528
rect 50620 9580 50672 9586
rect 50620 9522 50672 9528
rect 46296 9512 46348 9518
rect 46296 9454 46348 9460
rect 46204 9444 46256 9450
rect 46204 9386 46256 9392
rect 47768 9444 47820 9450
rect 47768 9386 47820 9392
rect 45560 9376 45612 9382
rect 45560 9318 45612 9324
rect 46112 9376 46164 9382
rect 46112 9318 46164 9324
rect 45468 8968 45520 8974
rect 45468 8910 45520 8916
rect 43996 6792 44048 6798
rect 43996 6734 44048 6740
rect 43904 6656 43956 6662
rect 43904 6598 43956 6604
rect 43916 6390 43944 6598
rect 43904 6384 43956 6390
rect 43904 6326 43956 6332
rect 43626 5808 43682 5817
rect 43626 5743 43682 5752
rect 43640 5710 43668 5743
rect 43628 5704 43680 5710
rect 43720 5704 43772 5710
rect 43628 5646 43680 5652
rect 43718 5672 43720 5681
rect 43772 5672 43774 5681
rect 43536 5364 43588 5370
rect 43536 5306 43588 5312
rect 43352 5296 43404 5302
rect 43352 5238 43404 5244
rect 43640 5284 43668 5646
rect 43718 5607 43774 5616
rect 43720 5296 43772 5302
rect 43640 5256 43720 5284
rect 43260 4616 43312 4622
rect 43260 4558 43312 4564
rect 43076 4480 43128 4486
rect 43076 4422 43128 4428
rect 42984 1284 43036 1290
rect 42984 1226 43036 1232
rect 43088 1222 43116 4422
rect 43364 1494 43392 5238
rect 43640 4622 43668 5256
rect 43720 5238 43772 5244
rect 43812 5228 43864 5234
rect 43812 5170 43864 5176
rect 43824 5001 43852 5170
rect 43810 4992 43866 5001
rect 43810 4927 43866 4936
rect 43628 4616 43680 4622
rect 43628 4558 43680 4564
rect 43352 1488 43404 1494
rect 43352 1430 43404 1436
rect 43260 1352 43312 1358
rect 43260 1294 43312 1300
rect 43076 1216 43128 1222
rect 43076 1158 43128 1164
rect 43272 649 43300 1294
rect 43916 678 43944 6326
rect 44008 4554 44036 6734
rect 45572 6390 45600 9318
rect 45928 9104 45980 9110
rect 45928 9046 45980 9052
rect 45744 7948 45796 7954
rect 45744 7890 45796 7896
rect 45756 6390 45784 7890
rect 45008 6384 45060 6390
rect 45008 6326 45060 6332
rect 45560 6384 45612 6390
rect 45560 6326 45612 6332
rect 45744 6384 45796 6390
rect 45744 6326 45796 6332
rect 44732 6248 44784 6254
rect 44086 6216 44142 6225
rect 44732 6190 44784 6196
rect 44086 6151 44088 6160
rect 44140 6151 44142 6160
rect 44088 6122 44140 6128
rect 44744 5778 44772 6190
rect 44732 5772 44784 5778
rect 44732 5714 44784 5720
rect 44364 5704 44416 5710
rect 44284 5664 44364 5692
rect 44284 5137 44312 5664
rect 44364 5646 44416 5652
rect 44546 5672 44602 5681
rect 44546 5607 44602 5616
rect 44560 5574 44588 5607
rect 44456 5568 44508 5574
rect 44456 5510 44508 5516
rect 44548 5568 44600 5574
rect 44548 5510 44600 5516
rect 44364 5296 44416 5302
rect 44364 5238 44416 5244
rect 44468 5250 44496 5510
rect 44270 5128 44326 5137
rect 44270 5063 44326 5072
rect 43996 4548 44048 4554
rect 43996 4490 44048 4496
rect 44272 4480 44324 4486
rect 44272 4422 44324 4428
rect 44284 4321 44312 4422
rect 44270 4312 44326 4321
rect 44270 4247 44326 4256
rect 43996 1352 44048 1358
rect 43996 1294 44048 1300
rect 43904 672 43956 678
rect 41418 640 41474 649
rect 41418 575 41474 584
rect 42062 640 42118 649
rect 42062 575 42118 584
rect 43258 640 43314 649
rect 44008 649 44036 1294
rect 44376 1057 44404 5238
rect 44468 5222 44588 5250
rect 44560 1834 44588 5222
rect 44744 5166 44772 5714
rect 44732 5160 44784 5166
rect 44638 5128 44694 5137
rect 44732 5102 44784 5108
rect 44638 5063 44640 5072
rect 44692 5063 44694 5072
rect 44640 5034 44692 5040
rect 44744 4690 44772 5102
rect 44732 4684 44784 4690
rect 44732 4626 44784 4632
rect 44548 1828 44600 1834
rect 44548 1770 44600 1776
rect 44640 1352 44692 1358
rect 44640 1294 44692 1300
rect 44362 1048 44418 1057
rect 44362 983 44418 992
rect 44652 649 44680 1294
rect 45020 1222 45048 6326
rect 45376 6316 45428 6322
rect 45376 6258 45428 6264
rect 45388 5817 45416 6258
rect 45374 5808 45430 5817
rect 45374 5743 45430 5752
rect 45388 5370 45416 5743
rect 45376 5364 45428 5370
rect 45376 5306 45428 5312
rect 45836 5296 45888 5302
rect 45836 5238 45888 5244
rect 45468 1964 45520 1970
rect 45468 1906 45520 1912
rect 45008 1216 45060 1222
rect 45008 1158 45060 1164
rect 45480 649 45508 1906
rect 45848 1222 45876 5238
rect 45940 5234 45968 9046
rect 46018 6488 46074 6497
rect 46018 6423 46020 6432
rect 46072 6423 46074 6432
rect 46020 6394 46072 6400
rect 46020 6248 46072 6254
rect 46020 6190 46072 6196
rect 46032 5778 46060 6190
rect 46020 5772 46072 5778
rect 46020 5714 46072 5720
rect 46124 5302 46152 9318
rect 46216 9110 46244 9386
rect 46848 9376 46900 9382
rect 46848 9318 46900 9324
rect 47124 9376 47176 9382
rect 47124 9318 47176 9324
rect 46204 9104 46256 9110
rect 46204 9046 46256 9052
rect 46860 5710 46888 9318
rect 46848 5704 46900 5710
rect 46848 5646 46900 5652
rect 46940 5704 46992 5710
rect 46940 5646 46992 5652
rect 46664 5568 46716 5574
rect 46664 5510 46716 5516
rect 46112 5296 46164 5302
rect 46112 5238 46164 5244
rect 46296 5296 46348 5302
rect 46296 5238 46348 5244
rect 45928 5228 45980 5234
rect 45928 5170 45980 5176
rect 45928 1352 45980 1358
rect 45928 1294 45980 1300
rect 45836 1216 45888 1222
rect 45836 1158 45888 1164
rect 45940 649 45968 1294
rect 46308 746 46336 5238
rect 46676 4162 46704 5510
rect 46848 5364 46900 5370
rect 46952 5352 46980 5646
rect 46900 5324 46980 5352
rect 46848 5306 46900 5312
rect 46860 4554 46888 5306
rect 46848 4548 46900 4554
rect 46848 4490 46900 4496
rect 46940 4480 46992 4486
rect 46938 4448 46940 4457
rect 46992 4448 46994 4457
rect 46938 4383 46994 4392
rect 46676 4134 46888 4162
rect 46664 3460 46716 3466
rect 46664 3402 46716 3408
rect 46572 1352 46624 1358
rect 46572 1294 46624 1300
rect 46296 740 46348 746
rect 46296 682 46348 688
rect 46584 649 46612 1294
rect 46676 1290 46704 3402
rect 46664 1284 46716 1290
rect 46664 1226 46716 1232
rect 46860 1222 46888 4134
rect 46940 3460 46992 3466
rect 47136 3448 47164 9318
rect 47308 8084 47360 8090
rect 47308 8026 47360 8032
rect 47320 5710 47348 8026
rect 47584 6248 47636 6254
rect 47584 6190 47636 6196
rect 47596 5778 47624 6190
rect 47584 5772 47636 5778
rect 47584 5714 47636 5720
rect 47308 5704 47360 5710
rect 47308 5646 47360 5652
rect 47676 5568 47728 5574
rect 47676 5510 47728 5516
rect 47216 4548 47268 4554
rect 47216 4490 47268 4496
rect 47228 3466 47256 4490
rect 47400 3936 47452 3942
rect 47400 3878 47452 3884
rect 47412 3466 47440 3878
rect 46992 3420 47164 3448
rect 47216 3460 47268 3466
rect 46940 3402 46992 3408
rect 47216 3402 47268 3408
rect 47400 3460 47452 3466
rect 47400 3402 47452 3408
rect 47216 1352 47268 1358
rect 47216 1294 47268 1300
rect 46848 1216 46900 1222
rect 46848 1158 46900 1164
rect 47228 649 47256 1294
rect 47688 1018 47716 5510
rect 47780 4622 47808 9386
rect 49240 9376 49292 9382
rect 49240 9318 49292 9324
rect 50436 9376 50488 9382
rect 50436 9318 50488 9324
rect 48228 8016 48280 8022
rect 48228 7958 48280 7964
rect 47860 6792 47912 6798
rect 47860 6734 47912 6740
rect 47872 5914 47900 6734
rect 47860 5908 47912 5914
rect 47860 5850 47912 5856
rect 48044 5772 48096 5778
rect 48044 5714 48096 5720
rect 47950 5400 48006 5409
rect 47950 5335 48006 5344
rect 47964 5234 47992 5335
rect 47952 5228 48004 5234
rect 47952 5170 48004 5176
rect 48056 5166 48084 5714
rect 48044 5160 48096 5166
rect 48044 5102 48096 5108
rect 47860 5024 47912 5030
rect 47860 4966 47912 4972
rect 47768 4616 47820 4622
rect 47768 4558 47820 4564
rect 47872 4554 47900 4966
rect 48056 4690 48084 5102
rect 48044 4684 48096 4690
rect 48044 4626 48096 4632
rect 47860 4548 47912 4554
rect 47860 4490 47912 4496
rect 48056 4214 48084 4626
rect 48136 4616 48188 4622
rect 48136 4558 48188 4564
rect 48148 4457 48176 4558
rect 48240 4554 48268 7958
rect 48228 4548 48280 4554
rect 48228 4490 48280 4496
rect 48872 4548 48924 4554
rect 48872 4490 48924 4496
rect 48596 4480 48648 4486
rect 48134 4448 48190 4457
rect 48596 4422 48648 4428
rect 48134 4383 48190 4392
rect 48608 4282 48636 4422
rect 48596 4276 48648 4282
rect 48596 4218 48648 4224
rect 48044 4208 48096 4214
rect 48044 4150 48096 4156
rect 48056 3602 48084 4150
rect 48044 3596 48096 3602
rect 48044 3538 48096 3544
rect 48320 1352 48372 1358
rect 48320 1294 48372 1300
rect 47676 1012 47728 1018
rect 47676 954 47728 960
rect 48332 649 48360 1294
rect 48884 1222 48912 4490
rect 49056 4276 49108 4282
rect 49056 4218 49108 4224
rect 49068 2009 49096 4218
rect 49252 4214 49280 9318
rect 49884 6724 49936 6730
rect 49884 6666 49936 6672
rect 49332 5228 49384 5234
rect 49332 5170 49384 5176
rect 49344 4214 49372 5170
rect 49896 4214 49924 6666
rect 50448 5710 50476 9318
rect 51092 5710 51120 9658
rect 51368 9586 51396 10231
rect 52104 9586 52132 10231
rect 53024 9586 53052 10231
rect 51356 9580 51408 9586
rect 51356 9522 51408 9528
rect 52092 9580 52144 9586
rect 52092 9522 52144 9528
rect 53012 9580 53064 9586
rect 53012 9522 53064 9528
rect 51172 9376 51224 9382
rect 51172 9318 51224 9324
rect 51264 9376 51316 9382
rect 51264 9318 51316 9324
rect 52276 9376 52328 9382
rect 52276 9318 52328 9324
rect 50436 5704 50488 5710
rect 50436 5646 50488 5652
rect 51080 5704 51132 5710
rect 51080 5646 51132 5652
rect 50988 5636 51040 5642
rect 50988 5578 51040 5584
rect 50528 5568 50580 5574
rect 50528 5510 50580 5516
rect 49148 4208 49200 4214
rect 49148 4150 49200 4156
rect 49240 4208 49292 4214
rect 49240 4150 49292 4156
rect 49332 4208 49384 4214
rect 49332 4150 49384 4156
rect 49884 4208 49936 4214
rect 49884 4150 49936 4156
rect 49160 2774 49188 4150
rect 49792 4072 49844 4078
rect 49790 4040 49792 4049
rect 49844 4040 49846 4049
rect 49790 3975 49846 3984
rect 49160 2746 49648 2774
rect 49054 2000 49110 2009
rect 49054 1935 49110 1944
rect 49148 1352 49200 1358
rect 49148 1294 49200 1300
rect 48872 1216 48924 1222
rect 48872 1158 48924 1164
rect 49160 649 49188 1294
rect 49620 1222 49648 2746
rect 50540 1834 50568 5510
rect 50712 5296 50764 5302
rect 50712 5238 50764 5244
rect 50620 1964 50672 1970
rect 50620 1906 50672 1912
rect 50528 1828 50580 1834
rect 50528 1770 50580 1776
rect 49792 1352 49844 1358
rect 49792 1294 49844 1300
rect 49608 1216 49660 1222
rect 49608 1158 49660 1164
rect 49804 649 49832 1294
rect 50632 649 50660 1906
rect 50724 1222 50752 5238
rect 51000 5234 51028 5578
rect 51184 5302 51212 9318
rect 51172 5296 51224 5302
rect 51172 5238 51224 5244
rect 50988 5228 51040 5234
rect 50988 5170 51040 5176
rect 51000 4486 51028 5170
rect 51172 4752 51224 4758
rect 51172 4694 51224 4700
rect 50988 4480 51040 4486
rect 50988 4422 51040 4428
rect 51184 4282 51212 4694
rect 51172 4276 51224 4282
rect 51172 4218 51224 4224
rect 51276 4146 51304 9318
rect 51356 8288 51408 8294
rect 51356 8230 51408 8236
rect 51368 5302 51396 8230
rect 51724 7812 51776 7818
rect 51724 7754 51776 7760
rect 51632 5772 51684 5778
rect 51632 5714 51684 5720
rect 51356 5296 51408 5302
rect 51356 5238 51408 5244
rect 51448 5296 51500 5302
rect 51448 5238 51500 5244
rect 51356 4480 51408 4486
rect 51356 4422 51408 4428
rect 51368 4146 51396 4422
rect 51264 4140 51316 4146
rect 51264 4082 51316 4088
rect 51356 4140 51408 4146
rect 51356 4082 51408 4088
rect 51080 1352 51132 1358
rect 51080 1294 51132 1300
rect 50712 1216 50764 1222
rect 50712 1158 50764 1164
rect 51092 649 51120 1294
rect 51460 882 51488 5238
rect 51644 5166 51672 5714
rect 51632 5160 51684 5166
rect 51632 5102 51684 5108
rect 51540 4208 51592 4214
rect 51540 4150 51592 4156
rect 51552 1222 51580 4150
rect 51644 4078 51672 5102
rect 51736 4214 51764 7754
rect 52092 5296 52144 5302
rect 52092 5238 52144 5244
rect 51908 5024 51960 5030
rect 51908 4966 51960 4972
rect 52000 5024 52052 5030
rect 52000 4966 52052 4972
rect 51724 4208 51776 4214
rect 51724 4150 51776 4156
rect 51816 4208 51868 4214
rect 51816 4150 51868 4156
rect 51632 4072 51684 4078
rect 51630 4040 51632 4049
rect 51684 4040 51686 4049
rect 51630 3975 51686 3984
rect 51724 1352 51776 1358
rect 51724 1294 51776 1300
rect 51540 1216 51592 1222
rect 51540 1158 51592 1164
rect 51448 876 51500 882
rect 51448 818 51500 824
rect 51736 649 51764 1294
rect 43904 614 43956 620
rect 43994 640 44050 649
rect 43258 575 43314 584
rect 43994 575 44050 584
rect 44638 640 44694 649
rect 44638 575 44694 584
rect 45466 640 45522 649
rect 45466 575 45522 584
rect 45926 640 45982 649
rect 45926 575 45982 584
rect 46570 640 46626 649
rect 46570 575 46626 584
rect 47214 640 47270 649
rect 47214 575 47270 584
rect 48318 640 48374 649
rect 48318 575 48374 584
rect 49146 640 49202 649
rect 49146 575 49202 584
rect 49790 640 49846 649
rect 49790 575 49846 584
rect 50618 640 50674 649
rect 50618 575 50674 584
rect 51078 640 51134 649
rect 51078 575 51134 584
rect 51722 640 51778 649
rect 51722 575 51778 584
rect 51828 542 51856 4150
rect 51920 3534 51948 4966
rect 52012 4758 52040 4966
rect 52104 4826 52132 5238
rect 52092 4820 52144 4826
rect 52092 4762 52144 4768
rect 52000 4752 52052 4758
rect 52000 4694 52052 4700
rect 52288 4554 52316 9318
rect 53208 9178 53236 10231
rect 54680 9722 54708 10367
rect 57164 10334 57192 10406
rect 57152 10328 57204 10334
rect 54758 10296 54814 10305
rect 54758 10231 54814 10240
rect 55494 10296 55550 10305
rect 55494 10231 55550 10240
rect 56230 10296 56286 10305
rect 56230 10231 56286 10240
rect 57058 10296 57114 10305
rect 57152 10270 57204 10276
rect 57794 10296 57850 10305
rect 57058 10231 57114 10240
rect 54668 9716 54720 9722
rect 54668 9658 54720 9664
rect 54024 9580 54076 9586
rect 54024 9522 54076 9528
rect 54116 9580 54168 9586
rect 54116 9522 54168 9528
rect 53748 9444 53800 9450
rect 53748 9386 53800 9392
rect 53380 9376 53432 9382
rect 53380 9318 53432 9324
rect 53196 9172 53248 9178
rect 53196 9114 53248 9120
rect 53392 8974 53420 9318
rect 53380 8968 53432 8974
rect 53380 8910 53432 8916
rect 53472 8968 53524 8974
rect 53472 8910 53524 8916
rect 52828 7880 52880 7886
rect 52828 7822 52880 7828
rect 52840 4554 52868 7822
rect 53104 5772 53156 5778
rect 53104 5714 53156 5720
rect 53116 5370 53144 5714
rect 53104 5364 53156 5370
rect 53104 5306 53156 5312
rect 53116 4690 53144 5306
rect 53104 4684 53156 4690
rect 53104 4626 53156 4632
rect 52276 4548 52328 4554
rect 52276 4490 52328 4496
rect 52460 4548 52512 4554
rect 52460 4490 52512 4496
rect 52828 4548 52880 4554
rect 52828 4490 52880 4496
rect 52000 4480 52052 4486
rect 52000 4422 52052 4428
rect 51908 3528 51960 3534
rect 51908 3470 51960 3476
rect 52012 1222 52040 4422
rect 52472 4146 52500 4490
rect 53196 4480 53248 4486
rect 53196 4422 53248 4428
rect 53380 4480 53432 4486
rect 53380 4422 53432 4428
rect 52460 4140 52512 4146
rect 52460 4082 52512 4088
rect 52276 3936 52328 3942
rect 52276 3878 52328 3884
rect 52288 3194 52316 3878
rect 52276 3188 52328 3194
rect 52276 3130 52328 3136
rect 52920 1964 52972 1970
rect 52920 1906 52972 1912
rect 52368 1352 52420 1358
rect 52368 1294 52420 1300
rect 52000 1216 52052 1222
rect 52000 1158 52052 1164
rect 52380 649 52408 1294
rect 52932 1290 52960 1906
rect 52920 1284 52972 1290
rect 52920 1226 52972 1232
rect 53208 950 53236 4422
rect 53392 4282 53420 4422
rect 53380 4276 53432 4282
rect 53380 4218 53432 4224
rect 53484 2446 53512 8910
rect 53760 2514 53788 9386
rect 54036 8906 54064 9522
rect 54024 8900 54076 8906
rect 54024 8842 54076 8848
rect 54036 8498 54064 8842
rect 54128 8634 54156 9522
rect 54392 8968 54444 8974
rect 54392 8910 54444 8916
rect 54116 8628 54168 8634
rect 54116 8570 54168 8576
rect 54024 8492 54076 8498
rect 54024 8434 54076 8440
rect 54116 8424 54168 8430
rect 54116 8366 54168 8372
rect 54128 3058 54156 8366
rect 54404 3097 54432 8910
rect 54576 8832 54628 8838
rect 54576 8774 54628 8780
rect 54588 8498 54616 8774
rect 54772 8634 54800 10231
rect 55404 10056 55456 10062
rect 55404 9998 55456 10004
rect 55416 9110 55444 9998
rect 55404 9104 55456 9110
rect 55404 9046 55456 9052
rect 55416 8974 55444 9046
rect 55404 8968 55456 8974
rect 55404 8910 55456 8916
rect 55312 8832 55364 8838
rect 55312 8774 55364 8780
rect 54760 8628 54812 8634
rect 54760 8570 54812 8576
rect 55324 8498 55352 8774
rect 54576 8492 54628 8498
rect 54576 8434 54628 8440
rect 55312 8492 55364 8498
rect 55312 8434 55364 8440
rect 54390 3088 54446 3097
rect 54116 3052 54168 3058
rect 54390 3023 54446 3032
rect 54116 2994 54168 3000
rect 53748 2508 53800 2514
rect 53748 2450 53800 2456
rect 53472 2440 53524 2446
rect 53472 2382 53524 2388
rect 54024 2440 54076 2446
rect 54024 2382 54076 2388
rect 53484 1902 53512 2382
rect 53840 2304 53892 2310
rect 53840 2246 53892 2252
rect 53472 1896 53524 1902
rect 53472 1838 53524 1844
rect 53484 1766 53512 1838
rect 53472 1760 53524 1766
rect 53472 1702 53524 1708
rect 53484 1426 53512 1702
rect 53472 1420 53524 1426
rect 53472 1362 53524 1368
rect 53852 1358 53880 2246
rect 54036 1970 54064 2382
rect 54024 1964 54076 1970
rect 54024 1906 54076 1912
rect 53932 1828 53984 1834
rect 53932 1770 53984 1776
rect 53944 1465 53972 1770
rect 53930 1456 53986 1465
rect 53930 1391 53986 1400
rect 54036 1358 54064 1906
rect 54128 1494 54156 2994
rect 54208 2440 54260 2446
rect 54208 2382 54260 2388
rect 54220 2038 54248 2382
rect 54208 2032 54260 2038
rect 54404 2009 54432 3023
rect 55036 2440 55088 2446
rect 55036 2382 55088 2388
rect 54852 2304 54904 2310
rect 54852 2246 54904 2252
rect 54208 1974 54260 1980
rect 54390 2000 54446 2009
rect 54390 1935 54446 1944
rect 54404 1902 54432 1935
rect 54392 1896 54444 1902
rect 54392 1838 54444 1844
rect 54116 1488 54168 1494
rect 54206 1456 54262 1465
rect 54168 1436 54206 1442
rect 54116 1430 54206 1436
rect 54128 1414 54206 1430
rect 54206 1391 54262 1400
rect 53840 1352 53892 1358
rect 53840 1294 53892 1300
rect 54024 1352 54076 1358
rect 54024 1294 54076 1300
rect 53380 1216 53432 1222
rect 53380 1158 53432 1164
rect 53196 944 53248 950
rect 53196 886 53248 892
rect 53392 649 53420 1158
rect 54864 649 54892 2246
rect 55048 2038 55076 2382
rect 55036 2032 55088 2038
rect 55036 1974 55088 1980
rect 55416 1970 55444 8910
rect 55508 8634 55536 10231
rect 55864 9512 55916 9518
rect 55864 9454 55916 9460
rect 55876 9042 55904 9454
rect 55864 9036 55916 9042
rect 55864 8978 55916 8984
rect 56048 8832 56100 8838
rect 56048 8774 56100 8780
rect 55496 8628 55548 8634
rect 55496 8570 55548 8576
rect 56060 8498 56088 8774
rect 56244 8634 56272 10231
rect 56416 10124 56468 10130
rect 56416 10066 56468 10072
rect 56428 9178 56456 10066
rect 56416 9172 56468 9178
rect 56416 9114 56468 9120
rect 56428 8974 56456 9114
rect 56416 8968 56468 8974
rect 56416 8910 56468 8916
rect 56232 8628 56284 8634
rect 56232 8570 56284 8576
rect 56048 8492 56100 8498
rect 56048 8434 56100 8440
rect 56428 2774 56456 8910
rect 56876 8832 56928 8838
rect 56876 8774 56928 8780
rect 56888 8498 56916 8774
rect 57072 8634 57100 10231
rect 57164 8974 57192 10270
rect 57794 10231 57850 10240
rect 58622 10296 58678 10305
rect 58622 10231 58678 10240
rect 59266 10296 59322 10305
rect 60002 10296 60058 10305
rect 59266 10231 59322 10240
rect 59636 10260 59688 10266
rect 57808 9722 57836 10231
rect 57796 9716 57848 9722
rect 57796 9658 57848 9664
rect 57520 9580 57572 9586
rect 57520 9522 57572 9528
rect 57532 9178 57560 9522
rect 57520 9172 57572 9178
rect 57520 9114 57572 9120
rect 57152 8968 57204 8974
rect 57152 8910 57204 8916
rect 57060 8628 57112 8634
rect 57060 8570 57112 8576
rect 56876 8492 56928 8498
rect 56876 8434 56928 8440
rect 56336 2746 56456 2774
rect 55680 2304 55732 2310
rect 55680 2246 55732 2252
rect 55404 1964 55456 1970
rect 55404 1906 55456 1912
rect 55692 649 55720 2246
rect 56336 1970 56364 2746
rect 57164 1970 57192 8910
rect 58532 8900 58584 8906
rect 58532 8842 58584 8848
rect 58440 8832 58492 8838
rect 58440 8774 58492 8780
rect 58452 8498 58480 8774
rect 58440 8492 58492 8498
rect 58440 8434 58492 8440
rect 57520 2440 57572 2446
rect 57520 2382 57572 2388
rect 57532 2106 57560 2382
rect 57796 2304 57848 2310
rect 57796 2246 57848 2252
rect 57520 2100 57572 2106
rect 57520 2042 57572 2048
rect 56324 1964 56376 1970
rect 56324 1906 56376 1912
rect 57152 1964 57204 1970
rect 57152 1906 57204 1912
rect 56048 1760 56100 1766
rect 56048 1702 56100 1708
rect 56876 1760 56928 1766
rect 56876 1702 56928 1708
rect 56060 1358 56088 1702
rect 56888 1358 56916 1702
rect 56048 1352 56100 1358
rect 56048 1294 56100 1300
rect 56876 1352 56928 1358
rect 56876 1294 56928 1300
rect 56232 1216 56284 1222
rect 56232 1158 56284 1164
rect 57060 1216 57112 1222
rect 57060 1158 57112 1164
rect 56244 649 56272 1158
rect 57072 649 57100 1158
rect 57808 649 57836 2246
rect 58544 2106 58572 8842
rect 58636 8634 58664 10231
rect 58900 9920 58952 9926
rect 58900 9862 58952 9868
rect 58912 8974 58940 9862
rect 59280 9722 59308 10231
rect 60002 10231 60058 10240
rect 59636 10202 59688 10208
rect 59268 9716 59320 9722
rect 59268 9658 59320 9664
rect 59176 9580 59228 9586
rect 59176 9522 59228 9528
rect 59188 9178 59216 9522
rect 59648 9382 59676 10202
rect 60016 9722 60044 10231
rect 60004 9716 60056 9722
rect 60004 9658 60056 9664
rect 60108 9654 60136 10474
rect 60096 9648 60148 9654
rect 60096 9590 60148 9596
rect 60004 9580 60056 9586
rect 60004 9522 60056 9528
rect 59636 9376 59688 9382
rect 59636 9318 59688 9324
rect 59176 9172 59228 9178
rect 59176 9114 59228 9120
rect 59648 8974 59676 9318
rect 60016 9178 60044 9522
rect 60004 9172 60056 9178
rect 60004 9114 60056 9120
rect 60108 8974 60136 9590
rect 58900 8968 58952 8974
rect 58900 8910 58952 8916
rect 59636 8968 59688 8974
rect 59636 8910 59688 8916
rect 59820 8968 59872 8974
rect 59820 8910 59872 8916
rect 60096 8968 60148 8974
rect 60096 8910 60148 8916
rect 58624 8628 58676 8634
rect 58624 8570 58676 8576
rect 58912 2650 58940 8910
rect 59648 2774 59676 8910
rect 59832 8634 59860 8910
rect 59820 8628 59872 8634
rect 59820 8570 59872 8576
rect 60384 8430 60412 10542
rect 62396 10396 62448 10402
rect 62396 10338 62448 10344
rect 61476 10328 61528 10334
rect 60830 10296 60886 10305
rect 61476 10270 61528 10276
rect 61566 10296 61622 10305
rect 60830 10231 60886 10240
rect 60844 9722 60872 10231
rect 60832 9716 60884 9722
rect 60832 9658 60884 9664
rect 60740 9580 60792 9586
rect 60740 9522 60792 9528
rect 60648 8968 60700 8974
rect 60648 8910 60700 8916
rect 60372 8424 60424 8430
rect 60372 8366 60424 8372
rect 60384 7478 60412 8366
rect 59820 7472 59872 7478
rect 59820 7414 59872 7420
rect 60372 7472 60424 7478
rect 60372 7414 60424 7420
rect 59648 2746 59768 2774
rect 58900 2644 58952 2650
rect 58900 2586 58952 2592
rect 58532 2100 58584 2106
rect 58532 2042 58584 2048
rect 58544 1902 58572 2042
rect 58912 1902 58940 2586
rect 59268 2440 59320 2446
rect 59268 2382 59320 2388
rect 59280 2106 59308 2382
rect 59360 2304 59412 2310
rect 59360 2246 59412 2252
rect 59268 2100 59320 2106
rect 59268 2042 59320 2048
rect 58532 1896 58584 1902
rect 58532 1838 58584 1844
rect 58900 1896 58952 1902
rect 58900 1838 58952 1844
rect 58440 1760 58492 1766
rect 58440 1702 58492 1708
rect 58452 1358 58480 1702
rect 58912 1562 58940 1838
rect 59372 1601 59400 2246
rect 59358 1592 59414 1601
rect 58900 1556 58952 1562
rect 59358 1527 59414 1536
rect 58900 1498 58952 1504
rect 59740 1358 59768 2746
rect 59832 1970 59860 7414
rect 60004 2440 60056 2446
rect 60004 2382 60056 2388
rect 59820 1964 59872 1970
rect 59820 1906 59872 1912
rect 59912 1896 59964 1902
rect 59912 1838 59964 1844
rect 59924 1358 59952 1838
rect 60016 1562 60044 2382
rect 60660 1970 60688 8910
rect 60752 8634 60780 9522
rect 61488 9518 61516 10270
rect 61566 10231 61622 10240
rect 62302 10296 62358 10305
rect 62302 10231 62358 10240
rect 61476 9512 61528 9518
rect 61476 9454 61528 9460
rect 61488 8974 61516 9454
rect 60924 8968 60976 8974
rect 60924 8910 60976 8916
rect 61476 8968 61528 8974
rect 61476 8910 61528 8916
rect 60740 8628 60792 8634
rect 60740 8570 60792 8576
rect 60936 8498 60964 8910
rect 61384 8832 61436 8838
rect 61384 8774 61436 8780
rect 61396 8498 61424 8774
rect 60924 8492 60976 8498
rect 60924 8434 60976 8440
rect 61384 8492 61436 8498
rect 61384 8434 61436 8440
rect 61488 6914 61516 8910
rect 61580 8634 61608 10231
rect 62120 8832 62172 8838
rect 62120 8774 62172 8780
rect 61568 8628 61620 8634
rect 61568 8570 61620 8576
rect 62132 8498 62160 8774
rect 62316 8634 62344 10231
rect 62408 8974 62436 10338
rect 62764 9580 62816 9586
rect 62764 9522 62816 9528
rect 62776 9178 62804 9522
rect 62764 9172 62816 9178
rect 62764 9114 62816 9120
rect 63236 8974 63264 10610
rect 63406 10296 63462 10305
rect 63406 10231 63462 10240
rect 63774 10296 63830 10305
rect 63774 10231 63830 10240
rect 64602 10296 64658 10305
rect 64602 10231 64658 10240
rect 65430 10296 65486 10305
rect 65430 10231 65486 10240
rect 63420 9722 63448 10231
rect 63408 9716 63460 9722
rect 63408 9658 63460 9664
rect 62396 8968 62448 8974
rect 62396 8910 62448 8916
rect 63224 8968 63276 8974
rect 63224 8910 63276 8916
rect 62304 8628 62356 8634
rect 62304 8570 62356 8576
rect 62120 8492 62172 8498
rect 62120 8434 62172 8440
rect 61488 6886 61608 6914
rect 60738 4312 60794 4321
rect 60738 4247 60794 4256
rect 60752 3670 60780 4247
rect 60740 3664 60792 3670
rect 60740 3606 60792 3612
rect 60738 2816 60794 2825
rect 60738 2751 60794 2760
rect 60752 2650 60780 2751
rect 60740 2644 60792 2650
rect 60740 2586 60792 2592
rect 61580 1970 61608 6886
rect 62408 1970 62436 8910
rect 62672 2440 62724 2446
rect 62672 2382 62724 2388
rect 62684 2106 62712 2382
rect 62948 2304 63000 2310
rect 62948 2246 63000 2252
rect 62672 2100 62724 2106
rect 62672 2042 62724 2048
rect 60648 1964 60700 1970
rect 60648 1906 60700 1912
rect 61568 1964 61620 1970
rect 61568 1906 61620 1912
rect 62396 1964 62448 1970
rect 62396 1906 62448 1912
rect 60648 1760 60700 1766
rect 60648 1702 60700 1708
rect 61384 1760 61436 1766
rect 61384 1702 61436 1708
rect 61844 1760 61896 1766
rect 61844 1702 61896 1708
rect 60004 1556 60056 1562
rect 60004 1498 60056 1504
rect 60660 1358 60688 1702
rect 61396 1358 61424 1702
rect 61856 1358 61884 1702
rect 58440 1352 58492 1358
rect 58440 1294 58492 1300
rect 59728 1352 59780 1358
rect 59728 1294 59780 1300
rect 59912 1352 59964 1358
rect 59912 1294 59964 1300
rect 60648 1352 60700 1358
rect 60648 1294 60700 1300
rect 61384 1352 61436 1358
rect 61384 1294 61436 1300
rect 61844 1352 61896 1358
rect 61844 1294 61896 1300
rect 58624 1216 58676 1222
rect 58624 1158 58676 1164
rect 60832 1216 60884 1222
rect 60832 1158 60884 1164
rect 61568 1216 61620 1222
rect 61568 1158 61620 1164
rect 62304 1216 62356 1222
rect 62304 1158 62356 1164
rect 58636 649 58664 1158
rect 60844 649 60872 1158
rect 61580 649 61608 1158
rect 62316 649 62344 1158
rect 62960 649 62988 2246
rect 63236 1970 63264 8910
rect 63592 8832 63644 8838
rect 63592 8774 63644 8780
rect 63604 8498 63632 8774
rect 63788 8634 63816 10231
rect 64052 10192 64104 10198
rect 64052 10134 64104 10140
rect 64064 9178 64092 10134
rect 64052 9172 64104 9178
rect 64052 9114 64104 9120
rect 64064 8974 64092 9114
rect 64052 8968 64104 8974
rect 64052 8910 64104 8916
rect 63776 8628 63828 8634
rect 63776 8570 63828 8576
rect 63592 8492 63644 8498
rect 63592 8434 63644 8440
rect 64064 1970 64092 8910
rect 64420 8832 64472 8838
rect 64420 8774 64472 8780
rect 64432 8498 64460 8774
rect 64616 8634 64644 10231
rect 64972 9988 65024 9994
rect 64972 9930 65024 9936
rect 64696 9104 64748 9110
rect 64696 9046 64748 9052
rect 64708 8634 64736 9046
rect 64984 8974 65012 9930
rect 64972 8968 65024 8974
rect 64972 8910 65024 8916
rect 64604 8628 64656 8634
rect 64604 8570 64656 8576
rect 64696 8628 64748 8634
rect 64696 8570 64748 8576
rect 64420 8492 64472 8498
rect 64420 8434 64472 8440
rect 64984 6914 65012 8910
rect 65248 8832 65300 8838
rect 65248 8774 65300 8780
rect 65260 8498 65288 8774
rect 65248 8492 65300 8498
rect 65248 8434 65300 8440
rect 65444 8362 65472 10231
rect 65996 8974 66024 10678
rect 75000 10668 75052 10674
rect 75000 10610 75052 10616
rect 71318 10568 71374 10577
rect 71318 10503 71374 10512
rect 74262 10568 74318 10577
rect 74262 10503 74318 10512
rect 66166 10296 66222 10305
rect 66076 10260 66128 10266
rect 66166 10231 66222 10240
rect 66902 10296 66958 10305
rect 66902 10231 66958 10240
rect 66076 10202 66128 10208
rect 66088 9994 66116 10202
rect 66076 9988 66128 9994
rect 66076 9930 66128 9936
rect 66180 9722 66208 10231
rect 66916 9722 66944 10231
rect 68546 9820 68854 9829
rect 68546 9818 68552 9820
rect 68608 9818 68632 9820
rect 68688 9818 68712 9820
rect 68768 9818 68792 9820
rect 68848 9818 68854 9820
rect 68608 9766 68610 9818
rect 68790 9766 68792 9818
rect 68546 9764 68552 9766
rect 68608 9764 68632 9766
rect 68688 9764 68712 9766
rect 68768 9764 68792 9766
rect 68848 9764 68854 9766
rect 68546 9755 68854 9764
rect 66168 9716 66220 9722
rect 66168 9658 66220 9664
rect 66904 9716 66956 9722
rect 66904 9658 66956 9664
rect 69110 9616 69166 9625
rect 66352 9580 66404 9586
rect 66352 9522 66404 9528
rect 66996 9580 67048 9586
rect 69110 9551 69112 9560
rect 66996 9522 67048 9528
rect 69164 9551 69166 9560
rect 70306 9616 70362 9625
rect 70306 9551 70308 9560
rect 69112 9522 69164 9528
rect 70360 9551 70362 9560
rect 70308 9522 70360 9528
rect 66364 9178 66392 9522
rect 66352 9172 66404 9178
rect 66352 9114 66404 9120
rect 65984 8968 66036 8974
rect 65984 8910 66036 8916
rect 66904 8968 66956 8974
rect 66904 8910 66956 8916
rect 65996 8566 66024 8910
rect 66812 8832 66864 8838
rect 66812 8774 66864 8780
rect 65708 8560 65760 8566
rect 65708 8502 65760 8508
rect 65984 8560 66036 8566
rect 65984 8502 66036 8508
rect 65432 8356 65484 8362
rect 65432 8298 65484 8304
rect 64892 6886 65012 6914
rect 63224 1964 63276 1970
rect 63224 1906 63276 1912
rect 64052 1964 64104 1970
rect 64052 1906 64104 1912
rect 64892 1902 64920 6886
rect 65248 2440 65300 2446
rect 65248 2382 65300 2388
rect 65260 2106 65288 2382
rect 65616 2304 65668 2310
rect 65616 2246 65668 2252
rect 65248 2100 65300 2106
rect 65248 2042 65300 2048
rect 64880 1896 64932 1902
rect 64880 1838 64932 1844
rect 63592 1760 63644 1766
rect 63592 1702 63644 1708
rect 64328 1760 64380 1766
rect 64328 1702 64380 1708
rect 63604 1358 63632 1702
rect 64340 1358 64368 1702
rect 63592 1352 63644 1358
rect 63592 1294 63644 1300
rect 64328 1352 64380 1358
rect 64328 1294 64380 1300
rect 63776 1216 63828 1222
rect 63776 1158 63828 1164
rect 64512 1216 64564 1222
rect 64512 1158 64564 1164
rect 63788 649 63816 1158
rect 64524 649 64552 1158
rect 65628 649 65656 2246
rect 65720 1970 65748 8502
rect 66824 8498 66852 8774
rect 66812 8492 66864 8498
rect 66812 8434 66864 8440
rect 66916 8362 66944 8910
rect 67008 8566 67036 9522
rect 67272 9172 67324 9178
rect 67272 9114 67324 9120
rect 67180 9036 67232 9042
rect 67284 9024 67312 9114
rect 67232 8996 67312 9024
rect 69570 9072 69626 9081
rect 69570 9007 69572 9016
rect 67180 8978 67232 8984
rect 69624 9007 69626 9016
rect 69572 8978 69624 8984
rect 69848 8968 69900 8974
rect 69848 8910 69900 8916
rect 68546 8732 68854 8741
rect 68546 8730 68552 8732
rect 68608 8730 68632 8732
rect 68688 8730 68712 8732
rect 68768 8730 68792 8732
rect 68848 8730 68854 8732
rect 68608 8678 68610 8730
rect 68790 8678 68792 8730
rect 68546 8676 68552 8678
rect 68608 8676 68632 8678
rect 68688 8676 68712 8678
rect 68768 8676 68792 8678
rect 68848 8676 68854 8678
rect 68546 8667 68854 8676
rect 66996 8560 67048 8566
rect 66996 8502 67048 8508
rect 66904 8356 66956 8362
rect 66904 8298 66956 8304
rect 66916 7546 66944 8298
rect 69860 7818 69888 8910
rect 71332 8498 71360 10503
rect 72054 10432 72110 10441
rect 72054 10367 72110 10376
rect 72068 9042 72096 10367
rect 72146 9616 72202 9625
rect 72146 9551 72148 9560
rect 72200 9551 72202 9560
rect 72148 9522 72200 9528
rect 72424 9376 72476 9382
rect 72424 9318 72476 9324
rect 72056 9036 72108 9042
rect 72056 8978 72108 8984
rect 72436 8906 72464 9318
rect 73434 9072 73490 9081
rect 73434 9007 73436 9016
rect 73488 9007 73490 9016
rect 73436 8978 73488 8984
rect 73712 8968 73764 8974
rect 73712 8910 73764 8916
rect 72424 8900 72476 8906
rect 72424 8842 72476 8848
rect 71320 8492 71372 8498
rect 71320 8434 71372 8440
rect 71596 8424 71648 8430
rect 71596 8366 71648 8372
rect 69848 7812 69900 7818
rect 69848 7754 69900 7760
rect 68546 7644 68854 7653
rect 68546 7642 68552 7644
rect 68608 7642 68632 7644
rect 68688 7642 68712 7644
rect 68768 7642 68792 7644
rect 68848 7642 68854 7644
rect 68608 7590 68610 7642
rect 68790 7590 68792 7642
rect 68546 7588 68552 7590
rect 68608 7588 68632 7590
rect 68688 7588 68712 7590
rect 68768 7588 68792 7590
rect 68848 7588 68854 7590
rect 68546 7579 68854 7588
rect 66904 7540 66956 7546
rect 66904 7482 66956 7488
rect 68546 6556 68854 6565
rect 68546 6554 68552 6556
rect 68608 6554 68632 6556
rect 68688 6554 68712 6556
rect 68768 6554 68792 6556
rect 68848 6554 68854 6556
rect 68608 6502 68610 6554
rect 68790 6502 68792 6554
rect 68546 6500 68552 6502
rect 68608 6500 68632 6502
rect 68688 6500 68712 6502
rect 68768 6500 68792 6502
rect 68848 6500 68854 6502
rect 68546 6491 68854 6500
rect 71608 6254 71636 8366
rect 73724 8022 73752 8910
rect 74276 8498 74304 10503
rect 74722 9616 74778 9625
rect 74722 9551 74724 9560
rect 74776 9551 74778 9560
rect 74724 9522 74776 9528
rect 74722 9072 74778 9081
rect 75012 9042 75040 10610
rect 84566 10568 84622 10577
rect 84566 10503 84622 10512
rect 86774 10568 86830 10577
rect 90836 10538 90864 10746
rect 94964 10600 95016 10606
rect 94964 10542 95016 10548
rect 86774 10503 86830 10512
rect 90824 10532 90876 10538
rect 77206 10432 77262 10441
rect 77206 10367 77262 10376
rect 82358 10432 82414 10441
rect 82358 10367 82414 10376
rect 83830 10432 83886 10441
rect 83830 10367 83886 10376
rect 76748 9988 76800 9994
rect 76748 9930 76800 9936
rect 76470 9752 76526 9761
rect 76470 9687 76526 9696
rect 75828 9512 75880 9518
rect 75828 9454 75880 9460
rect 74722 9007 74724 9016
rect 74776 9007 74778 9016
rect 75000 9036 75052 9042
rect 74724 8978 74776 8984
rect 75000 8978 75052 8984
rect 74264 8492 74316 8498
rect 74264 8434 74316 8440
rect 74540 8424 74592 8430
rect 74540 8366 74592 8372
rect 73712 8016 73764 8022
rect 73712 7958 73764 7964
rect 72332 6452 72384 6458
rect 72332 6394 72384 6400
rect 71596 6248 71648 6254
rect 71596 6190 71648 6196
rect 68546 5468 68854 5477
rect 68546 5466 68552 5468
rect 68608 5466 68632 5468
rect 68688 5466 68712 5468
rect 68768 5466 68792 5468
rect 68848 5466 68854 5468
rect 68608 5414 68610 5466
rect 68790 5414 68792 5466
rect 68546 5412 68552 5414
rect 68608 5412 68632 5414
rect 68688 5412 68712 5414
rect 68768 5412 68792 5414
rect 68848 5412 68854 5414
rect 68546 5403 68854 5412
rect 67546 5264 67602 5273
rect 67546 5199 67602 5208
rect 66720 3732 66772 3738
rect 66720 3674 66772 3680
rect 66628 2304 66680 2310
rect 66628 2246 66680 2252
rect 66640 1970 66668 2246
rect 66732 1970 66760 3674
rect 66996 3528 67048 3534
rect 67180 3528 67232 3534
rect 67048 3476 67180 3482
rect 66996 3470 67232 3476
rect 67008 3454 67220 3470
rect 67560 2990 67588 5199
rect 68546 4380 68854 4389
rect 68546 4378 68552 4380
rect 68608 4378 68632 4380
rect 68688 4378 68712 4380
rect 68768 4378 68792 4380
rect 68848 4378 68854 4380
rect 68608 4326 68610 4378
rect 68790 4326 68792 4378
rect 68546 4324 68552 4326
rect 68608 4324 68632 4326
rect 68688 4324 68712 4326
rect 68768 4324 68792 4326
rect 68848 4324 68854 4326
rect 68546 4315 68854 4324
rect 68546 3292 68854 3301
rect 68546 3290 68552 3292
rect 68608 3290 68632 3292
rect 68688 3290 68712 3292
rect 68768 3290 68792 3292
rect 68848 3290 68854 3292
rect 68608 3238 68610 3290
rect 68790 3238 68792 3290
rect 68546 3236 68552 3238
rect 68608 3236 68632 3238
rect 68688 3236 68712 3238
rect 68768 3236 68792 3238
rect 68848 3236 68854 3238
rect 68546 3227 68854 3236
rect 67548 2984 67600 2990
rect 67548 2926 67600 2932
rect 70860 2576 70912 2582
rect 70860 2518 70912 2524
rect 68546 2204 68854 2213
rect 68546 2202 68552 2204
rect 68608 2202 68632 2204
rect 68688 2202 68712 2204
rect 68768 2202 68792 2204
rect 68848 2202 68854 2204
rect 68608 2150 68610 2202
rect 68790 2150 68792 2202
rect 68546 2148 68552 2150
rect 68608 2148 68632 2150
rect 68688 2148 68712 2150
rect 68768 2148 68792 2150
rect 68848 2148 68854 2150
rect 68546 2139 68854 2148
rect 70872 1970 70900 2518
rect 71320 2440 71372 2446
rect 71320 2382 71372 2388
rect 65708 1964 65760 1970
rect 65708 1906 65760 1912
rect 66628 1964 66680 1970
rect 66628 1906 66680 1912
rect 66720 1964 66772 1970
rect 66720 1906 66772 1912
rect 70860 1964 70912 1970
rect 70860 1906 70912 1912
rect 70584 1896 70636 1902
rect 70584 1838 70636 1844
rect 65984 1760 66036 1766
rect 65984 1702 66036 1708
rect 67548 1760 67600 1766
rect 67548 1702 67600 1708
rect 65996 1358 66024 1702
rect 65984 1352 66036 1358
rect 65984 1294 66036 1300
rect 66168 1216 66220 1222
rect 66168 1158 66220 1164
rect 52366 640 52422 649
rect 52366 575 52422 584
rect 53378 640 53434 649
rect 53378 575 53434 584
rect 54850 640 54906 649
rect 54850 575 54906 584
rect 55678 640 55734 649
rect 55678 575 55734 584
rect 56230 640 56286 649
rect 56230 575 56286 584
rect 57058 640 57114 649
rect 57058 575 57114 584
rect 57794 640 57850 649
rect 57794 575 57850 584
rect 58622 640 58678 649
rect 58622 575 58678 584
rect 60830 640 60886 649
rect 60830 575 60886 584
rect 61566 640 61622 649
rect 61566 575 61622 584
rect 62302 640 62358 649
rect 62302 575 62358 584
rect 62946 640 63002 649
rect 62946 575 63002 584
rect 63774 640 63830 649
rect 63774 575 63830 584
rect 64510 640 64566 649
rect 64510 575 64566 584
rect 65614 640 65670 649
rect 65614 575 65670 584
rect 51816 536 51868 542
rect 66180 513 66208 1158
rect 67560 513 67588 1702
rect 69112 1420 69164 1426
rect 69112 1362 69164 1368
rect 68546 1116 68854 1125
rect 68546 1114 68552 1116
rect 68608 1114 68632 1116
rect 68688 1114 68712 1116
rect 68768 1114 68792 1116
rect 68848 1114 68854 1116
rect 68608 1062 68610 1114
rect 68790 1062 68792 1114
rect 68546 1060 68552 1062
rect 68608 1060 68632 1062
rect 68688 1060 68712 1062
rect 68768 1060 68792 1062
rect 68848 1060 68854 1062
rect 68546 1051 68854 1060
rect 69124 785 69152 1362
rect 69572 1352 69624 1358
rect 69572 1294 69624 1300
rect 69848 1352 69900 1358
rect 69848 1294 69900 1300
rect 69584 785 69612 1294
rect 69860 1018 69888 1294
rect 70596 1057 70624 1838
rect 71332 1329 71360 2382
rect 72344 1970 72372 6394
rect 74552 4826 74580 8366
rect 75840 6866 75868 9454
rect 76484 8498 76512 9687
rect 76760 8498 76788 9930
rect 77220 9042 77248 10367
rect 77484 10192 77536 10198
rect 77484 10134 77536 10140
rect 77298 9616 77354 9625
rect 77298 9551 77300 9560
rect 77352 9551 77354 9560
rect 77300 9522 77352 9528
rect 77496 9042 77524 10134
rect 79414 9752 79470 9761
rect 79414 9687 79470 9696
rect 81622 9752 81678 9761
rect 81622 9687 81678 9696
rect 77576 9512 77628 9518
rect 77576 9454 77628 9460
rect 77208 9036 77260 9042
rect 77208 8978 77260 8984
rect 77484 9036 77536 9042
rect 77484 8978 77536 8984
rect 76472 8492 76524 8498
rect 76472 8434 76524 8440
rect 76748 8492 76800 8498
rect 76748 8434 76800 8440
rect 77588 7478 77616 9454
rect 78586 9072 78642 9081
rect 78586 9007 78588 9016
rect 78640 9007 78642 9016
rect 78588 8978 78640 8984
rect 78864 8968 78916 8974
rect 78864 8910 78916 8916
rect 78220 7540 78272 7546
rect 78220 7482 78272 7488
rect 77576 7472 77628 7478
rect 77576 7414 77628 7420
rect 75828 6860 75880 6866
rect 75828 6802 75880 6808
rect 77300 5840 77352 5846
rect 77300 5782 77352 5788
rect 74540 4820 74592 4826
rect 74540 4762 74592 4768
rect 77312 3602 77340 5782
rect 78128 5024 78180 5030
rect 78128 4966 78180 4972
rect 78140 4690 78168 4966
rect 78128 4684 78180 4690
rect 78128 4626 78180 4632
rect 77300 3596 77352 3602
rect 77300 3538 77352 3544
rect 73160 2916 73212 2922
rect 73160 2858 73212 2864
rect 73172 2446 73200 2858
rect 78232 2514 78260 7482
rect 78876 7274 78904 8910
rect 79428 8498 79456 9687
rect 79966 9616 80022 9625
rect 79966 9551 79968 9560
rect 80020 9551 80022 9560
rect 79968 9522 80020 9528
rect 81348 9512 81400 9518
rect 81348 9454 81400 9460
rect 79966 9072 80022 9081
rect 79966 9007 79968 9016
rect 80020 9007 80022 9016
rect 79968 8978 80020 8984
rect 80152 8968 80204 8974
rect 80152 8910 80204 8916
rect 79416 8492 79468 8498
rect 79416 8434 79468 8440
rect 79416 7404 79468 7410
rect 79416 7346 79468 7352
rect 78864 7268 78916 7274
rect 78864 7210 78916 7216
rect 79428 7002 79456 7346
rect 80164 7342 80192 8910
rect 80152 7336 80204 7342
rect 80152 7278 80204 7284
rect 79600 7200 79652 7206
rect 79600 7142 79652 7148
rect 80152 7200 80204 7206
rect 80152 7142 80204 7148
rect 79048 6996 79100 7002
rect 79048 6938 79100 6944
rect 79416 6996 79468 7002
rect 79416 6938 79468 6944
rect 79060 6186 79088 6938
rect 79322 6760 79378 6769
rect 79152 6730 79322 6746
rect 79140 6724 79322 6730
rect 79192 6718 79322 6724
rect 79322 6695 79378 6704
rect 79140 6666 79192 6672
rect 79336 6390 79364 6695
rect 79416 6656 79468 6662
rect 79416 6598 79468 6604
rect 79324 6384 79376 6390
rect 79324 6326 79376 6332
rect 79048 6180 79100 6186
rect 79048 6122 79100 6128
rect 79060 5914 79088 6122
rect 79048 5908 79100 5914
rect 79048 5850 79100 5856
rect 79336 5778 79364 6326
rect 79428 6118 79456 6598
rect 79612 6458 79640 7142
rect 79692 6860 79744 6866
rect 79692 6802 79744 6808
rect 79600 6452 79652 6458
rect 79600 6394 79652 6400
rect 79704 6186 79732 6802
rect 80060 6656 80112 6662
rect 80060 6598 80112 6604
rect 79692 6180 79744 6186
rect 79692 6122 79744 6128
rect 79416 6112 79468 6118
rect 79416 6054 79468 6060
rect 79324 5772 79376 5778
rect 79324 5714 79376 5720
rect 79428 5574 79456 6054
rect 79416 5568 79468 5574
rect 80072 5522 80100 6598
rect 79416 5510 79468 5516
rect 79980 5494 80100 5522
rect 79232 3732 79284 3738
rect 79232 3674 79284 3680
rect 79244 3466 79272 3674
rect 79232 3460 79284 3466
rect 79232 3402 79284 3408
rect 78220 2508 78272 2514
rect 78220 2450 78272 2456
rect 79980 2446 80008 5494
rect 73160 2440 73212 2446
rect 73160 2382 73212 2388
rect 73528 2440 73580 2446
rect 73528 2382 73580 2388
rect 73804 2440 73856 2446
rect 73804 2382 73856 2388
rect 76472 2440 76524 2446
rect 76472 2382 76524 2388
rect 76748 2440 76800 2446
rect 76748 2382 76800 2388
rect 77944 2440 77996 2446
rect 77944 2382 77996 2388
rect 79416 2440 79468 2446
rect 79416 2382 79468 2388
rect 79968 2440 80020 2446
rect 79968 2382 80020 2388
rect 72332 1964 72384 1970
rect 72332 1906 72384 1912
rect 72056 1896 72108 1902
rect 72056 1838 72108 1844
rect 71318 1320 71374 1329
rect 71318 1255 71374 1264
rect 72068 1057 72096 1838
rect 72148 1352 72200 1358
rect 72148 1294 72200 1300
rect 72424 1352 72476 1358
rect 73540 1329 73568 2382
rect 72424 1294 72476 1300
rect 73526 1320 73582 1329
rect 70582 1048 70638 1057
rect 69848 1012 69900 1018
rect 70582 983 70638 992
rect 72054 1048 72110 1057
rect 72054 983 72110 992
rect 69848 954 69900 960
rect 69110 776 69166 785
rect 69110 711 69166 720
rect 69570 776 69626 785
rect 69570 711 69626 720
rect 72160 649 72188 1294
rect 72146 640 72202 649
rect 72146 575 72202 584
rect 51816 478 51868 484
rect 66166 504 66222 513
rect 66166 439 66222 448
rect 67546 504 67602 513
rect 72436 474 72464 1294
rect 73526 1255 73582 1264
rect 73816 678 73844 2382
rect 74264 1896 74316 1902
rect 74264 1838 74316 1844
rect 75736 1896 75788 1902
rect 75736 1838 75788 1844
rect 74276 1057 74304 1838
rect 74724 1352 74776 1358
rect 74724 1294 74776 1300
rect 75000 1352 75052 1358
rect 75000 1294 75052 1300
rect 74262 1048 74318 1057
rect 74262 983 74318 992
rect 73804 672 73856 678
rect 74736 649 74764 1294
rect 73804 614 73856 620
rect 74722 640 74778 649
rect 75012 610 75040 1294
rect 75748 1057 75776 1838
rect 76484 1329 76512 2382
rect 76470 1320 76526 1329
rect 76470 1255 76526 1264
rect 75734 1048 75790 1057
rect 75734 983 75790 992
rect 76760 746 76788 2382
rect 77208 1896 77260 1902
rect 77208 1838 77260 1844
rect 77220 1057 77248 1838
rect 77576 1352 77628 1358
rect 77956 1329 77984 2382
rect 79428 1329 79456 2382
rect 80164 1970 80192 7142
rect 81360 6390 81388 9454
rect 81636 8498 81664 9687
rect 82372 9042 82400 10367
rect 82634 9616 82690 9625
rect 82634 9551 82636 9560
rect 82688 9551 82690 9560
rect 82636 9522 82688 9528
rect 82728 9512 82780 9518
rect 82728 9454 82780 9460
rect 82360 9036 82412 9042
rect 82360 8978 82412 8984
rect 82636 8968 82688 8974
rect 82636 8910 82688 8916
rect 81624 8492 81676 8498
rect 81624 8434 81676 8440
rect 81900 8424 81952 8430
rect 81900 8366 81952 8372
rect 81912 7954 81940 8366
rect 82176 8016 82228 8022
rect 82176 7958 82228 7964
rect 81900 7948 81952 7954
rect 81900 7890 81952 7896
rect 81348 6384 81400 6390
rect 81348 6326 81400 6332
rect 81990 5808 82046 5817
rect 80796 5772 80848 5778
rect 81990 5743 81992 5752
rect 80796 5714 80848 5720
rect 82044 5743 82046 5752
rect 81992 5714 82044 5720
rect 80336 5296 80388 5302
rect 80334 5264 80336 5273
rect 80388 5264 80390 5273
rect 80808 5234 80836 5714
rect 81440 5704 81492 5710
rect 81440 5646 81492 5652
rect 81898 5672 81954 5681
rect 81348 5296 81400 5302
rect 80886 5264 80942 5273
rect 80334 5199 80390 5208
rect 80796 5228 80848 5234
rect 81452 5250 81480 5646
rect 81898 5607 81954 5616
rect 81400 5244 81480 5250
rect 81348 5238 81480 5244
rect 81624 5296 81676 5302
rect 81624 5238 81676 5244
rect 81360 5222 81480 5238
rect 80886 5199 80888 5208
rect 80796 5170 80848 5176
rect 80940 5199 80942 5208
rect 80888 5170 80940 5176
rect 80900 4214 80928 5170
rect 81452 4729 81480 5222
rect 81438 4720 81494 4729
rect 81438 4655 81494 4664
rect 81636 4554 81664 5238
rect 81912 4690 81940 5607
rect 81900 4684 81952 4690
rect 81900 4626 81952 4632
rect 81624 4548 81676 4554
rect 81624 4490 81676 4496
rect 81636 4214 81664 4490
rect 80888 4208 80940 4214
rect 80888 4150 80940 4156
rect 81624 4208 81676 4214
rect 81624 4150 81676 4156
rect 81440 4072 81492 4078
rect 81440 4014 81492 4020
rect 81452 3194 81480 4014
rect 82188 3233 82216 7958
rect 82648 7449 82676 8910
rect 82740 7857 82768 9454
rect 83844 9042 83872 10367
rect 84580 9586 84608 10503
rect 85394 9888 85450 9897
rect 85394 9823 85450 9832
rect 86498 9888 86554 9897
rect 86498 9823 86554 9832
rect 84568 9580 84620 9586
rect 84568 9522 84620 9528
rect 84844 9512 84896 9518
rect 84844 9454 84896 9460
rect 83832 9036 83884 9042
rect 83832 8978 83884 8984
rect 84108 8968 84160 8974
rect 84108 8910 84160 8916
rect 84120 7993 84148 8910
rect 84856 8294 84884 9454
rect 85408 8974 85436 9823
rect 86512 8974 86540 9823
rect 86788 9586 86816 10503
rect 90824 10474 90876 10480
rect 91008 10532 91060 10538
rect 91008 10474 91060 10480
rect 94044 10532 94096 10538
rect 94044 10474 94096 10480
rect 90362 10296 90418 10305
rect 90362 10231 90418 10240
rect 90376 9722 90404 10231
rect 91020 10130 91048 10474
rect 92388 10464 92440 10470
rect 92388 10406 92440 10412
rect 91008 10124 91060 10130
rect 91008 10066 91060 10072
rect 90272 9716 90324 9722
rect 90272 9658 90324 9664
rect 90364 9716 90416 9722
rect 90364 9658 90416 9664
rect 86776 9580 86828 9586
rect 86776 9522 86828 9528
rect 89168 9580 89220 9586
rect 89168 9522 89220 9528
rect 90180 9580 90232 9586
rect 90180 9522 90232 9528
rect 87052 9512 87104 9518
rect 87052 9454 87104 9460
rect 87788 9512 87840 9518
rect 87788 9454 87840 9460
rect 85396 8968 85448 8974
rect 85396 8910 85448 8916
rect 86500 8968 86552 8974
rect 86500 8910 86552 8916
rect 85580 8900 85632 8906
rect 85580 8842 85632 8848
rect 84200 8288 84252 8294
rect 84200 8230 84252 8236
rect 84844 8288 84896 8294
rect 84844 8230 84896 8236
rect 84106 7984 84162 7993
rect 84106 7919 84162 7928
rect 82726 7848 82782 7857
rect 82726 7783 82782 7792
rect 82634 7440 82690 7449
rect 82634 7375 82690 7384
rect 84212 5846 84240 8230
rect 85592 8022 85620 8842
rect 86592 8832 86644 8838
rect 86592 8774 86644 8780
rect 85580 8016 85632 8022
rect 85580 7958 85632 7964
rect 85672 7812 85724 7818
rect 85672 7754 85724 7760
rect 84200 5840 84252 5846
rect 84200 5782 84252 5788
rect 84936 5772 84988 5778
rect 84936 5714 84988 5720
rect 84948 5642 84976 5714
rect 85578 5672 85634 5681
rect 84936 5636 84988 5642
rect 85578 5607 85580 5616
rect 84936 5578 84988 5584
rect 85632 5607 85634 5616
rect 85580 5578 85632 5584
rect 84948 5302 84976 5578
rect 82912 5296 82964 5302
rect 82912 5238 82964 5244
rect 84752 5296 84804 5302
rect 84936 5296 84988 5302
rect 84804 5244 84884 5250
rect 84752 5238 84884 5244
rect 84936 5238 84988 5244
rect 82924 4826 82952 5238
rect 84764 5222 84884 5238
rect 84660 5160 84712 5166
rect 84660 5102 84712 5108
rect 84752 5160 84804 5166
rect 84752 5102 84804 5108
rect 84672 5030 84700 5102
rect 84660 5024 84712 5030
rect 84660 4966 84712 4972
rect 84672 4826 84700 4966
rect 82912 4820 82964 4826
rect 82912 4762 82964 4768
rect 84660 4820 84712 4826
rect 84660 4762 84712 4768
rect 84764 4758 84792 5102
rect 84856 5030 84884 5222
rect 84844 5024 84896 5030
rect 84844 4966 84896 4972
rect 84752 4752 84804 4758
rect 84752 4694 84804 4700
rect 84016 4616 84068 4622
rect 84016 4558 84068 4564
rect 83648 4208 83700 4214
rect 83648 4150 83700 4156
rect 83660 3466 83688 4150
rect 83924 3936 83976 3942
rect 83924 3878 83976 3884
rect 83648 3460 83700 3466
rect 83700 3420 83780 3448
rect 83648 3402 83700 3408
rect 82174 3224 82230 3233
rect 81440 3188 81492 3194
rect 82174 3159 82230 3168
rect 81440 3130 81492 3136
rect 82358 3088 82414 3097
rect 82358 3023 82360 3032
rect 82412 3023 82414 3032
rect 82360 2994 82412 3000
rect 82084 2984 82136 2990
rect 82084 2926 82136 2932
rect 80152 1964 80204 1970
rect 80152 1906 80204 1912
rect 80060 1896 80112 1902
rect 80060 1838 80112 1844
rect 81348 1896 81400 1902
rect 81348 1838 81400 1844
rect 81440 1896 81492 1902
rect 81440 1838 81492 1844
rect 80072 1601 80100 1838
rect 81360 1601 81388 1838
rect 80058 1592 80114 1601
rect 80058 1527 80114 1536
rect 81346 1592 81402 1601
rect 81346 1527 81402 1536
rect 79968 1352 80020 1358
rect 77576 1294 77628 1300
rect 77942 1320 77998 1329
rect 77206 1048 77262 1057
rect 77206 983 77262 992
rect 77588 921 77616 1294
rect 79414 1320 79470 1329
rect 77942 1255 77998 1264
rect 78588 1284 78640 1290
rect 79968 1294 80020 1300
rect 79414 1255 79470 1264
rect 78588 1226 78640 1232
rect 77574 912 77630 921
rect 77574 847 77630 856
rect 78600 785 78628 1226
rect 79980 785 80008 1294
rect 81452 814 81480 1838
rect 82096 1329 82124 2926
rect 82360 2440 82412 2446
rect 82360 2382 82412 2388
rect 82082 1320 82138 1329
rect 82082 1255 82138 1264
rect 82372 950 82400 2382
rect 83752 2378 83780 3420
rect 83004 2372 83056 2378
rect 83004 2314 83056 2320
rect 83740 2372 83792 2378
rect 83740 2314 83792 2320
rect 82636 1896 82688 1902
rect 82636 1838 82688 1844
rect 82360 944 82412 950
rect 82360 886 82412 892
rect 82648 882 82676 1838
rect 83016 1601 83044 2314
rect 83740 1964 83792 1970
rect 83740 1906 83792 1912
rect 83752 1601 83780 1906
rect 83832 1896 83884 1902
rect 83832 1838 83884 1844
rect 83844 1737 83872 1838
rect 83830 1728 83886 1737
rect 83830 1663 83886 1672
rect 83002 1592 83058 1601
rect 83002 1527 83058 1536
rect 83738 1592 83794 1601
rect 83738 1527 83794 1536
rect 82728 1352 82780 1358
rect 82728 1294 82780 1300
rect 82636 876 82688 882
rect 82636 818 82688 824
rect 81440 808 81492 814
rect 78586 776 78642 785
rect 76748 740 76800 746
rect 78586 711 78642 720
rect 79966 776 80022 785
rect 81440 750 81492 756
rect 79966 711 80022 720
rect 76748 682 76800 688
rect 82740 649 82768 1294
rect 82726 640 82782 649
rect 74722 575 74778 584
rect 75000 604 75052 610
rect 82726 575 82782 584
rect 75000 546 75052 552
rect 83936 513 83964 3878
rect 84028 3738 84056 4558
rect 84948 4214 84976 5238
rect 85580 4752 85632 4758
rect 85580 4694 85632 4700
rect 85592 4554 85620 4694
rect 85580 4548 85632 4554
rect 85580 4490 85632 4496
rect 84936 4208 84988 4214
rect 84936 4150 84988 4156
rect 84016 3732 84068 3738
rect 84016 3674 84068 3680
rect 84948 3466 84976 4150
rect 85684 3641 85712 7754
rect 86604 7721 86632 8774
rect 86590 7712 86646 7721
rect 86590 7647 86646 7656
rect 87064 7585 87092 9454
rect 87800 9382 87828 9454
rect 88248 9444 88300 9450
rect 88248 9386 88300 9392
rect 87788 9376 87840 9382
rect 87788 9318 87840 9324
rect 87050 7576 87106 7585
rect 87050 7511 87106 7520
rect 86590 6624 86646 6633
rect 86590 6559 86646 6568
rect 86604 5302 86632 6559
rect 87696 6316 87748 6322
rect 87696 6258 87748 6264
rect 86776 5704 86828 5710
rect 86776 5646 86828 5652
rect 86592 5296 86644 5302
rect 86592 5238 86644 5244
rect 86788 4758 86816 5646
rect 86776 4752 86828 4758
rect 86776 4694 86828 4700
rect 86408 4548 86460 4554
rect 86684 4548 86736 4554
rect 86460 4508 86684 4536
rect 86408 4490 86460 4496
rect 86684 4490 86736 4496
rect 85670 3632 85726 3641
rect 85670 3567 85726 3576
rect 86590 3496 86646 3505
rect 84476 3460 84528 3466
rect 84476 3402 84528 3408
rect 84936 3460 84988 3466
rect 84936 3402 84988 3408
rect 85396 3460 85448 3466
rect 85448 3420 85620 3448
rect 86590 3431 86646 3440
rect 85396 3402 85448 3408
rect 84488 2990 84516 3402
rect 85592 3346 85620 3420
rect 85672 3392 85724 3398
rect 85670 3360 85672 3369
rect 86040 3392 86092 3398
rect 85724 3360 85726 3369
rect 85592 3318 85670 3346
rect 86040 3334 86092 3340
rect 85670 3295 85726 3304
rect 86052 3126 86080 3334
rect 86040 3120 86092 3126
rect 86040 3062 86092 3068
rect 86604 3058 86632 3431
rect 86592 3052 86644 3058
rect 86592 2994 86644 3000
rect 86788 2990 86816 4694
rect 87512 4480 87564 4486
rect 87512 4422 87564 4428
rect 87524 4282 87552 4422
rect 87512 4276 87564 4282
rect 87512 4218 87564 4224
rect 87708 3942 87736 6258
rect 87696 3936 87748 3942
rect 87696 3878 87748 3884
rect 87512 3732 87564 3738
rect 87512 3674 87564 3680
rect 84292 2984 84344 2990
rect 84292 2926 84344 2932
rect 84476 2984 84528 2990
rect 84476 2926 84528 2932
rect 86776 2984 86828 2990
rect 86776 2926 86828 2932
rect 84304 2417 84332 2926
rect 85396 2644 85448 2650
rect 85396 2586 85448 2592
rect 84290 2408 84346 2417
rect 84016 2372 84068 2378
rect 85408 2378 85436 2586
rect 84290 2343 84346 2352
rect 85396 2372 85448 2378
rect 84016 2314 84068 2320
rect 85396 2314 85448 2320
rect 84028 1902 84056 2314
rect 86406 2136 86462 2145
rect 86406 2071 86462 2080
rect 86420 1970 86448 2071
rect 86408 1964 86460 1970
rect 86408 1906 86460 1912
rect 84016 1896 84068 1902
rect 84016 1838 84068 1844
rect 86040 1896 86092 1902
rect 86040 1838 86092 1844
rect 86132 1896 86184 1902
rect 86132 1838 86184 1844
rect 86052 1766 86080 1838
rect 86040 1760 86092 1766
rect 86040 1702 86092 1708
rect 86052 1494 86080 1702
rect 86040 1488 86092 1494
rect 86040 1430 86092 1436
rect 85028 1352 85080 1358
rect 85028 1294 85080 1300
rect 85304 1352 85356 1358
rect 85304 1294 85356 1300
rect 84476 1284 84528 1290
rect 84476 1226 84528 1232
rect 84488 785 84516 1226
rect 85040 785 85068 1294
rect 85316 1193 85344 1294
rect 85302 1184 85358 1193
rect 85302 1119 85358 1128
rect 86144 1057 86172 1838
rect 86776 1352 86828 1358
rect 86776 1294 86828 1300
rect 87052 1352 87104 1358
rect 87524 1329 87552 3674
rect 87604 2304 87656 2310
rect 87604 2246 87656 2252
rect 87052 1294 87104 1300
rect 87510 1320 87566 1329
rect 86130 1048 86186 1057
rect 86130 983 86186 992
rect 86788 785 86816 1294
rect 84474 776 84530 785
rect 84474 711 84530 720
rect 85026 776 85082 785
rect 85026 711 85082 720
rect 86774 776 86830 785
rect 86774 711 86830 720
rect 83922 504 83978 513
rect 67546 439 67602 448
rect 72424 468 72476 474
rect 83922 439 83978 448
rect 72424 410 72476 416
rect 38842 303 38898 312
rect 41052 332 41104 338
rect 9404 274 9456 280
rect 41052 274 41104 280
rect 87064 241 87092 1294
rect 87510 1255 87566 1264
rect 87616 1193 87644 2246
rect 87800 1426 87828 9318
rect 88260 9178 88288 9386
rect 88800 9376 88852 9382
rect 88800 9318 88852 9324
rect 88338 9208 88394 9217
rect 88248 9172 88300 9178
rect 88338 9143 88340 9152
rect 88248 9114 88300 9120
rect 88392 9143 88394 9152
rect 88340 9114 88392 9120
rect 88338 8664 88394 8673
rect 88338 8599 88340 8608
rect 88392 8599 88394 8608
rect 88340 8570 88392 8576
rect 88812 8498 88840 9318
rect 89180 8974 89208 9522
rect 90192 9178 90220 9522
rect 90180 9172 90232 9178
rect 90180 9114 90232 9120
rect 88984 8968 89036 8974
rect 88984 8910 89036 8916
rect 89168 8968 89220 8974
rect 89168 8910 89220 8916
rect 89904 8968 89956 8974
rect 89904 8910 89956 8916
rect 88800 8492 88852 8498
rect 88800 8434 88852 8440
rect 88156 8424 88208 8430
rect 88156 8366 88208 8372
rect 87880 6792 87932 6798
rect 87880 6734 87932 6740
rect 87892 4622 87920 6734
rect 88064 5568 88116 5574
rect 88064 5510 88116 5516
rect 87880 4616 87932 4622
rect 87880 4558 87932 4564
rect 88076 4554 88104 5510
rect 88064 4548 88116 4554
rect 88064 4490 88116 4496
rect 88168 3482 88196 8366
rect 88076 3454 88196 3482
rect 88248 3528 88300 3534
rect 88248 3470 88300 3476
rect 88076 2530 88104 3454
rect 87984 2514 88104 2530
rect 87972 2508 88104 2514
rect 88024 2502 88104 2508
rect 87972 2450 88024 2456
rect 88076 1970 88104 2502
rect 88064 1964 88116 1970
rect 88064 1906 88116 1912
rect 88260 1442 88288 3470
rect 88340 2440 88392 2446
rect 88340 2382 88392 2388
rect 88352 1873 88380 2382
rect 88524 1896 88576 1902
rect 88338 1864 88394 1873
rect 88524 1838 88576 1844
rect 88338 1799 88394 1808
rect 87788 1420 87840 1426
rect 88260 1414 88380 1442
rect 88536 1426 88564 1838
rect 88996 1442 89024 8910
rect 89180 8498 89208 8910
rect 89628 8832 89680 8838
rect 89628 8774 89680 8780
rect 89168 8492 89220 8498
rect 89168 8434 89220 8440
rect 89640 6730 89668 8774
rect 89718 8120 89774 8129
rect 89718 8055 89774 8064
rect 89732 7750 89760 8055
rect 89720 7744 89772 7750
rect 89720 7686 89772 7692
rect 89628 6724 89680 6730
rect 89628 6666 89680 6672
rect 89916 5896 89944 8910
rect 89996 8560 90048 8566
rect 89996 8502 90048 8508
rect 89732 5868 89944 5896
rect 89536 5092 89588 5098
rect 89536 5034 89588 5040
rect 89168 3052 89220 3058
rect 89168 2994 89220 3000
rect 89074 2000 89130 2009
rect 89180 1970 89208 2994
rect 89352 2848 89404 2854
rect 89352 2790 89404 2796
rect 89260 2304 89312 2310
rect 89260 2246 89312 2252
rect 89074 1935 89130 1944
rect 89168 1964 89220 1970
rect 89088 1902 89116 1935
rect 89168 1906 89220 1912
rect 89076 1896 89128 1902
rect 89076 1838 89128 1844
rect 89074 1456 89130 1465
rect 87788 1362 87840 1368
rect 88352 1358 88380 1414
rect 88524 1420 88576 1426
rect 88996 1414 89074 1442
rect 89074 1391 89130 1400
rect 88524 1362 88576 1368
rect 89088 1358 89116 1391
rect 89272 1358 89300 2246
rect 88340 1352 88392 1358
rect 88340 1294 88392 1300
rect 89076 1352 89128 1358
rect 89076 1294 89128 1300
rect 89260 1352 89312 1358
rect 89364 1329 89392 2790
rect 89548 2378 89576 5034
rect 89732 2666 89760 5868
rect 89904 5024 89956 5030
rect 89904 4966 89956 4972
rect 89812 3392 89864 3398
rect 89812 3334 89864 3340
rect 89824 2922 89852 3334
rect 89812 2916 89864 2922
rect 89812 2858 89864 2864
rect 89640 2638 89760 2666
rect 89536 2372 89588 2378
rect 89536 2314 89588 2320
rect 89640 2009 89668 2638
rect 89824 2281 89852 2858
rect 89916 2553 89944 4966
rect 89902 2544 89958 2553
rect 89902 2479 89958 2488
rect 89904 2440 89956 2446
rect 89904 2382 89956 2388
rect 89810 2272 89866 2281
rect 89810 2207 89866 2216
rect 89626 2000 89682 2009
rect 89916 1970 89944 2382
rect 90008 1970 90036 8502
rect 90088 8288 90140 8294
rect 90088 8230 90140 8236
rect 90100 7886 90128 8230
rect 90088 7880 90140 7886
rect 90088 7822 90140 7828
rect 90284 6118 90312 9658
rect 91020 8974 91048 10066
rect 92400 10062 92428 10406
rect 94056 10402 94084 10474
rect 94044 10396 94096 10402
rect 94044 10338 94096 10344
rect 93216 10124 93268 10130
rect 93216 10066 93268 10072
rect 92388 10056 92440 10062
rect 92388 9998 92440 10004
rect 92204 9376 92256 9382
rect 92204 9318 92256 9324
rect 90732 8968 90784 8974
rect 91008 8968 91060 8974
rect 90732 8910 90784 8916
rect 90836 8928 91008 8956
rect 90454 8664 90510 8673
rect 90454 8599 90456 8608
rect 90508 8599 90510 8608
rect 90456 8570 90508 8576
rect 90744 8566 90772 8910
rect 90732 8560 90784 8566
rect 90732 8502 90784 8508
rect 90272 6112 90324 6118
rect 90272 6054 90324 6060
rect 90088 2984 90140 2990
rect 90086 2952 90088 2961
rect 90272 2984 90324 2990
rect 90140 2952 90142 2961
rect 90272 2926 90324 2932
rect 90086 2887 90142 2896
rect 90284 2310 90312 2926
rect 90836 2774 90864 8928
rect 91008 8910 91060 8916
rect 92020 8968 92072 8974
rect 92020 8910 92072 8916
rect 90916 8832 90968 8838
rect 90916 8774 90968 8780
rect 91652 8832 91704 8838
rect 91652 8774 91704 8780
rect 91834 8800 91890 8809
rect 90928 8498 90956 8774
rect 91664 8498 91692 8774
rect 91834 8735 91890 8744
rect 91848 8634 91876 8735
rect 91926 8664 91982 8673
rect 91836 8628 91888 8634
rect 91926 8599 91928 8608
rect 91836 8570 91888 8576
rect 91980 8599 91982 8608
rect 91928 8570 91980 8576
rect 90916 8492 90968 8498
rect 90916 8434 90968 8440
rect 91652 8492 91704 8498
rect 91652 8434 91704 8440
rect 91468 6384 91520 6390
rect 91468 6326 91520 6332
rect 91480 5409 91508 6326
rect 91466 5400 91522 5409
rect 91466 5335 91522 5344
rect 91744 5160 91796 5166
rect 91742 5128 91744 5137
rect 91928 5160 91980 5166
rect 91796 5128 91798 5137
rect 91928 5102 91980 5108
rect 91742 5063 91798 5072
rect 91008 4820 91060 4826
rect 91008 4762 91060 4768
rect 91020 4146 91048 4762
rect 91008 4140 91060 4146
rect 91008 4082 91060 4088
rect 91940 3466 91968 5102
rect 91652 3460 91704 3466
rect 91652 3402 91704 3408
rect 91928 3460 91980 3466
rect 91928 3402 91980 3408
rect 91664 2990 91692 3402
rect 91652 2984 91704 2990
rect 91652 2926 91704 2932
rect 90744 2746 90864 2774
rect 90272 2304 90324 2310
rect 90272 2246 90324 2252
rect 90744 1970 90772 2746
rect 91100 2440 91152 2446
rect 91100 2382 91152 2388
rect 91008 2372 91060 2378
rect 91008 2314 91060 2320
rect 90824 2304 90876 2310
rect 90824 2246 90876 2252
rect 89626 1935 89682 1944
rect 89904 1964 89956 1970
rect 89904 1906 89956 1912
rect 89996 1964 90048 1970
rect 89996 1906 90048 1912
rect 90732 1964 90784 1970
rect 90732 1906 90784 1912
rect 89536 1896 89588 1902
rect 89536 1838 89588 1844
rect 89548 1426 89576 1838
rect 90456 1760 90508 1766
rect 90456 1702 90508 1708
rect 89536 1420 89588 1426
rect 89536 1362 89588 1368
rect 90468 1358 90496 1702
rect 90456 1352 90508 1358
rect 89260 1294 89312 1300
rect 89350 1320 89406 1329
rect 90456 1294 90508 1300
rect 89350 1255 89406 1264
rect 90640 1216 90692 1222
rect 87602 1184 87658 1193
rect 90640 1158 90692 1164
rect 87602 1119 87658 1128
rect 90652 785 90680 1158
rect 90638 776 90694 785
rect 90638 711 90694 720
rect 90836 377 90864 2246
rect 91020 2106 91048 2314
rect 91112 2106 91140 2382
rect 91744 2304 91796 2310
rect 91744 2246 91796 2252
rect 91008 2100 91060 2106
rect 91008 2042 91060 2048
rect 91100 2100 91152 2106
rect 91100 2042 91152 2048
rect 91756 377 91784 2246
rect 92032 1902 92060 8910
rect 92216 2774 92244 9318
rect 92400 8974 92428 9998
rect 92848 9920 92900 9926
rect 92848 9862 92900 9868
rect 92940 9920 92992 9926
rect 92940 9862 92992 9868
rect 92860 9518 92888 9862
rect 92848 9512 92900 9518
rect 92848 9454 92900 9460
rect 92388 8968 92440 8974
rect 92388 8910 92440 8916
rect 92388 8832 92440 8838
rect 92388 8774 92440 8780
rect 92400 8498 92428 8774
rect 92388 8492 92440 8498
rect 92388 8434 92440 8440
rect 92952 8430 92980 9862
rect 93228 9382 93256 10066
rect 93490 9752 93546 9761
rect 93490 9687 93492 9696
rect 93544 9687 93546 9696
rect 93492 9658 93544 9664
rect 94136 9648 94188 9654
rect 94136 9590 94188 9596
rect 93676 9580 93728 9586
rect 93676 9522 93728 9528
rect 93400 9512 93452 9518
rect 93400 9454 93452 9460
rect 93216 9376 93268 9382
rect 93216 9318 93268 9324
rect 93228 8498 93256 9318
rect 93412 8974 93440 9454
rect 93688 8974 93716 9522
rect 93400 8968 93452 8974
rect 93400 8910 93452 8916
rect 93492 8968 93544 8974
rect 93492 8910 93544 8916
rect 93676 8968 93728 8974
rect 93676 8910 93728 8916
rect 93216 8492 93268 8498
rect 93216 8434 93268 8440
rect 92940 8424 92992 8430
rect 92940 8366 92992 8372
rect 93306 8392 93362 8401
rect 93306 8327 93362 8336
rect 93124 8288 93176 8294
rect 93124 8230 93176 8236
rect 93136 7886 93164 8230
rect 93320 8022 93348 8327
rect 93308 8016 93360 8022
rect 93308 7958 93360 7964
rect 93124 7880 93176 7886
rect 93412 7834 93440 8910
rect 93504 8498 93532 8910
rect 93492 8492 93544 8498
rect 93492 8434 93544 8440
rect 93124 7822 93176 7828
rect 93320 7806 93440 7834
rect 92848 6860 92900 6866
rect 92848 6802 92900 6808
rect 92480 6792 92532 6798
rect 92480 6734 92532 6740
rect 92492 5574 92520 6734
rect 92756 6248 92808 6254
rect 92662 6216 92718 6225
rect 92860 6202 92888 6802
rect 92808 6196 92888 6202
rect 92756 6190 92888 6196
rect 92768 6174 92888 6190
rect 92662 6151 92718 6160
rect 92676 5710 92704 6151
rect 92664 5704 92716 5710
rect 92664 5646 92716 5652
rect 92860 5642 92888 6174
rect 92848 5636 92900 5642
rect 92848 5578 92900 5584
rect 92480 5568 92532 5574
rect 92480 5510 92532 5516
rect 92664 5160 92716 5166
rect 92860 5148 92888 5578
rect 92716 5120 92888 5148
rect 92664 5102 92716 5108
rect 92676 4690 92704 5102
rect 92664 4684 92716 4690
rect 92664 4626 92716 4632
rect 92480 4480 92532 4486
rect 92478 4448 92480 4457
rect 92532 4448 92534 4457
rect 92478 4383 92534 4392
rect 92296 4004 92348 4010
rect 92296 3946 92348 3952
rect 92308 3058 92336 3946
rect 92296 3052 92348 3058
rect 92296 2994 92348 3000
rect 92308 2922 92336 2994
rect 92296 2916 92348 2922
rect 92296 2858 92348 2864
rect 92216 2746 92336 2774
rect 92308 1970 92336 2746
rect 92756 2440 92808 2446
rect 92756 2382 92808 2388
rect 92768 2106 92796 2382
rect 93032 2304 93084 2310
rect 93032 2246 93084 2252
rect 92756 2100 92808 2106
rect 92756 2042 92808 2048
rect 92296 1964 92348 1970
rect 92296 1906 92348 1912
rect 92020 1896 92072 1902
rect 92020 1838 92072 1844
rect 92020 1760 92072 1766
rect 92020 1702 92072 1708
rect 92032 1358 92060 1702
rect 92020 1352 92072 1358
rect 92020 1294 92072 1300
rect 92204 1216 92256 1222
rect 92204 1158 92256 1164
rect 92216 785 92244 1158
rect 92202 776 92258 785
rect 92202 711 92258 720
rect 93044 377 93072 2246
rect 93320 1970 93348 7806
rect 93400 6248 93452 6254
rect 93400 6190 93452 6196
rect 93412 5642 93440 6190
rect 93860 5840 93912 5846
rect 93860 5782 93912 5788
rect 93400 5636 93452 5642
rect 93400 5578 93452 5584
rect 93872 5302 93900 5782
rect 93860 5296 93912 5302
rect 93860 5238 93912 5244
rect 94148 5030 94176 9590
rect 94976 9382 95004 10542
rect 94320 9376 94372 9382
rect 94320 9318 94372 9324
rect 94964 9376 95016 9382
rect 94964 9318 95016 9324
rect 94332 8974 94360 9318
rect 94976 9042 95004 9318
rect 95068 9042 95096 10746
rect 97000 10606 97028 10746
rect 96988 10600 97040 10606
rect 96988 10542 97040 10548
rect 96712 10532 96764 10538
rect 96712 10474 96764 10480
rect 96436 10396 96488 10402
rect 96436 10338 96488 10344
rect 95974 9752 96030 9761
rect 95974 9687 95976 9696
rect 96028 9687 96030 9696
rect 96342 9752 96398 9761
rect 96342 9687 96344 9696
rect 95976 9658 96028 9664
rect 96396 9687 96398 9696
rect 96344 9658 96396 9664
rect 96160 9580 96212 9586
rect 96160 9522 96212 9528
rect 96172 9178 96200 9522
rect 96160 9172 96212 9178
rect 96160 9114 96212 9120
rect 94964 9036 95016 9042
rect 94964 8978 95016 8984
rect 95056 9036 95108 9042
rect 95056 8978 95108 8984
rect 94320 8968 94372 8974
rect 94320 8910 94372 8916
rect 94228 8900 94280 8906
rect 94228 8842 94280 8848
rect 94240 8362 94268 8842
rect 94412 8832 94464 8838
rect 94412 8774 94464 8780
rect 94424 8498 94452 8774
rect 94594 8664 94650 8673
rect 94594 8599 94596 8608
rect 94648 8599 94650 8608
rect 94870 8664 94926 8673
rect 94870 8599 94872 8608
rect 94596 8570 94648 8576
rect 94924 8599 94926 8608
rect 94872 8570 94924 8576
rect 94412 8492 94464 8498
rect 94412 8434 94464 8440
rect 94228 8356 94280 8362
rect 94228 8298 94280 8304
rect 94136 5024 94188 5030
rect 94136 4966 94188 4972
rect 94240 4842 94268 8298
rect 94976 8106 95004 8978
rect 95068 8242 95096 8978
rect 95148 8832 95200 8838
rect 95148 8774 95200 8780
rect 95160 8498 95188 8774
rect 96448 8498 96476 10338
rect 96724 9042 96752 10474
rect 97644 10266 97672 10814
rect 98368 10396 98420 10402
rect 98368 10338 98420 10344
rect 97632 10260 97684 10266
rect 97632 10202 97684 10208
rect 97540 10192 97592 10198
rect 97540 10134 97592 10140
rect 96804 9580 96856 9586
rect 96804 9522 96856 9528
rect 96712 9036 96764 9042
rect 96712 8978 96764 8984
rect 96620 8900 96672 8906
rect 96620 8842 96672 8848
rect 96632 8498 96660 8842
rect 96816 8634 96844 9522
rect 97172 9172 97224 9178
rect 97172 9114 97224 9120
rect 96896 9036 96948 9042
rect 96896 8978 96948 8984
rect 96804 8628 96856 8634
rect 96804 8570 96856 8576
rect 95148 8492 95200 8498
rect 95148 8434 95200 8440
rect 95976 8492 96028 8498
rect 95976 8434 96028 8440
rect 96436 8492 96488 8498
rect 96436 8434 96488 8440
rect 96620 8492 96672 8498
rect 96620 8434 96672 8440
rect 95068 8214 95188 8242
rect 94884 8078 95004 8106
rect 94320 7744 94372 7750
rect 94320 7686 94372 7692
rect 94332 7478 94360 7686
rect 94320 7472 94372 7478
rect 94320 7414 94372 7420
rect 94412 7472 94464 7478
rect 94412 7414 94464 7420
rect 94424 7274 94452 7414
rect 94412 7268 94464 7274
rect 94412 7210 94464 7216
rect 94502 6216 94558 6225
rect 94502 6151 94558 6160
rect 94516 5710 94544 6151
rect 94504 5704 94556 5710
rect 94504 5646 94556 5652
rect 94148 4814 94268 4842
rect 93768 4072 93820 4078
rect 93768 4014 93820 4020
rect 93780 2990 93808 4014
rect 93768 2984 93820 2990
rect 93768 2926 93820 2932
rect 93676 2440 93728 2446
rect 93676 2382 93728 2388
rect 93688 2106 93716 2382
rect 93860 2304 93912 2310
rect 93860 2246 93912 2252
rect 93676 2100 93728 2106
rect 93676 2042 93728 2048
rect 93308 1964 93360 1970
rect 93308 1906 93360 1912
rect 93308 1760 93360 1766
rect 93308 1702 93360 1708
rect 93320 1358 93348 1702
rect 93308 1352 93360 1358
rect 93308 1294 93360 1300
rect 93492 1216 93544 1222
rect 93872 1193 93900 2246
rect 94148 1970 94176 4814
rect 94410 4720 94466 4729
rect 94410 4655 94466 4664
rect 94424 4622 94452 4655
rect 94412 4616 94464 4622
rect 94318 4584 94374 4593
rect 94412 4558 94464 4564
rect 94318 4519 94374 4528
rect 94332 4146 94360 4519
rect 94320 4140 94372 4146
rect 94320 4082 94372 4088
rect 94228 3664 94280 3670
rect 94228 3606 94280 3612
rect 94240 3058 94268 3606
rect 94228 3052 94280 3058
rect 94228 2994 94280 3000
rect 94412 2440 94464 2446
rect 94412 2382 94464 2388
rect 94136 1964 94188 1970
rect 94136 1906 94188 1912
rect 94424 1562 94452 2382
rect 94596 2304 94648 2310
rect 94596 2246 94648 2252
rect 94412 1556 94464 1562
rect 94412 1498 94464 1504
rect 94608 1193 94636 2246
rect 94884 1358 94912 8078
rect 94964 7948 95016 7954
rect 94964 7890 95016 7896
rect 94976 4622 95004 7890
rect 95056 5568 95108 5574
rect 95056 5510 95108 5516
rect 94964 4616 95016 4622
rect 94964 4558 95016 4564
rect 95068 4554 95096 5510
rect 95056 4548 95108 4554
rect 95056 4490 95108 4496
rect 95068 3466 95096 4490
rect 95056 3460 95108 3466
rect 95056 3402 95108 3408
rect 95160 1970 95188 8214
rect 95238 6352 95294 6361
rect 95238 6287 95294 6296
rect 95252 4690 95280 6287
rect 95240 4684 95292 4690
rect 95240 4626 95292 4632
rect 95884 3528 95936 3534
rect 95882 3496 95884 3505
rect 95936 3496 95938 3505
rect 95882 3431 95938 3440
rect 95424 2440 95476 2446
rect 95424 2382 95476 2388
rect 95332 2304 95384 2310
rect 95332 2246 95384 2252
rect 95148 1964 95200 1970
rect 95148 1906 95200 1912
rect 94964 1896 95016 1902
rect 94964 1838 95016 1844
rect 94976 1358 95004 1838
rect 95240 1828 95292 1834
rect 95240 1770 95292 1776
rect 95252 1562 95280 1770
rect 95240 1556 95292 1562
rect 95240 1498 95292 1504
rect 94872 1352 94924 1358
rect 94872 1294 94924 1300
rect 94964 1352 95016 1358
rect 94964 1294 95016 1300
rect 95344 1193 95372 2246
rect 95436 2106 95464 2382
rect 95424 2100 95476 2106
rect 95424 2042 95476 2048
rect 95988 1834 96016 8434
rect 96448 8378 96476 8434
rect 96448 8362 96660 8378
rect 96448 8356 96672 8362
rect 96448 8350 96620 8356
rect 96620 8298 96672 8304
rect 96804 6112 96856 6118
rect 96804 6054 96856 6060
rect 96068 4208 96120 4214
rect 96068 4150 96120 4156
rect 96080 3058 96108 4150
rect 96160 4072 96212 4078
rect 96158 4040 96160 4049
rect 96212 4040 96214 4049
rect 96158 3975 96214 3984
rect 96618 3632 96674 3641
rect 96618 3567 96620 3576
rect 96672 3567 96674 3576
rect 96620 3538 96672 3544
rect 96712 3528 96764 3534
rect 96712 3470 96764 3476
rect 96068 3052 96120 3058
rect 96068 2994 96120 3000
rect 96344 2508 96396 2514
rect 96344 2450 96396 2456
rect 96252 2440 96304 2446
rect 96252 2382 96304 2388
rect 96068 2304 96120 2310
rect 96068 2246 96120 2252
rect 95976 1828 96028 1834
rect 95976 1770 96028 1776
rect 96080 1193 96108 2246
rect 96264 2106 96292 2382
rect 96356 2106 96384 2450
rect 96252 2100 96304 2106
rect 96252 2042 96304 2048
rect 96344 2100 96396 2106
rect 96344 2042 96396 2048
rect 96620 1760 96672 1766
rect 96620 1702 96672 1708
rect 96632 1358 96660 1702
rect 96620 1352 96672 1358
rect 96620 1294 96672 1300
rect 96528 1216 96580 1222
rect 93492 1158 93544 1164
rect 93858 1184 93914 1193
rect 93504 785 93532 1158
rect 93858 1119 93914 1128
rect 94594 1184 94650 1193
rect 94594 1119 94650 1128
rect 95330 1184 95386 1193
rect 95330 1119 95386 1128
rect 96066 1184 96122 1193
rect 96528 1158 96580 1164
rect 96066 1119 96122 1128
rect 93490 776 93546 785
rect 93490 711 93546 720
rect 96540 513 96568 1158
rect 96724 1018 96752 3470
rect 96816 2938 96844 6054
rect 96908 4026 96936 8978
rect 96908 3998 97028 4026
rect 96896 3936 96948 3942
rect 96896 3878 96948 3884
rect 96908 3058 96936 3878
rect 96896 3052 96948 3058
rect 96896 2994 96948 3000
rect 96816 2910 96936 2938
rect 96804 2848 96856 2854
rect 96804 2790 96856 2796
rect 96816 1834 96844 2790
rect 96908 2582 96936 2910
rect 97000 2854 97028 3998
rect 97184 2990 97212 9114
rect 97264 8832 97316 8838
rect 97264 8774 97316 8780
rect 97276 8498 97304 8774
rect 97446 8664 97502 8673
rect 97446 8599 97448 8608
rect 97500 8599 97502 8608
rect 97448 8570 97500 8576
rect 97264 8492 97316 8498
rect 97264 8434 97316 8440
rect 97552 3602 97580 10134
rect 97644 9042 97672 10202
rect 97998 9752 98054 9761
rect 97998 9687 98000 9696
rect 98052 9687 98054 9696
rect 98276 9716 98328 9722
rect 98000 9658 98052 9664
rect 98276 9658 98328 9664
rect 98000 9580 98052 9586
rect 98000 9522 98052 9528
rect 98012 9178 98040 9522
rect 98092 9512 98144 9518
rect 98092 9454 98144 9460
rect 98104 9178 98132 9454
rect 98288 9382 98316 9658
rect 98276 9376 98328 9382
rect 98276 9318 98328 9324
rect 98000 9172 98052 9178
rect 98000 9114 98052 9120
rect 98092 9172 98144 9178
rect 98092 9114 98144 9120
rect 97632 9036 97684 9042
rect 97632 8978 97684 8984
rect 98276 9036 98328 9042
rect 98276 8978 98328 8984
rect 97264 3596 97316 3602
rect 97264 3538 97316 3544
rect 97540 3596 97592 3602
rect 97540 3538 97592 3544
rect 97276 3398 97304 3538
rect 97644 3482 97672 8978
rect 98090 4312 98146 4321
rect 98090 4247 98146 4256
rect 97552 3454 97672 3482
rect 97816 3528 97868 3534
rect 98104 3516 98132 4247
rect 98184 3936 98236 3942
rect 98184 3878 98236 3884
rect 97868 3488 98132 3516
rect 97816 3470 97868 3476
rect 97264 3392 97316 3398
rect 97264 3334 97316 3340
rect 97172 2984 97224 2990
rect 97172 2926 97224 2932
rect 96988 2848 97040 2854
rect 96988 2790 97040 2796
rect 97356 2848 97408 2854
rect 97356 2790 97408 2796
rect 97368 2582 97396 2790
rect 96896 2576 96948 2582
rect 96896 2518 96948 2524
rect 97356 2576 97408 2582
rect 97356 2518 97408 2524
rect 97448 2508 97500 2514
rect 97448 2450 97500 2456
rect 96804 1828 96856 1834
rect 96804 1770 96856 1776
rect 97172 1760 97224 1766
rect 97172 1702 97224 1708
rect 97184 1358 97212 1702
rect 97172 1352 97224 1358
rect 97460 1329 97488 2450
rect 97552 1902 97580 3454
rect 98104 3058 98132 3488
rect 98092 3052 98144 3058
rect 98012 3012 98092 3040
rect 97630 2680 97686 2689
rect 97630 2615 97686 2624
rect 97644 2446 97672 2615
rect 98012 2496 98040 3012
rect 98092 2994 98144 3000
rect 97920 2480 98040 2496
rect 97908 2474 98040 2480
rect 97632 2440 97684 2446
rect 97960 2468 98040 2474
rect 98092 2508 98144 2514
rect 98196 2496 98224 3878
rect 98144 2468 98224 2496
rect 98092 2450 98144 2456
rect 97908 2416 97960 2422
rect 97632 2382 97684 2388
rect 97540 1896 97592 1902
rect 97540 1838 97592 1844
rect 98288 1426 98316 8978
rect 98380 1902 98408 10338
rect 98472 9042 98500 10814
rect 132868 10804 132920 10810
rect 132868 10746 132920 10752
rect 133696 10804 133748 10810
rect 133696 10746 133748 10752
rect 99380 10736 99432 10742
rect 99380 10678 99432 10684
rect 104348 10736 104400 10742
rect 104348 10678 104400 10684
rect 130568 10736 130620 10742
rect 130568 10678 130620 10684
rect 99288 10396 99340 10402
rect 99288 10338 99340 10344
rect 99300 9586 99328 10338
rect 99288 9580 99340 9586
rect 99288 9522 99340 9528
rect 99392 9466 99420 10678
rect 104360 10402 104388 10678
rect 104808 10668 104860 10674
rect 104808 10610 104860 10616
rect 103520 10396 103572 10402
rect 103520 10338 103572 10344
rect 104348 10396 104400 10402
rect 104348 10338 104400 10344
rect 103336 10328 103388 10334
rect 103242 10296 103298 10305
rect 103336 10270 103388 10276
rect 103242 10231 103298 10240
rect 102416 10056 102468 10062
rect 102416 9998 102468 10004
rect 101680 9988 101732 9994
rect 101680 9930 101732 9936
rect 100666 9752 100722 9761
rect 100666 9687 100668 9696
rect 100720 9687 100722 9696
rect 100668 9658 100720 9664
rect 99472 9580 99524 9586
rect 99472 9522 99524 9528
rect 100208 9580 100260 9586
rect 100208 9522 100260 9528
rect 99300 9438 99420 9466
rect 99300 9042 99328 9438
rect 99380 9376 99432 9382
rect 99380 9318 99432 9324
rect 98460 9036 98512 9042
rect 98460 8978 98512 8984
rect 99288 9036 99340 9042
rect 99288 8978 99340 8984
rect 99300 8838 99328 8978
rect 98460 8832 98512 8838
rect 98460 8774 98512 8780
rect 99288 8832 99340 8838
rect 99288 8774 99340 8780
rect 98472 8498 98500 8774
rect 98642 8664 98698 8673
rect 98642 8599 98644 8608
rect 98696 8599 98698 8608
rect 98644 8570 98696 8576
rect 98460 8492 98512 8498
rect 98460 8434 98512 8440
rect 99286 8256 99342 8265
rect 99286 8191 99342 8200
rect 99300 8022 99328 8191
rect 99288 8016 99340 8022
rect 99288 7958 99340 7964
rect 99392 7886 99420 9318
rect 99484 8974 99512 9522
rect 100116 9172 100168 9178
rect 100116 9114 100168 9120
rect 100024 9036 100076 9042
rect 100024 8978 100076 8984
rect 99472 8968 99524 8974
rect 99472 8910 99524 8916
rect 99564 8832 99616 8838
rect 99564 8774 99616 8780
rect 99380 7880 99432 7886
rect 99380 7822 99432 7828
rect 99012 6860 99064 6866
rect 99012 6802 99064 6808
rect 99024 6662 99052 6802
rect 99012 6656 99064 6662
rect 99012 6598 99064 6604
rect 99024 6458 99052 6598
rect 99012 6452 99064 6458
rect 99012 6394 99064 6400
rect 99380 4752 99432 4758
rect 99380 4694 99432 4700
rect 98552 4072 98604 4078
rect 98552 4014 98604 4020
rect 98460 3392 98512 3398
rect 98460 3334 98512 3340
rect 98472 2514 98500 3334
rect 98564 2650 98592 4014
rect 98920 4004 98972 4010
rect 98920 3946 98972 3952
rect 98932 3738 98960 3946
rect 98828 3732 98880 3738
rect 98828 3674 98880 3680
rect 98920 3732 98972 3738
rect 98920 3674 98972 3680
rect 98644 3664 98696 3670
rect 98644 3606 98696 3612
rect 98656 3398 98684 3606
rect 98736 3528 98788 3534
rect 98736 3470 98788 3476
rect 98644 3392 98696 3398
rect 98644 3334 98696 3340
rect 98656 3194 98684 3334
rect 98748 3194 98776 3470
rect 98644 3188 98696 3194
rect 98644 3130 98696 3136
rect 98736 3188 98788 3194
rect 98736 3130 98788 3136
rect 98840 2650 98868 3674
rect 99104 3664 99156 3670
rect 99104 3606 99156 3612
rect 99116 3466 99144 3606
rect 99104 3460 99156 3466
rect 99104 3402 99156 3408
rect 99392 2961 99420 4694
rect 99472 4548 99524 4554
rect 99472 4490 99524 4496
rect 99484 4321 99512 4490
rect 99470 4312 99526 4321
rect 99470 4247 99526 4256
rect 99472 3664 99524 3670
rect 99472 3606 99524 3612
rect 99484 3398 99512 3606
rect 99472 3392 99524 3398
rect 99472 3334 99524 3340
rect 99472 2984 99524 2990
rect 99378 2952 99434 2961
rect 99472 2926 99524 2932
rect 99378 2887 99434 2896
rect 98552 2644 98604 2650
rect 98552 2586 98604 2592
rect 98828 2644 98880 2650
rect 98828 2586 98880 2592
rect 98644 2576 98696 2582
rect 98644 2518 98696 2524
rect 98460 2508 98512 2514
rect 98460 2450 98512 2456
rect 98656 2106 98684 2518
rect 99010 2408 99066 2417
rect 99010 2343 99066 2352
rect 99196 2372 99248 2378
rect 99024 2310 99052 2343
rect 99196 2314 99248 2320
rect 99012 2304 99064 2310
rect 99012 2246 99064 2252
rect 98644 2100 98696 2106
rect 98644 2042 98696 2048
rect 98552 1964 98604 1970
rect 98552 1906 98604 1912
rect 98368 1896 98420 1902
rect 98368 1838 98420 1844
rect 98564 1766 98592 1906
rect 98552 1760 98604 1766
rect 98552 1702 98604 1708
rect 98276 1420 98328 1426
rect 98276 1362 98328 1368
rect 98564 1358 98592 1702
rect 99024 1494 99052 2246
rect 99208 1562 99236 2314
rect 99380 2032 99432 2038
rect 99380 1974 99432 1980
rect 99392 1562 99420 1974
rect 99484 1873 99512 2926
rect 99470 1864 99526 1873
rect 99470 1799 99526 1808
rect 99196 1556 99248 1562
rect 99196 1498 99248 1504
rect 99380 1556 99432 1562
rect 99380 1498 99432 1504
rect 99012 1488 99064 1494
rect 99012 1430 99064 1436
rect 99576 1426 99604 8774
rect 100036 8498 100064 8978
rect 100128 8974 100156 9114
rect 100116 8968 100168 8974
rect 100116 8910 100168 8916
rect 99932 8492 99984 8498
rect 99932 8434 99984 8440
rect 100024 8492 100076 8498
rect 100024 8434 100076 8440
rect 99944 7954 99972 8434
rect 100128 8378 100156 8910
rect 100220 8634 100248 9522
rect 100392 9376 100444 9382
rect 100392 9318 100444 9324
rect 100298 8664 100354 8673
rect 100208 8628 100260 8634
rect 100298 8599 100300 8608
rect 100208 8570 100260 8576
rect 100352 8599 100354 8608
rect 100300 8570 100352 8576
rect 100036 8350 100156 8378
rect 99932 7948 99984 7954
rect 99932 7890 99984 7896
rect 100036 7206 100064 8350
rect 100208 7404 100260 7410
rect 100208 7346 100260 7352
rect 100024 7200 100076 7206
rect 100024 7142 100076 7148
rect 99840 6928 99892 6934
rect 99840 6870 99892 6876
rect 99748 6180 99800 6186
rect 99748 6122 99800 6128
rect 99760 5914 99788 6122
rect 99748 5908 99800 5914
rect 99748 5850 99800 5856
rect 99656 5024 99708 5030
rect 99656 4966 99708 4972
rect 99668 3058 99696 4966
rect 99852 4758 99880 6870
rect 100114 6760 100170 6769
rect 100114 6695 100170 6704
rect 100128 6458 100156 6695
rect 100220 6458 100248 7346
rect 100300 6860 100352 6866
rect 100404 6848 100432 9318
rect 101692 8974 101720 9930
rect 102428 9926 102456 9998
rect 102416 9920 102468 9926
rect 102416 9862 102468 9868
rect 103256 9586 103284 10231
rect 103244 9580 103296 9586
rect 103244 9522 103296 9528
rect 102345 9276 102653 9285
rect 102345 9274 102351 9276
rect 102407 9274 102431 9276
rect 102487 9274 102511 9276
rect 102567 9274 102591 9276
rect 102647 9274 102653 9276
rect 102407 9222 102409 9274
rect 102589 9222 102591 9274
rect 102345 9220 102351 9222
rect 102407 9220 102431 9222
rect 102487 9220 102511 9222
rect 102567 9220 102591 9222
rect 102647 9220 102653 9222
rect 102345 9211 102653 9220
rect 102692 9172 102744 9178
rect 102692 9114 102744 9120
rect 101680 8968 101732 8974
rect 101680 8910 101732 8916
rect 100484 8900 100536 8906
rect 100484 8842 100536 8848
rect 100352 6820 100432 6848
rect 100300 6802 100352 6808
rect 100116 6452 100168 6458
rect 100116 6394 100168 6400
rect 100208 6452 100260 6458
rect 100208 6394 100260 6400
rect 99932 6316 99984 6322
rect 99932 6258 99984 6264
rect 99944 5778 99972 6258
rect 100116 6112 100168 6118
rect 100116 6054 100168 6060
rect 100128 5846 100156 6054
rect 100116 5840 100168 5846
rect 100116 5782 100168 5788
rect 99932 5772 99984 5778
rect 99932 5714 99984 5720
rect 99840 4752 99892 4758
rect 99892 4712 99972 4740
rect 99840 4694 99892 4700
rect 99748 4072 99800 4078
rect 99748 4014 99800 4020
rect 99760 3466 99788 4014
rect 99748 3460 99800 3466
rect 99748 3402 99800 3408
rect 99656 3052 99708 3058
rect 99656 2994 99708 3000
rect 99760 2514 99788 3402
rect 99840 2984 99892 2990
rect 99840 2926 99892 2932
rect 99748 2508 99800 2514
rect 99748 2450 99800 2456
rect 99852 1986 99880 2926
rect 99944 2922 99972 4712
rect 100208 4480 100260 4486
rect 100208 4422 100260 4428
rect 99932 2916 99984 2922
rect 99932 2858 99984 2864
rect 100220 2038 100248 4422
rect 100496 3074 100524 8842
rect 100668 8832 100720 8838
rect 100668 8774 100720 8780
rect 100680 8498 100708 8774
rect 100668 8492 100720 8498
rect 100668 8434 100720 8440
rect 102345 8188 102653 8197
rect 102345 8186 102351 8188
rect 102407 8186 102431 8188
rect 102487 8186 102511 8188
rect 102567 8186 102591 8188
rect 102647 8186 102653 8188
rect 102407 8134 102409 8186
rect 102589 8134 102591 8186
rect 102345 8132 102351 8134
rect 102407 8132 102431 8134
rect 102487 8132 102511 8134
rect 102567 8132 102591 8134
rect 102647 8132 102653 8134
rect 102345 8123 102653 8132
rect 102345 7100 102653 7109
rect 102345 7098 102351 7100
rect 102407 7098 102431 7100
rect 102487 7098 102511 7100
rect 102567 7098 102591 7100
rect 102647 7098 102653 7100
rect 102407 7046 102409 7098
rect 102589 7046 102591 7098
rect 102345 7044 102351 7046
rect 102407 7044 102431 7046
rect 102487 7044 102511 7046
rect 102567 7044 102591 7046
rect 102647 7044 102653 7046
rect 102345 7035 102653 7044
rect 100944 6996 100996 7002
rect 100944 6938 100996 6944
rect 100576 6792 100628 6798
rect 100628 6752 100892 6780
rect 100576 6734 100628 6740
rect 100760 6452 100812 6458
rect 100760 6394 100812 6400
rect 100668 6384 100720 6390
rect 100668 6326 100720 6332
rect 100574 5808 100630 5817
rect 100574 5743 100630 5752
rect 100588 5710 100616 5743
rect 100576 5704 100628 5710
rect 100576 5646 100628 5652
rect 100588 5137 100616 5646
rect 100680 5166 100708 6326
rect 100668 5160 100720 5166
rect 100574 5128 100630 5137
rect 100668 5102 100720 5108
rect 100574 5063 100630 5072
rect 100588 4690 100616 5063
rect 100576 4684 100628 4690
rect 100576 4626 100628 4632
rect 100576 3596 100628 3602
rect 100576 3538 100628 3544
rect 100404 3046 100524 3074
rect 100404 2990 100432 3046
rect 100392 2984 100444 2990
rect 100392 2926 100444 2932
rect 99760 1958 99880 1986
rect 100208 2032 100260 2038
rect 100208 1974 100260 1980
rect 100116 1964 100168 1970
rect 99564 1420 99616 1426
rect 99564 1362 99616 1368
rect 98552 1352 98604 1358
rect 97172 1294 97224 1300
rect 97446 1320 97502 1329
rect 98552 1294 98604 1300
rect 97446 1255 97502 1264
rect 97080 1216 97132 1222
rect 97080 1158 97132 1164
rect 98460 1216 98512 1222
rect 98460 1158 98512 1164
rect 96712 1012 96764 1018
rect 96712 954 96764 960
rect 97092 785 97120 1158
rect 98472 785 98500 1158
rect 97078 776 97134 785
rect 97078 711 97134 720
rect 98458 776 98514 785
rect 98458 711 98514 720
rect 98734 776 98790 785
rect 98734 711 98790 720
rect 96526 504 96582 513
rect 96526 439 96582 448
rect 98748 377 98776 711
rect 99760 474 99788 1958
rect 100116 1906 100168 1912
rect 99840 1896 99892 1902
rect 99840 1838 99892 1844
rect 99852 1358 99880 1838
rect 100128 1766 100156 1906
rect 100116 1760 100168 1766
rect 100116 1702 100168 1708
rect 100128 1358 100156 1702
rect 99840 1352 99892 1358
rect 99840 1294 99892 1300
rect 100116 1352 100168 1358
rect 100116 1294 100168 1300
rect 100588 1290 100616 3538
rect 100668 2984 100720 2990
rect 100668 2926 100720 2932
rect 100680 2106 100708 2926
rect 100772 2689 100800 6394
rect 100864 4321 100892 6752
rect 100956 5710 100984 6938
rect 101862 6896 101918 6905
rect 101862 6831 101918 6840
rect 101312 6792 101364 6798
rect 101312 6734 101364 6740
rect 100944 5704 100996 5710
rect 100944 5646 100996 5652
rect 100956 5234 100984 5646
rect 101324 5370 101352 6734
rect 101772 6656 101824 6662
rect 101772 6598 101824 6604
rect 101784 6322 101812 6598
rect 101772 6316 101824 6322
rect 101772 6258 101824 6264
rect 101876 5642 101904 6831
rect 102230 6624 102286 6633
rect 102230 6559 102286 6568
rect 102244 6254 102272 6559
rect 102232 6248 102284 6254
rect 102232 6190 102284 6196
rect 102345 6012 102653 6021
rect 102345 6010 102351 6012
rect 102407 6010 102431 6012
rect 102487 6010 102511 6012
rect 102567 6010 102591 6012
rect 102647 6010 102653 6012
rect 102407 5958 102409 6010
rect 102589 5958 102591 6010
rect 102345 5956 102351 5958
rect 102407 5956 102431 5958
rect 102487 5956 102511 5958
rect 102567 5956 102591 5958
rect 102647 5956 102653 5958
rect 102345 5947 102653 5956
rect 101864 5636 101916 5642
rect 101864 5578 101916 5584
rect 102048 5568 102100 5574
rect 102048 5510 102100 5516
rect 101312 5364 101364 5370
rect 101312 5306 101364 5312
rect 100944 5228 100996 5234
rect 100944 5170 100996 5176
rect 100956 4758 100984 5170
rect 102060 5098 102088 5510
rect 102048 5092 102100 5098
rect 102048 5034 102100 5040
rect 102345 4924 102653 4933
rect 102345 4922 102351 4924
rect 102407 4922 102431 4924
rect 102487 4922 102511 4924
rect 102567 4922 102591 4924
rect 102647 4922 102653 4924
rect 102407 4870 102409 4922
rect 102589 4870 102591 4922
rect 102345 4868 102351 4870
rect 102407 4868 102431 4870
rect 102487 4868 102511 4870
rect 102567 4868 102591 4870
rect 102647 4868 102653 4870
rect 102345 4859 102653 4868
rect 100944 4752 100996 4758
rect 100944 4694 100996 4700
rect 101312 4480 101364 4486
rect 101312 4422 101364 4428
rect 100850 4312 100906 4321
rect 100850 4247 100906 4256
rect 101324 3602 101352 4422
rect 101402 4312 101458 4321
rect 101402 4247 101458 4256
rect 101416 3602 101444 4247
rect 102048 4208 102100 4214
rect 102048 4150 102100 4156
rect 101588 3936 101640 3942
rect 101588 3878 101640 3884
rect 101312 3596 101364 3602
rect 101312 3538 101364 3544
rect 101404 3596 101456 3602
rect 101404 3538 101456 3544
rect 101324 3398 101352 3538
rect 101312 3392 101364 3398
rect 101312 3334 101364 3340
rect 101416 2990 101444 3538
rect 101496 3528 101548 3534
rect 101496 3470 101548 3476
rect 101508 3194 101536 3470
rect 101496 3188 101548 3194
rect 101496 3130 101548 3136
rect 101404 2984 101456 2990
rect 101404 2926 101456 2932
rect 100758 2680 100814 2689
rect 100758 2615 100814 2624
rect 101218 2408 101274 2417
rect 101218 2343 101220 2352
rect 101272 2343 101274 2352
rect 101220 2314 101272 2320
rect 100668 2100 100720 2106
rect 100668 2042 100720 2048
rect 100760 2100 100812 2106
rect 100760 2042 100812 2048
rect 100772 1601 100800 2042
rect 101312 1760 101364 1766
rect 101312 1702 101364 1708
rect 100758 1592 100814 1601
rect 100758 1527 100814 1536
rect 100576 1284 100628 1290
rect 100576 1226 100628 1232
rect 100024 1216 100076 1222
rect 100024 1158 100076 1164
rect 100574 1184 100630 1193
rect 100036 513 100064 1158
rect 100574 1119 100630 1128
rect 100588 921 100616 1119
rect 101324 921 101352 1702
rect 101600 1494 101628 3878
rect 101678 3224 101734 3233
rect 102060 3194 102088 4150
rect 102232 4072 102284 4078
rect 102232 4014 102284 4020
rect 101678 3159 101734 3168
rect 102048 3188 102100 3194
rect 101692 3058 101720 3159
rect 102048 3130 102100 3136
rect 101680 3052 101732 3058
rect 101680 2994 101732 3000
rect 102244 2990 102272 4014
rect 102345 3836 102653 3845
rect 102345 3834 102351 3836
rect 102407 3834 102431 3836
rect 102487 3834 102511 3836
rect 102567 3834 102591 3836
rect 102647 3834 102653 3836
rect 102407 3782 102409 3834
rect 102589 3782 102591 3834
rect 102345 3780 102351 3782
rect 102407 3780 102431 3782
rect 102487 3780 102511 3782
rect 102567 3780 102591 3782
rect 102647 3780 102653 3782
rect 102345 3771 102653 3780
rect 102704 3720 102732 9114
rect 103348 6730 103376 10270
rect 103532 10266 103560 10338
rect 103886 10296 103942 10305
rect 103520 10260 103572 10266
rect 103886 10231 103942 10240
rect 103520 10202 103572 10208
rect 103704 10192 103756 10198
rect 103704 10134 103756 10140
rect 103716 9722 103744 10134
rect 103704 9716 103756 9722
rect 103704 9658 103756 9664
rect 103900 9586 103928 10231
rect 104716 9716 104768 9722
rect 104716 9658 104768 9664
rect 103888 9580 103940 9586
rect 103888 9522 103940 9528
rect 104348 9036 104400 9042
rect 104348 8978 104400 8984
rect 104164 8900 104216 8906
rect 104164 8842 104216 8848
rect 104176 8430 104204 8842
rect 104164 8424 104216 8430
rect 104164 8366 104216 8372
rect 104164 7744 104216 7750
rect 104164 7686 104216 7692
rect 104176 7546 104204 7686
rect 104164 7540 104216 7546
rect 104164 7482 104216 7488
rect 102784 6724 102836 6730
rect 102784 6666 102836 6672
rect 103336 6724 103388 6730
rect 103336 6666 103388 6672
rect 102796 5710 102824 6666
rect 103152 6112 103204 6118
rect 103152 6054 103204 6060
rect 102784 5704 102836 5710
rect 102784 5646 102836 5652
rect 103164 5642 103192 6054
rect 103152 5636 103204 5642
rect 103152 5578 103204 5584
rect 102876 4004 102928 4010
rect 102876 3946 102928 3952
rect 102612 3692 102732 3720
rect 102612 3024 102640 3692
rect 102888 3602 102916 3946
rect 102876 3596 102928 3602
rect 102876 3538 102928 3544
rect 102888 3058 102916 3538
rect 103164 3398 103192 5578
rect 103520 5024 103572 5030
rect 103520 4966 103572 4972
rect 103152 3392 103204 3398
rect 103152 3334 103204 3340
rect 102876 3052 102928 3058
rect 102600 3018 102652 3024
rect 101864 2984 101916 2990
rect 101864 2926 101916 2932
rect 102232 2984 102284 2990
rect 102876 2994 102928 3000
rect 102600 2960 102652 2966
rect 102232 2926 102284 2932
rect 101588 1488 101640 1494
rect 101588 1430 101640 1436
rect 100574 912 100630 921
rect 100574 847 100630 856
rect 101310 912 101366 921
rect 101310 847 101366 856
rect 100392 740 100444 746
rect 100392 682 100444 688
rect 100022 504 100078 513
rect 99748 468 99800 474
rect 100404 474 100432 682
rect 101876 610 101904 2926
rect 103336 2848 103388 2854
rect 103336 2790 103388 2796
rect 102345 2748 102653 2757
rect 102345 2746 102351 2748
rect 102407 2746 102431 2748
rect 102487 2746 102511 2748
rect 102567 2746 102591 2748
rect 102647 2746 102653 2748
rect 102407 2694 102409 2746
rect 102589 2694 102591 2746
rect 102345 2692 102351 2694
rect 102407 2692 102431 2694
rect 102487 2692 102511 2694
rect 102567 2692 102591 2694
rect 102647 2692 102653 2694
rect 102345 2683 102653 2692
rect 103348 2582 103376 2790
rect 103336 2576 103388 2582
rect 103336 2518 103388 2524
rect 103426 2544 103482 2553
rect 103426 2479 103428 2488
rect 103480 2479 103482 2488
rect 103428 2450 103480 2456
rect 103532 2310 103560 4966
rect 104164 3664 104216 3670
rect 104164 3606 104216 3612
rect 103796 3596 103848 3602
rect 103796 3538 103848 3544
rect 103520 2304 103572 2310
rect 103808 2281 103836 3538
rect 104176 3534 104204 3606
rect 104164 3528 104216 3534
rect 104164 3470 104216 3476
rect 104176 2582 104204 3470
rect 104164 2576 104216 2582
rect 104164 2518 104216 2524
rect 104360 2514 104388 8978
rect 104440 6860 104492 6866
rect 104440 6802 104492 6808
rect 104452 2774 104480 6802
rect 104728 6458 104756 9658
rect 104820 8378 104848 10610
rect 129464 10600 129516 10606
rect 129464 10542 129516 10548
rect 125048 10464 125100 10470
rect 125048 10406 125100 10412
rect 125322 10432 125378 10441
rect 104898 10296 104954 10305
rect 104898 10231 104954 10240
rect 105634 10296 105690 10305
rect 105634 10231 105690 10240
rect 106278 10296 106334 10305
rect 106278 10231 106334 10240
rect 107198 10296 107254 10305
rect 107198 10231 107254 10240
rect 107750 10296 107806 10305
rect 107750 10231 107806 10240
rect 108394 10296 108450 10305
rect 108394 10231 108450 10240
rect 109038 10296 109094 10305
rect 109038 10231 109094 10240
rect 110050 10296 110106 10305
rect 110050 10231 110106 10240
rect 110786 10296 110842 10305
rect 110786 10231 110842 10240
rect 111522 10296 111578 10305
rect 111522 10231 111578 10240
rect 112350 10296 112406 10305
rect 112350 10231 112406 10240
rect 112902 10296 112958 10305
rect 112902 10231 112958 10240
rect 113546 10296 113602 10305
rect 113546 10231 113602 10240
rect 114190 10296 114246 10305
rect 114190 10231 114246 10240
rect 115202 10296 115258 10305
rect 115202 10231 115258 10240
rect 115938 10296 115994 10305
rect 115938 10231 115994 10240
rect 116674 10296 116730 10305
rect 116674 10231 116730 10240
rect 117318 10296 117374 10305
rect 117318 10231 117374 10240
rect 118054 10296 118110 10305
rect 118054 10231 118110 10240
rect 118698 10296 118754 10305
rect 118698 10231 118754 10240
rect 119342 10296 119398 10305
rect 119342 10231 119398 10240
rect 120354 10296 120410 10305
rect 120354 10231 120410 10240
rect 121090 10296 121146 10305
rect 121090 10231 121146 10240
rect 121366 10296 121422 10305
rect 121366 10231 121422 10240
rect 122654 10296 122710 10305
rect 122654 10231 122710 10240
rect 123206 10296 123262 10305
rect 123206 10231 123262 10240
rect 123942 10296 123998 10305
rect 123942 10231 123998 10240
rect 104912 9586 104940 10231
rect 105452 9716 105504 9722
rect 105452 9658 105504 9664
rect 104900 9580 104952 9586
rect 104900 9522 104952 9528
rect 105464 9110 105492 9658
rect 105648 9586 105676 10231
rect 105912 9716 105964 9722
rect 105912 9658 105964 9664
rect 105636 9580 105688 9586
rect 105636 9522 105688 9528
rect 105452 9104 105504 9110
rect 105452 9046 105504 9052
rect 104820 8350 105032 8378
rect 104900 8288 104952 8294
rect 104900 8230 104952 8236
rect 104716 6452 104768 6458
rect 104716 6394 104768 6400
rect 104716 6248 104768 6254
rect 104716 6190 104768 6196
rect 104728 5642 104756 6190
rect 104716 5636 104768 5642
rect 104716 5578 104768 5584
rect 104532 3936 104584 3942
rect 104532 3878 104584 3884
rect 104544 3738 104572 3878
rect 104532 3732 104584 3738
rect 104532 3674 104584 3680
rect 104544 3602 104572 3674
rect 104532 3596 104584 3602
rect 104532 3538 104584 3544
rect 104728 3482 104756 5578
rect 104912 5545 104940 8230
rect 104898 5536 104954 5545
rect 104898 5471 104954 5480
rect 105004 4146 105032 8350
rect 105728 8288 105780 8294
rect 105728 8230 105780 8236
rect 105176 7948 105228 7954
rect 105176 7890 105228 7896
rect 105188 7274 105216 7890
rect 105740 7886 105768 8230
rect 105636 7880 105688 7886
rect 105636 7822 105688 7828
rect 105728 7880 105780 7886
rect 105728 7822 105780 7828
rect 105648 7750 105676 7822
rect 105636 7744 105688 7750
rect 105636 7686 105688 7692
rect 105176 7268 105228 7274
rect 105176 7210 105228 7216
rect 105820 5024 105872 5030
rect 105820 4966 105872 4972
rect 105544 4752 105596 4758
rect 105544 4694 105596 4700
rect 105452 4548 105504 4554
rect 105452 4490 105504 4496
rect 104992 4140 105044 4146
rect 104992 4082 105044 4088
rect 105084 4072 105136 4078
rect 105084 4014 105136 4020
rect 104728 3466 104940 3482
rect 104728 3460 104952 3466
rect 104728 3454 104900 3460
rect 104900 3402 104952 3408
rect 104624 3392 104676 3398
rect 104624 3334 104676 3340
rect 104636 2990 104664 3334
rect 104624 2984 104676 2990
rect 104624 2926 104676 2932
rect 104452 2746 104848 2774
rect 104348 2508 104400 2514
rect 104348 2450 104400 2456
rect 104624 2440 104676 2446
rect 104624 2382 104676 2388
rect 104636 2310 104664 2382
rect 104624 2304 104676 2310
rect 103520 2246 103572 2252
rect 103794 2272 103850 2281
rect 104624 2246 104676 2252
rect 103794 2207 103850 2216
rect 102345 1660 102653 1669
rect 102345 1658 102351 1660
rect 102407 1658 102431 1660
rect 102487 1658 102511 1660
rect 102567 1658 102591 1660
rect 102647 1658 102653 1660
rect 102407 1606 102409 1658
rect 102589 1606 102591 1658
rect 102345 1604 102351 1606
rect 102407 1604 102431 1606
rect 102487 1604 102511 1606
rect 102567 1604 102591 1606
rect 102647 1604 102653 1606
rect 102345 1595 102653 1604
rect 103244 1420 103296 1426
rect 103244 1362 103296 1368
rect 101864 604 101916 610
rect 101864 546 101916 552
rect 103256 513 103284 1362
rect 103888 1352 103940 1358
rect 104716 1352 104768 1358
rect 103888 1294 103940 1300
rect 104622 1320 104678 1329
rect 103900 513 103928 1294
rect 104256 1284 104308 1290
rect 104716 1294 104768 1300
rect 104622 1255 104678 1264
rect 104256 1226 104308 1232
rect 104268 814 104296 1226
rect 104636 1222 104664 1255
rect 104624 1216 104676 1222
rect 104624 1158 104676 1164
rect 104256 808 104308 814
rect 104256 750 104308 756
rect 104728 513 104756 1294
rect 104820 1290 104848 2746
rect 104808 1284 104860 1290
rect 104808 1226 104860 1232
rect 105096 542 105124 4014
rect 105464 3670 105492 4490
rect 105556 4078 105584 4694
rect 105832 4622 105860 4966
rect 105820 4616 105872 4622
rect 105820 4558 105872 4564
rect 105924 4434 105952 9658
rect 106292 9586 106320 10231
rect 106280 9580 106332 9586
rect 106280 9522 106332 9528
rect 106096 9104 106148 9110
rect 106096 9046 106148 9052
rect 106108 7954 106136 9046
rect 107212 8974 107240 10231
rect 107764 9586 107792 10231
rect 108408 9586 108436 10231
rect 108948 9716 109000 9722
rect 108948 9658 109000 9664
rect 107752 9580 107804 9586
rect 107752 9522 107804 9528
rect 108396 9580 108448 9586
rect 108396 9522 108448 9528
rect 107568 9376 107620 9382
rect 107568 9318 107620 9324
rect 108212 9376 108264 9382
rect 108212 9318 108264 9324
rect 107580 9178 107608 9318
rect 107568 9172 107620 9178
rect 107568 9114 107620 9120
rect 107660 9172 107712 9178
rect 107660 9114 107712 9120
rect 106280 8968 106332 8974
rect 106280 8910 106332 8916
rect 107200 8968 107252 8974
rect 107200 8910 107252 8916
rect 106096 7948 106148 7954
rect 106096 7890 106148 7896
rect 106292 4622 106320 8910
rect 107108 8832 107160 8838
rect 107028 8792 107108 8820
rect 106556 7812 106608 7818
rect 106556 7754 106608 7760
rect 106372 7744 106424 7750
rect 106372 7686 106424 7692
rect 106384 6322 106412 7686
rect 106372 6316 106424 6322
rect 106372 6258 106424 6264
rect 106372 4684 106424 4690
rect 106372 4626 106424 4632
rect 106280 4616 106332 4622
rect 106280 4558 106332 4564
rect 105832 4406 105952 4434
rect 106280 4480 106332 4486
rect 106280 4422 106332 4428
rect 105832 4146 105860 4406
rect 105820 4140 105872 4146
rect 105820 4082 105872 4088
rect 105544 4072 105596 4078
rect 105544 4014 105596 4020
rect 106004 4072 106056 4078
rect 106004 4014 106056 4020
rect 105452 3664 105504 3670
rect 105452 3606 105504 3612
rect 105268 3596 105320 3602
rect 105268 3538 105320 3544
rect 105280 2650 105308 3538
rect 105268 2644 105320 2650
rect 105268 2586 105320 2592
rect 105450 1864 105506 1873
rect 105450 1799 105506 1808
rect 105464 1222 105492 1799
rect 105636 1352 105688 1358
rect 105636 1294 105688 1300
rect 105452 1216 105504 1222
rect 105452 1158 105504 1164
rect 105084 536 105136 542
rect 103242 504 103298 513
rect 100022 439 100078 448
rect 100392 468 100444 474
rect 99748 410 99800 416
rect 103242 439 103298 448
rect 103886 504 103942 513
rect 103886 439 103942 448
rect 104714 504 104770 513
rect 105648 513 105676 1294
rect 106016 1018 106044 4014
rect 106292 3194 106320 4422
rect 106280 3188 106332 3194
rect 106280 3130 106332 3136
rect 106188 2916 106240 2922
rect 106188 2858 106240 2864
rect 106200 1442 106228 2858
rect 106200 1414 106320 1442
rect 106188 1352 106240 1358
rect 106188 1294 106240 1300
rect 106004 1012 106056 1018
rect 106004 954 106056 960
rect 106200 513 106228 1294
rect 106292 1222 106320 1414
rect 106280 1216 106332 1222
rect 106280 1158 106332 1164
rect 105084 478 105136 484
rect 105634 504 105690 513
rect 104714 439 104770 448
rect 105634 439 105690 448
rect 106186 504 106242 513
rect 106384 474 106412 4626
rect 106568 2106 106596 7754
rect 106832 7336 106884 7342
rect 106832 7278 106884 7284
rect 106740 6724 106792 6730
rect 106740 6666 106792 6672
rect 106648 5092 106700 5098
rect 106648 5034 106700 5040
rect 106660 4758 106688 5034
rect 106648 4752 106700 4758
rect 106648 4694 106700 4700
rect 106752 4146 106780 6666
rect 106740 4140 106792 4146
rect 106740 4082 106792 4088
rect 106556 2100 106608 2106
rect 106556 2042 106608 2048
rect 106844 1193 106872 7278
rect 107028 5234 107056 8792
rect 107108 8774 107160 8780
rect 107672 7426 107700 9114
rect 108224 9042 108252 9318
rect 108212 9036 108264 9042
rect 108212 8978 108264 8984
rect 107936 8288 107988 8294
rect 107936 8230 107988 8236
rect 107948 8022 107976 8230
rect 107936 8016 107988 8022
rect 107856 7976 107936 8004
rect 107752 7948 107804 7954
rect 107752 7890 107804 7896
rect 107396 7410 107700 7426
rect 107384 7404 107700 7410
rect 107436 7398 107700 7404
rect 107384 7346 107436 7352
rect 107568 7336 107620 7342
rect 107568 7278 107620 7284
rect 107108 7268 107160 7274
rect 107108 7210 107160 7216
rect 107120 6934 107148 7210
rect 107108 6928 107160 6934
rect 107108 6870 107160 6876
rect 107292 6452 107344 6458
rect 107292 6394 107344 6400
rect 107304 5234 107332 6394
rect 107016 5228 107068 5234
rect 107016 5170 107068 5176
rect 107200 5228 107252 5234
rect 107200 5170 107252 5176
rect 107292 5228 107344 5234
rect 107292 5170 107344 5176
rect 106924 4004 106976 4010
rect 106924 3946 106976 3952
rect 106936 3398 106964 3946
rect 107108 3936 107160 3942
rect 107108 3878 107160 3884
rect 106924 3392 106976 3398
rect 106924 3334 106976 3340
rect 107120 3058 107148 3878
rect 107108 3052 107160 3058
rect 107108 2994 107160 3000
rect 107108 1964 107160 1970
rect 107108 1906 107160 1912
rect 106830 1184 106886 1193
rect 106830 1119 106886 1128
rect 107120 513 107148 1906
rect 107212 746 107240 5170
rect 107304 4078 107332 5170
rect 107292 4072 107344 4078
rect 107292 4014 107344 4020
rect 107384 4072 107436 4078
rect 107384 4014 107436 4020
rect 107292 2984 107344 2990
rect 107292 2926 107344 2932
rect 107304 2378 107332 2926
rect 107292 2372 107344 2378
rect 107292 2314 107344 2320
rect 107396 1562 107424 4014
rect 107476 2508 107528 2514
rect 107476 2450 107528 2456
rect 107384 1556 107436 1562
rect 107384 1498 107436 1504
rect 107488 1290 107516 2450
rect 107476 1284 107528 1290
rect 107476 1226 107528 1232
rect 107200 740 107252 746
rect 107200 682 107252 688
rect 107580 678 107608 7278
rect 107764 6934 107792 7890
rect 107856 7342 107884 7976
rect 107936 7958 107988 7964
rect 108396 7812 108448 7818
rect 108396 7754 108448 7760
rect 108408 7410 108436 7754
rect 108764 7744 108816 7750
rect 108764 7686 108816 7692
rect 108396 7404 108448 7410
rect 108396 7346 108448 7352
rect 107844 7336 107896 7342
rect 107844 7278 107896 7284
rect 107752 6928 107804 6934
rect 107752 6870 107804 6876
rect 107660 6112 107712 6118
rect 107660 6054 107712 6060
rect 107672 4758 107700 6054
rect 107660 4752 107712 4758
rect 107660 4694 107712 4700
rect 107764 4010 107792 6870
rect 107856 5794 107884 7278
rect 108120 6792 108172 6798
rect 108120 6734 108172 6740
rect 108132 6390 108160 6734
rect 108120 6384 108172 6390
rect 108120 6326 108172 6332
rect 107856 5766 108252 5794
rect 107936 5024 107988 5030
rect 107936 4966 107988 4972
rect 107752 4004 107804 4010
rect 107752 3946 107804 3952
rect 107660 2984 107712 2990
rect 107660 2926 107712 2932
rect 107672 2650 107700 2926
rect 107660 2644 107712 2650
rect 107660 2586 107712 2592
rect 107948 2514 107976 4966
rect 108224 4622 108252 5766
rect 108408 5273 108436 7346
rect 108580 7200 108632 7206
rect 108580 7142 108632 7148
rect 108592 6458 108620 7142
rect 108776 6866 108804 7686
rect 108764 6860 108816 6866
rect 108764 6802 108816 6808
rect 108580 6452 108632 6458
rect 108580 6394 108632 6400
rect 108672 6316 108724 6322
rect 108672 6258 108724 6264
rect 108684 6225 108712 6258
rect 108670 6216 108726 6225
rect 108670 6151 108726 6160
rect 108776 6118 108804 6802
rect 108764 6112 108816 6118
rect 108764 6054 108816 6060
rect 108854 5808 108910 5817
rect 108854 5743 108856 5752
rect 108908 5743 108910 5752
rect 108856 5714 108908 5720
rect 108764 5364 108816 5370
rect 108764 5306 108816 5312
rect 108394 5264 108450 5273
rect 108394 5199 108450 5208
rect 108396 5160 108448 5166
rect 108396 5102 108448 5108
rect 108408 4690 108436 5102
rect 108396 4684 108448 4690
rect 108396 4626 108448 4632
rect 108120 4616 108172 4622
rect 108120 4558 108172 4564
rect 108212 4616 108264 4622
rect 108264 4564 108436 4570
rect 108212 4558 108436 4564
rect 107936 2508 107988 2514
rect 107936 2450 107988 2456
rect 107752 1352 107804 1358
rect 107752 1294 107804 1300
rect 107568 672 107620 678
rect 107568 614 107620 620
rect 107764 513 107792 1294
rect 108132 1290 108160 4558
rect 108224 4542 108436 4558
rect 108776 4554 108804 5306
rect 108408 4146 108436 4542
rect 108764 4548 108816 4554
rect 108764 4490 108816 4496
rect 108856 4480 108908 4486
rect 108856 4422 108908 4428
rect 108396 4140 108448 4146
rect 108396 4082 108448 4088
rect 108408 2310 108436 4082
rect 108868 3602 108896 4422
rect 108960 3942 108988 9658
rect 109052 9586 109080 10231
rect 110064 9586 110092 10231
rect 110800 9586 110828 10231
rect 111536 9586 111564 10231
rect 109040 9580 109092 9586
rect 109040 9522 109092 9528
rect 110052 9580 110104 9586
rect 110052 9522 110104 9528
rect 110788 9580 110840 9586
rect 110788 9522 110840 9528
rect 111524 9580 111576 9586
rect 111524 9522 111576 9528
rect 111708 9444 111760 9450
rect 111708 9386 111760 9392
rect 111892 9444 111944 9450
rect 111892 9386 111944 9392
rect 109868 9376 109920 9382
rect 109868 9318 109920 9324
rect 110604 9376 110656 9382
rect 110604 9318 110656 9324
rect 109880 8838 109908 9318
rect 109868 8832 109920 8838
rect 109868 8774 109920 8780
rect 109868 7880 109920 7886
rect 109868 7822 109920 7828
rect 109132 7268 109184 7274
rect 109132 7210 109184 7216
rect 109040 6792 109092 6798
rect 109040 6734 109092 6740
rect 109052 6662 109080 6734
rect 109040 6656 109092 6662
rect 109040 6598 109092 6604
rect 109144 6440 109172 7210
rect 109224 6792 109276 6798
rect 109224 6734 109276 6740
rect 109316 6792 109368 6798
rect 109316 6734 109368 6740
rect 109052 6412 109172 6440
rect 109052 5778 109080 6412
rect 109040 5772 109092 5778
rect 109040 5714 109092 5720
rect 108948 3936 109000 3942
rect 108948 3878 109000 3884
rect 108856 3596 108908 3602
rect 108856 3538 108908 3544
rect 109038 3496 109094 3505
rect 109038 3431 109094 3440
rect 109052 2514 109080 3431
rect 109040 2508 109092 2514
rect 109040 2450 109092 2456
rect 108396 2304 108448 2310
rect 108396 2246 108448 2252
rect 109236 1358 109264 6734
rect 109328 6458 109356 6734
rect 109316 6452 109368 6458
rect 109316 6394 109368 6400
rect 109316 6248 109368 6254
rect 109316 6190 109368 6196
rect 109328 5642 109356 6190
rect 109316 5636 109368 5642
rect 109316 5578 109368 5584
rect 109406 5400 109462 5409
rect 109406 5335 109462 5344
rect 109420 4758 109448 5335
rect 109408 4752 109460 4758
rect 109408 4694 109460 4700
rect 109880 4554 109908 7822
rect 110512 7744 110564 7750
rect 110512 7686 110564 7692
rect 110524 7410 110552 7686
rect 110512 7404 110564 7410
rect 110512 7346 110564 7352
rect 110236 7268 110288 7274
rect 110236 7210 110288 7216
rect 109960 6656 110012 6662
rect 109960 6598 110012 6604
rect 109972 6322 110000 6598
rect 109960 6316 110012 6322
rect 109960 6258 110012 6264
rect 110248 5030 110276 7210
rect 110616 5166 110644 9318
rect 111720 8498 111748 9386
rect 111708 8492 111760 8498
rect 111708 8434 111760 8440
rect 111904 7750 111932 9386
rect 112364 8974 112392 10231
rect 112916 9586 112944 10231
rect 113560 9586 113588 10231
rect 113824 9920 113876 9926
rect 113824 9862 113876 9868
rect 113836 9722 113864 9862
rect 113824 9716 113876 9722
rect 113824 9658 113876 9664
rect 114204 9586 114232 10231
rect 115216 9586 115244 10231
rect 115952 9586 115980 10231
rect 116688 9586 116716 10231
rect 112904 9580 112956 9586
rect 112904 9522 112956 9528
rect 113548 9580 113600 9586
rect 113548 9522 113600 9528
rect 114192 9580 114244 9586
rect 114192 9522 114244 9528
rect 115204 9580 115256 9586
rect 115204 9522 115256 9528
rect 115940 9580 115992 9586
rect 115940 9522 115992 9528
rect 116676 9580 116728 9586
rect 116676 9522 116728 9528
rect 114284 9444 114336 9450
rect 114284 9386 114336 9392
rect 115664 9444 115716 9450
rect 115664 9386 115716 9392
rect 112720 9376 112772 9382
rect 112720 9318 112772 9324
rect 113364 9376 113416 9382
rect 113364 9318 113416 9324
rect 112732 9178 112760 9318
rect 112720 9172 112772 9178
rect 112720 9114 112772 9120
rect 112352 8968 112404 8974
rect 112352 8910 112404 8916
rect 111892 7744 111944 7750
rect 111892 7686 111944 7692
rect 112350 7440 112406 7449
rect 112076 7404 112128 7410
rect 112350 7375 112406 7384
rect 112076 7346 112128 7352
rect 110972 7336 111024 7342
rect 110972 7278 111024 7284
rect 110696 5364 110748 5370
rect 110696 5306 110748 5312
rect 110604 5160 110656 5166
rect 110604 5102 110656 5108
rect 110236 5024 110288 5030
rect 110236 4966 110288 4972
rect 110248 4758 110276 4966
rect 110236 4752 110288 4758
rect 110236 4694 110288 4700
rect 110708 4690 110736 5306
rect 110696 4684 110748 4690
rect 110696 4626 110748 4632
rect 110984 4622 111012 7278
rect 111248 6452 111300 6458
rect 111248 6394 111300 6400
rect 111260 5846 111288 6394
rect 112088 6390 112116 7346
rect 112076 6384 112128 6390
rect 112076 6326 112128 6332
rect 112088 6118 112116 6326
rect 112076 6112 112128 6118
rect 112076 6054 112128 6060
rect 111248 5840 111300 5846
rect 111524 5840 111576 5846
rect 111248 5782 111300 5788
rect 111522 5808 111524 5817
rect 111576 5808 111578 5817
rect 111260 5710 111288 5782
rect 111522 5743 111578 5752
rect 111248 5704 111300 5710
rect 111248 5646 111300 5652
rect 111800 5704 111852 5710
rect 111800 5646 111852 5652
rect 111812 4758 111840 5646
rect 111984 5160 112036 5166
rect 111984 5102 112036 5108
rect 111800 4752 111852 4758
rect 111800 4694 111852 4700
rect 109960 4616 110012 4622
rect 109960 4558 110012 4564
rect 110972 4616 111024 4622
rect 110972 4558 111024 4564
rect 109868 4548 109920 4554
rect 109868 4490 109920 4496
rect 109880 4214 109908 4490
rect 109868 4208 109920 4214
rect 109868 4150 109920 4156
rect 109316 3460 109368 3466
rect 109316 3402 109368 3408
rect 109328 3058 109356 3402
rect 109500 3120 109552 3126
rect 109500 3062 109552 3068
rect 109316 3052 109368 3058
rect 109316 2994 109368 3000
rect 109328 2378 109356 2994
rect 109512 2972 109540 3062
rect 109684 2984 109736 2990
rect 109512 2944 109684 2972
rect 109684 2926 109736 2932
rect 109316 2372 109368 2378
rect 109316 2314 109368 2320
rect 108396 1352 108448 1358
rect 108396 1294 108448 1300
rect 109040 1352 109092 1358
rect 109040 1294 109092 1300
rect 109224 1352 109276 1358
rect 109224 1294 109276 1300
rect 108120 1284 108172 1290
rect 108120 1226 108172 1232
rect 108408 513 108436 1294
rect 108856 1216 108908 1222
rect 108856 1158 108908 1164
rect 108868 1018 108896 1158
rect 108856 1012 108908 1018
rect 108856 954 108908 960
rect 108948 1012 109000 1018
rect 108948 954 109000 960
rect 108960 762 108988 954
rect 108868 746 108988 762
rect 108856 740 108988 746
rect 108908 734 108988 740
rect 108856 682 108908 688
rect 109052 513 109080 1294
rect 109868 1216 109920 1222
rect 109868 1158 109920 1164
rect 109880 1018 109908 1158
rect 109868 1012 109920 1018
rect 109868 954 109920 960
rect 109972 814 110000 4558
rect 110984 4486 111012 4558
rect 110972 4480 111024 4486
rect 110972 4422 111024 4428
rect 111340 4072 111392 4078
rect 110510 4040 110566 4049
rect 111340 4014 111392 4020
rect 110510 3975 110566 3984
rect 110236 3936 110288 3942
rect 110236 3878 110288 3884
rect 110248 3058 110276 3878
rect 110524 3602 110552 3975
rect 110512 3596 110564 3602
rect 110512 3538 110564 3544
rect 110972 3596 111024 3602
rect 110972 3538 111024 3544
rect 110236 3052 110288 3058
rect 110236 2994 110288 3000
rect 110984 1426 111012 3538
rect 110972 1420 111024 1426
rect 110972 1362 111024 1368
rect 110052 1352 110104 1358
rect 110052 1294 110104 1300
rect 110788 1352 110840 1358
rect 110788 1294 110840 1300
rect 109960 808 110012 814
rect 109960 750 110012 756
rect 110064 513 110092 1294
rect 110800 513 110828 1294
rect 111352 1222 111380 4014
rect 111524 1352 111576 1358
rect 111524 1294 111576 1300
rect 111340 1216 111392 1222
rect 111340 1158 111392 1164
rect 111536 513 111564 1294
rect 111996 610 112024 5102
rect 112364 4146 112392 7375
rect 112628 7336 112680 7342
rect 112628 7278 112680 7284
rect 112444 7268 112496 7274
rect 112444 7210 112496 7216
rect 112456 6866 112484 7210
rect 112444 6860 112496 6866
rect 112444 6802 112496 6808
rect 112640 6730 112668 7278
rect 113088 7200 113140 7206
rect 113088 7142 113140 7148
rect 112628 6724 112680 6730
rect 112628 6666 112680 6672
rect 112640 6254 112668 6666
rect 112718 6352 112774 6361
rect 112718 6287 112720 6296
rect 112772 6287 112774 6296
rect 112720 6258 112772 6264
rect 112628 6248 112680 6254
rect 112628 6190 112680 6196
rect 112640 5642 112668 6190
rect 112628 5636 112680 5642
rect 112628 5578 112680 5584
rect 112812 5160 112864 5166
rect 112812 5102 112864 5108
rect 112444 5092 112496 5098
rect 112444 5034 112496 5040
rect 112352 4140 112404 4146
rect 112352 4082 112404 4088
rect 112456 4010 112484 5034
rect 112536 4616 112588 4622
rect 112536 4558 112588 4564
rect 112548 4214 112576 4558
rect 112536 4208 112588 4214
rect 112536 4150 112588 4156
rect 112536 4072 112588 4078
rect 112536 4014 112588 4020
rect 112444 4004 112496 4010
rect 112444 3946 112496 3952
rect 112548 3097 112576 4014
rect 112720 3664 112772 3670
rect 112720 3606 112772 3612
rect 112732 3126 112760 3606
rect 112720 3120 112772 3126
rect 112534 3088 112590 3097
rect 112720 3062 112772 3068
rect 112534 3023 112590 3032
rect 112260 1964 112312 1970
rect 112260 1906 112312 1912
rect 111984 604 112036 610
rect 111984 546 112036 552
rect 112272 513 112300 1906
rect 112824 1442 112852 5102
rect 112996 4752 113048 4758
rect 112996 4694 113048 4700
rect 113008 4282 113036 4694
rect 112996 4276 113048 4282
rect 112996 4218 113048 4224
rect 112996 4004 113048 4010
rect 112996 3946 113048 3952
rect 113008 3602 113036 3946
rect 112996 3596 113048 3602
rect 112996 3538 113048 3544
rect 112824 1414 113036 1442
rect 112904 1352 112956 1358
rect 112904 1294 112956 1300
rect 112720 1216 112772 1222
rect 112720 1158 112772 1164
rect 112732 746 112760 1158
rect 112720 740 112772 746
rect 112720 682 112772 688
rect 112916 513 112944 1294
rect 113008 1290 113036 1414
rect 113100 1358 113128 7142
rect 113180 6860 113232 6866
rect 113180 6802 113232 6808
rect 113192 6769 113220 6802
rect 113178 6760 113234 6769
rect 113178 6695 113234 6704
rect 113376 6662 113404 9318
rect 113364 6656 113416 6662
rect 113364 6598 113416 6604
rect 113180 5160 113232 5166
rect 113180 5102 113232 5108
rect 114192 5160 114244 5166
rect 114192 5102 114244 5108
rect 113192 4486 113220 5102
rect 113640 5024 113692 5030
rect 113640 4966 113692 4972
rect 113732 5024 113784 5030
rect 113732 4966 113784 4972
rect 113652 4690 113680 4966
rect 113744 4758 113772 4966
rect 113916 4820 113968 4826
rect 113916 4762 113968 4768
rect 113732 4752 113784 4758
rect 113732 4694 113784 4700
rect 113640 4684 113692 4690
rect 113640 4626 113692 4632
rect 113928 4622 113956 4762
rect 113916 4616 113968 4622
rect 113916 4558 113968 4564
rect 113180 4480 113232 4486
rect 113364 4480 113416 4486
rect 113232 4440 113312 4468
rect 113180 4422 113232 4428
rect 113284 4298 113312 4440
rect 113362 4448 113364 4457
rect 113416 4448 113418 4457
rect 113362 4383 113418 4392
rect 113180 4276 113232 4282
rect 113284 4270 113588 4298
rect 113180 4218 113232 4224
rect 113192 3398 113220 4218
rect 113560 4146 113588 4270
rect 114204 4146 114232 5102
rect 114296 5098 114324 9386
rect 115020 9376 115072 9382
rect 115020 9318 115072 9324
rect 114560 8424 114612 8430
rect 114560 8366 114612 8372
rect 114376 6724 114428 6730
rect 114376 6666 114428 6672
rect 114388 6186 114416 6666
rect 114376 6180 114428 6186
rect 114376 6122 114428 6128
rect 114376 5636 114428 5642
rect 114376 5578 114428 5584
rect 114388 5302 114416 5578
rect 114376 5296 114428 5302
rect 114376 5238 114428 5244
rect 114284 5092 114336 5098
rect 114284 5034 114336 5040
rect 114388 4690 114416 5238
rect 114376 4684 114428 4690
rect 114376 4626 114428 4632
rect 114468 4684 114520 4690
rect 114468 4626 114520 4632
rect 114480 4486 114508 4626
rect 114468 4480 114520 4486
rect 114468 4422 114520 4428
rect 113548 4140 113600 4146
rect 113548 4082 113600 4088
rect 114192 4140 114244 4146
rect 114192 4082 114244 4088
rect 113456 4072 113508 4078
rect 113456 4014 113508 4020
rect 113468 3738 113496 4014
rect 113456 3732 113508 3738
rect 113456 3674 113508 3680
rect 113180 3392 113232 3398
rect 113180 3334 113232 3340
rect 113560 2990 113588 4082
rect 114572 3942 114600 8366
rect 114928 8016 114980 8022
rect 114834 7984 114890 7993
rect 114928 7958 114980 7964
rect 114834 7919 114890 7928
rect 114742 7848 114798 7857
rect 114742 7783 114798 7792
rect 114652 4480 114704 4486
rect 114652 4422 114704 4428
rect 114560 3936 114612 3942
rect 114560 3878 114612 3884
rect 113548 2984 113600 2990
rect 113548 2926 113600 2932
rect 114664 2922 114692 4422
rect 114756 4146 114784 7783
rect 114848 5794 114876 7919
rect 114940 6866 114968 7958
rect 114928 6860 114980 6866
rect 114928 6802 114980 6808
rect 114848 5766 114968 5794
rect 114744 4140 114796 4146
rect 114744 4082 114796 4088
rect 114836 4072 114888 4078
rect 114836 4014 114888 4020
rect 114652 2916 114704 2922
rect 114652 2858 114704 2864
rect 113272 1556 113324 1562
rect 113272 1498 113324 1504
rect 113088 1352 113140 1358
rect 113088 1294 113140 1300
rect 112996 1284 113048 1290
rect 112996 1226 113048 1232
rect 113284 1222 113312 1498
rect 113376 1414 113680 1442
rect 113376 1290 113404 1414
rect 113652 1358 113680 1414
rect 113548 1352 113600 1358
rect 113548 1294 113600 1300
rect 113640 1352 113692 1358
rect 113640 1294 113692 1300
rect 114192 1352 114244 1358
rect 114192 1294 114244 1300
rect 113364 1284 113416 1290
rect 113364 1226 113416 1232
rect 113272 1216 113324 1222
rect 113272 1158 113324 1164
rect 107106 504 107162 513
rect 106186 439 106242 448
rect 106372 468 106424 474
rect 100392 410 100444 416
rect 107106 439 107162 448
rect 107750 504 107806 513
rect 107750 439 107806 448
rect 108394 504 108450 513
rect 108394 439 108450 448
rect 109038 504 109094 513
rect 109038 439 109094 448
rect 110050 504 110106 513
rect 110050 439 110106 448
rect 110786 504 110842 513
rect 110786 439 110842 448
rect 111522 504 111578 513
rect 111522 439 111578 448
rect 112258 504 112314 513
rect 112258 439 112314 448
rect 112902 504 112958 513
rect 112902 439 112958 448
rect 106372 410 106424 416
rect 113560 377 113588 1294
rect 114204 649 114232 1294
rect 114848 950 114876 4014
rect 114940 3534 114968 5766
rect 115032 5370 115060 9318
rect 115572 8832 115624 8838
rect 115572 8774 115624 8780
rect 115112 5840 115164 5846
rect 115112 5782 115164 5788
rect 115124 5710 115152 5782
rect 115112 5704 115164 5710
rect 115112 5646 115164 5652
rect 115020 5364 115072 5370
rect 115020 5306 115072 5312
rect 115296 5024 115348 5030
rect 115296 4966 115348 4972
rect 115020 4548 115072 4554
rect 115020 4490 115072 4496
rect 114928 3528 114980 3534
rect 114928 3470 114980 3476
rect 115032 1222 115060 4490
rect 115308 4010 115336 4966
rect 115584 4146 115612 8774
rect 115572 4140 115624 4146
rect 115572 4082 115624 4088
rect 115296 4004 115348 4010
rect 115296 3946 115348 3952
rect 115308 3602 115336 3946
rect 115676 3602 115704 9386
rect 115848 9376 115900 9382
rect 115848 9318 115900 9324
rect 115860 8430 115888 9318
rect 117332 8974 117360 10231
rect 118068 9586 118096 10231
rect 118712 9586 118740 10231
rect 119356 9586 119384 10231
rect 120368 9586 120396 10231
rect 121104 9586 121132 10231
rect 121276 9920 121328 9926
rect 121276 9862 121328 9868
rect 118056 9580 118108 9586
rect 118056 9522 118108 9528
rect 118700 9580 118752 9586
rect 118700 9522 118752 9528
rect 119344 9580 119396 9586
rect 119344 9522 119396 9528
rect 120356 9580 120408 9586
rect 120356 9522 120408 9528
rect 121092 9580 121144 9586
rect 121092 9522 121144 9528
rect 121288 9518 121316 9862
rect 121276 9512 121328 9518
rect 121276 9454 121328 9460
rect 118332 9376 118384 9382
rect 118332 9318 118384 9324
rect 119160 9376 119212 9382
rect 119160 9318 119212 9324
rect 120172 9376 120224 9382
rect 120172 9318 120224 9324
rect 121000 9376 121052 9382
rect 121000 9318 121052 9324
rect 117320 8968 117372 8974
rect 117320 8910 117372 8916
rect 115848 8424 115900 8430
rect 115848 8366 115900 8372
rect 118240 8084 118292 8090
rect 118240 8026 118292 8032
rect 115756 6656 115808 6662
rect 115756 6598 115808 6604
rect 115768 5846 115796 6598
rect 115938 6488 115994 6497
rect 115938 6423 115994 6432
rect 115952 6390 115980 6423
rect 115940 6384 115992 6390
rect 115940 6326 115992 6332
rect 115848 6112 115900 6118
rect 115848 6054 115900 6060
rect 115860 5846 115888 6054
rect 115756 5840 115808 5846
rect 115756 5782 115808 5788
rect 115848 5840 115900 5846
rect 115848 5782 115900 5788
rect 116768 5704 116820 5710
rect 116768 5646 116820 5652
rect 116308 5296 116360 5302
rect 116308 5238 116360 5244
rect 116216 4684 116268 4690
rect 116216 4626 116268 4632
rect 116228 4593 116256 4626
rect 116214 4584 116270 4593
rect 116214 4519 116270 4528
rect 116032 4072 116084 4078
rect 116084 4032 116164 4060
rect 116032 4014 116084 4020
rect 115848 3732 115900 3738
rect 115848 3674 115900 3680
rect 115940 3732 115992 3738
rect 115940 3674 115992 3680
rect 115296 3596 115348 3602
rect 115296 3538 115348 3544
rect 115664 3596 115716 3602
rect 115664 3538 115716 3544
rect 115112 3528 115164 3534
rect 115112 3470 115164 3476
rect 115020 1216 115072 1222
rect 115020 1158 115072 1164
rect 114836 944 114888 950
rect 114836 886 114888 892
rect 115124 882 115152 3470
rect 115754 2952 115810 2961
rect 115754 2887 115756 2896
rect 115808 2887 115810 2896
rect 115756 2858 115808 2864
rect 115204 1352 115256 1358
rect 115204 1294 115256 1300
rect 115756 1352 115808 1358
rect 115756 1294 115808 1300
rect 115112 876 115164 882
rect 115112 818 115164 824
rect 115216 649 115244 1294
rect 115768 649 115796 1294
rect 115860 1222 115888 3674
rect 115952 3058 115980 3674
rect 116136 3641 116164 4032
rect 116122 3632 116178 3641
rect 116122 3567 116178 3576
rect 116136 3534 116164 3567
rect 116124 3528 116176 3534
rect 116124 3470 116176 3476
rect 116136 3058 116164 3470
rect 115940 3052 115992 3058
rect 115940 2994 115992 3000
rect 116124 3052 116176 3058
rect 116124 2994 116176 3000
rect 116320 2990 116348 5238
rect 116780 5166 116808 5646
rect 117410 5536 117466 5545
rect 117410 5471 117466 5480
rect 117424 5234 117452 5471
rect 117412 5228 117464 5234
rect 117412 5170 117464 5176
rect 116768 5160 116820 5166
rect 116768 5102 116820 5108
rect 117424 5030 117452 5170
rect 117596 5160 117648 5166
rect 117596 5102 117648 5108
rect 117412 5024 117464 5030
rect 117412 4966 117464 4972
rect 116400 4480 116452 4486
rect 116400 4422 116452 4428
rect 116412 4214 116440 4422
rect 116400 4208 116452 4214
rect 116400 4150 116452 4156
rect 116768 4072 116820 4078
rect 116768 4014 116820 4020
rect 116400 3936 116452 3942
rect 116400 3878 116452 3884
rect 116492 3936 116544 3942
rect 116492 3878 116544 3884
rect 116676 3936 116728 3942
rect 116676 3878 116728 3884
rect 116308 2984 116360 2990
rect 116308 2926 116360 2932
rect 116412 2106 116440 3878
rect 116504 3058 116532 3878
rect 116688 3126 116716 3878
rect 116780 3738 116808 4014
rect 116768 3732 116820 3738
rect 116768 3674 116820 3680
rect 117228 3596 117280 3602
rect 117228 3538 117280 3544
rect 116676 3120 116728 3126
rect 116676 3062 116728 3068
rect 116492 3052 116544 3058
rect 116492 2994 116544 3000
rect 116952 2984 117004 2990
rect 116952 2926 117004 2932
rect 116964 2854 116992 2926
rect 116952 2848 117004 2854
rect 116952 2790 117004 2796
rect 116400 2100 116452 2106
rect 116400 2042 116452 2048
rect 116676 1352 116728 1358
rect 116676 1294 116728 1300
rect 115848 1216 115900 1222
rect 115848 1158 115900 1164
rect 116688 649 116716 1294
rect 117240 1222 117268 3538
rect 117320 1964 117372 1970
rect 117320 1906 117372 1912
rect 117332 1465 117360 1906
rect 117318 1456 117374 1465
rect 117318 1391 117374 1400
rect 117228 1216 117280 1222
rect 117228 1158 117280 1164
rect 117608 785 117636 5102
rect 118056 5092 118108 5098
rect 118056 5034 118108 5040
rect 118068 4622 118096 5034
rect 118252 4690 118280 8026
rect 118344 5166 118372 9318
rect 118974 7712 119030 7721
rect 118974 7647 119030 7656
rect 118332 5160 118384 5166
rect 118332 5102 118384 5108
rect 118516 5160 118568 5166
rect 118516 5102 118568 5108
rect 118240 4684 118292 4690
rect 118240 4626 118292 4632
rect 118056 4616 118108 4622
rect 118056 4558 118108 4564
rect 118424 4616 118476 4622
rect 118424 4558 118476 4564
rect 117688 4072 117740 4078
rect 117688 4014 117740 4020
rect 117700 3126 117728 4014
rect 117688 3120 117740 3126
rect 117688 3062 117740 3068
rect 118056 1352 118108 1358
rect 118056 1294 118108 1300
rect 117594 776 117650 785
rect 117594 711 117650 720
rect 118068 649 118096 1294
rect 118436 1057 118464 4558
rect 118528 1222 118556 5102
rect 118884 4820 118936 4826
rect 118884 4762 118936 4768
rect 118896 4486 118924 4762
rect 118884 4480 118936 4486
rect 118884 4422 118936 4428
rect 118988 3602 119016 7647
rect 119068 6248 119120 6254
rect 119068 6190 119120 6196
rect 119080 5710 119108 6190
rect 119068 5704 119120 5710
rect 119068 5646 119120 5652
rect 119172 4622 119200 9318
rect 119988 6384 120040 6390
rect 119988 6326 120040 6332
rect 120000 5778 120028 6326
rect 120080 6112 120132 6118
rect 120080 6054 120132 6060
rect 120092 5914 120120 6054
rect 120080 5908 120132 5914
rect 120080 5850 120132 5856
rect 119988 5772 120040 5778
rect 119988 5714 120040 5720
rect 120080 5704 120132 5710
rect 119434 5672 119490 5681
rect 120080 5646 120132 5652
rect 119434 5607 119436 5616
rect 119488 5607 119490 5616
rect 119436 5578 119488 5584
rect 120092 5370 120120 5646
rect 120080 5364 120132 5370
rect 120080 5306 120132 5312
rect 120184 5250 120212 9318
rect 120816 8968 120868 8974
rect 120816 8910 120868 8916
rect 120828 8634 120856 8910
rect 120816 8628 120868 8634
rect 120816 8570 120868 8576
rect 120354 7576 120410 7585
rect 120354 7511 120410 7520
rect 120264 7404 120316 7410
rect 120264 7346 120316 7352
rect 120276 6186 120304 7346
rect 120264 6180 120316 6186
rect 120264 6122 120316 6128
rect 120368 6066 120396 7511
rect 120276 6038 120396 6066
rect 120276 5302 120304 6038
rect 120092 5222 120212 5250
rect 120264 5296 120316 5302
rect 120264 5238 120316 5244
rect 121012 5234 121040 9318
rect 121380 9178 121408 10231
rect 122668 9722 122696 10231
rect 122748 10192 122800 10198
rect 122748 10134 122800 10140
rect 122760 10062 122788 10134
rect 122748 10056 122800 10062
rect 122748 9998 122800 10004
rect 122656 9716 122708 9722
rect 122656 9658 122708 9664
rect 122472 9580 122524 9586
rect 122472 9522 122524 9528
rect 121460 9512 121512 9518
rect 121460 9454 121512 9460
rect 121368 9172 121420 9178
rect 121368 9114 121420 9120
rect 121276 9104 121328 9110
rect 121276 9046 121328 9052
rect 121288 8498 121316 9046
rect 121276 8492 121328 8498
rect 121276 8434 121328 8440
rect 121000 5228 121052 5234
rect 119436 5160 119488 5166
rect 119436 5102 119488 5108
rect 119448 5030 119476 5102
rect 119436 5024 119488 5030
rect 119436 4966 119488 4972
rect 119448 4622 119476 4966
rect 119804 4684 119856 4690
rect 119804 4626 119856 4632
rect 119160 4616 119212 4622
rect 119160 4558 119212 4564
rect 119252 4616 119304 4622
rect 119252 4558 119304 4564
rect 119436 4616 119488 4622
rect 119436 4558 119488 4564
rect 118976 3596 119028 3602
rect 118976 3538 119028 3544
rect 118700 1352 118752 1358
rect 118700 1294 118752 1300
rect 118516 1216 118568 1222
rect 118516 1158 118568 1164
rect 118422 1048 118478 1057
rect 118422 983 118478 992
rect 118712 649 118740 1294
rect 119264 1222 119292 4558
rect 119816 3670 119844 4626
rect 119988 3936 120040 3942
rect 119986 3904 119988 3913
rect 120040 3904 120042 3913
rect 119986 3839 120042 3848
rect 119804 3664 119856 3670
rect 119804 3606 119856 3612
rect 120092 3602 120120 5222
rect 121000 5170 121052 5176
rect 120448 5160 120500 5166
rect 120448 5102 120500 5108
rect 120816 5160 120868 5166
rect 120816 5102 120868 5108
rect 120356 5024 120408 5030
rect 120356 4966 120408 4972
rect 120264 4480 120316 4486
rect 120264 4422 120316 4428
rect 120080 3596 120132 3602
rect 120080 3538 120132 3544
rect 119344 3528 119396 3534
rect 119344 3470 119396 3476
rect 120172 3528 120224 3534
rect 120172 3470 120224 3476
rect 119356 2145 119384 3470
rect 119342 2136 119398 2145
rect 119342 2071 119398 2080
rect 119344 1352 119396 1358
rect 119344 1294 119396 1300
rect 119252 1216 119304 1222
rect 119252 1158 119304 1164
rect 119356 649 119384 1294
rect 120184 1222 120212 3470
rect 120276 3058 120304 4422
rect 120368 3641 120396 4966
rect 120354 3632 120410 3641
rect 120354 3567 120356 3576
rect 120408 3567 120410 3576
rect 120356 3538 120408 3544
rect 120264 3052 120316 3058
rect 120264 2994 120316 3000
rect 120356 1352 120408 1358
rect 120356 1294 120408 1300
rect 120172 1216 120224 1222
rect 120172 1158 120224 1164
rect 120368 649 120396 1294
rect 114190 640 114246 649
rect 114190 575 114246 584
rect 115202 640 115258 649
rect 115202 575 115258 584
rect 115754 640 115810 649
rect 115754 575 115810 584
rect 116674 640 116730 649
rect 116674 575 116730 584
rect 118054 640 118110 649
rect 118054 575 118110 584
rect 118698 640 118754 649
rect 118698 575 118754 584
rect 119342 640 119398 649
rect 119342 575 119398 584
rect 120354 640 120410 649
rect 120354 575 120410 584
rect 120460 513 120488 5102
rect 120724 5092 120776 5098
rect 120724 5034 120776 5040
rect 120736 4758 120764 5034
rect 120724 4752 120776 4758
rect 120724 4694 120776 4700
rect 120630 3360 120686 3369
rect 120630 3295 120686 3304
rect 120644 3126 120672 3295
rect 120632 3120 120684 3126
rect 120632 3062 120684 3068
rect 120828 1222 120856 5102
rect 121000 4072 121052 4078
rect 121000 4014 121052 4020
rect 120908 4004 120960 4010
rect 120908 3946 120960 3952
rect 120816 1216 120868 1222
rect 120816 1158 120868 1164
rect 120920 921 120948 3946
rect 121012 3670 121040 4014
rect 121000 3664 121052 3670
rect 121000 3606 121052 3612
rect 121288 2774 121316 8434
rect 121472 7546 121500 9454
rect 121736 9376 121788 9382
rect 121736 9318 121788 9324
rect 121748 8974 121776 9318
rect 122484 9178 122512 9522
rect 122760 9178 122788 9998
rect 122472 9172 122524 9178
rect 122472 9114 122524 9120
rect 122748 9172 122800 9178
rect 122748 9114 122800 9120
rect 122760 9058 122788 9114
rect 122668 9030 122788 9058
rect 122668 8974 122696 9030
rect 121644 8968 121696 8974
rect 121644 8910 121696 8916
rect 121736 8968 121788 8974
rect 121736 8910 121788 8916
rect 122656 8968 122708 8974
rect 122656 8910 122708 8916
rect 121460 7540 121512 7546
rect 121460 7482 121512 7488
rect 121196 2746 121316 2774
rect 121196 2038 121224 2746
rect 121184 2032 121236 2038
rect 121184 1974 121236 1980
rect 121656 1902 121684 8910
rect 121748 8498 121776 8910
rect 121736 8492 121788 8498
rect 121736 8434 121788 8440
rect 122668 8106 122696 8910
rect 123024 8832 123076 8838
rect 123024 8774 123076 8780
rect 123036 8498 123064 8774
rect 123220 8634 123248 10231
rect 123300 8968 123352 8974
rect 123300 8910 123352 8916
rect 123208 8628 123260 8634
rect 123208 8570 123260 8576
rect 123024 8492 123076 8498
rect 123024 8434 123076 8440
rect 122484 8078 122696 8106
rect 122104 6316 122156 6322
rect 122104 6258 122156 6264
rect 122012 6248 122064 6254
rect 122012 6190 122064 6196
rect 122024 6066 122052 6190
rect 122116 6186 122144 6258
rect 122104 6180 122156 6186
rect 122104 6122 122156 6128
rect 122196 6180 122248 6186
rect 122196 6122 122248 6128
rect 122208 6066 122236 6122
rect 122024 6038 122236 6066
rect 122196 5568 122248 5574
rect 122196 5510 122248 5516
rect 122208 5273 122236 5510
rect 122194 5264 122250 5273
rect 122194 5199 122196 5208
rect 122248 5199 122250 5208
rect 122196 5170 122248 5176
rect 121920 5024 121972 5030
rect 121920 4966 121972 4972
rect 121932 4690 121960 4966
rect 121920 4684 121972 4690
rect 121920 4626 121972 4632
rect 121920 4072 121972 4078
rect 121920 4014 121972 4020
rect 121932 2990 121960 4014
rect 121920 2984 121972 2990
rect 121920 2926 121972 2932
rect 122012 2440 122064 2446
rect 122012 2382 122064 2388
rect 122024 2106 122052 2382
rect 122012 2100 122064 2106
rect 122012 2042 122064 2048
rect 122484 1902 122512 8078
rect 122564 6112 122616 6118
rect 122564 6054 122616 6060
rect 122576 3534 122604 6054
rect 122656 4548 122708 4554
rect 122656 4490 122708 4496
rect 122668 4078 122696 4490
rect 122656 4072 122708 4078
rect 122656 4014 122708 4020
rect 122564 3528 122616 3534
rect 122564 3470 122616 3476
rect 122840 3392 122892 3398
rect 122840 3334 122892 3340
rect 122656 2304 122708 2310
rect 122656 2246 122708 2252
rect 121644 1896 121696 1902
rect 121644 1838 121696 1844
rect 122472 1896 122524 1902
rect 122472 1838 122524 1844
rect 121184 1760 121236 1766
rect 121184 1702 121236 1708
rect 121196 1358 121224 1702
rect 121656 1601 121684 1838
rect 121642 1592 121698 1601
rect 121642 1527 121644 1536
rect 121696 1527 121698 1536
rect 121644 1498 121696 1504
rect 121092 1352 121144 1358
rect 121092 1294 121144 1300
rect 121184 1352 121236 1358
rect 121184 1294 121236 1300
rect 120906 912 120962 921
rect 120906 847 120962 856
rect 121104 649 121132 1294
rect 121828 1216 121880 1222
rect 121828 1158 121880 1164
rect 121840 649 121868 1158
rect 122668 649 122696 2246
rect 122852 1970 122880 3334
rect 123312 2009 123340 8910
rect 123760 8832 123812 8838
rect 123760 8774 123812 8780
rect 123772 8498 123800 8774
rect 123956 8634 123984 10231
rect 124128 9988 124180 9994
rect 124128 9930 124180 9936
rect 124140 8974 124168 9930
rect 124588 9580 124640 9586
rect 124588 9522 124640 9528
rect 124600 9178 124628 9522
rect 124588 9172 124640 9178
rect 124588 9114 124640 9120
rect 125060 8974 125088 10406
rect 125322 10367 125378 10376
rect 127806 10432 127862 10441
rect 127806 10367 127862 10376
rect 125230 10296 125286 10305
rect 125230 10231 125286 10240
rect 125244 9722 125272 10231
rect 125232 9716 125284 9722
rect 125232 9658 125284 9664
rect 124128 8968 124180 8974
rect 124128 8910 124180 8916
rect 125048 8968 125100 8974
rect 125048 8910 125100 8916
rect 123944 8628 123996 8634
rect 123944 8570 123996 8576
rect 124140 8566 124168 8910
rect 124128 8560 124180 8566
rect 124128 8502 124180 8508
rect 123760 8492 123812 8498
rect 123760 8434 123812 8440
rect 123484 6656 123536 6662
rect 123484 6598 123536 6604
rect 123496 5234 123524 6598
rect 123484 5228 123536 5234
rect 123484 5170 123536 5176
rect 123392 4276 123444 4282
rect 123392 4218 123444 4224
rect 123404 4162 123432 4218
rect 123668 4208 123720 4214
rect 123404 4156 123668 4162
rect 123404 4150 123720 4156
rect 124140 4162 124168 8502
rect 125060 8430 125088 8910
rect 125336 8634 125364 10367
rect 126334 10296 126390 10305
rect 126334 10231 126390 10240
rect 126794 10296 126850 10305
rect 126794 10231 126850 10240
rect 125876 9512 125928 9518
rect 125876 9454 125928 9460
rect 125888 8974 125916 9454
rect 125876 8968 125928 8974
rect 125876 8910 125928 8916
rect 125416 8832 125468 8838
rect 125416 8774 125468 8780
rect 125324 8628 125376 8634
rect 125324 8570 125376 8576
rect 125428 8498 125456 8774
rect 125888 8566 125916 8910
rect 126152 8832 126204 8838
rect 126152 8774 126204 8780
rect 125876 8560 125928 8566
rect 125876 8502 125928 8508
rect 125416 8492 125468 8498
rect 125416 8434 125468 8440
rect 125048 8424 125100 8430
rect 125048 8366 125100 8372
rect 123404 4134 123708 4150
rect 124140 4134 124260 4162
rect 124036 3936 124088 3942
rect 124036 3878 124088 3884
rect 123576 3120 123628 3126
rect 123576 3062 123628 3068
rect 123298 2000 123354 2009
rect 122840 1964 122892 1970
rect 123298 1935 123354 1944
rect 122840 1906 122892 1912
rect 123312 1902 123340 1935
rect 123300 1896 123352 1902
rect 123300 1838 123352 1844
rect 122932 1760 122984 1766
rect 122932 1702 122984 1708
rect 122944 1358 122972 1702
rect 122932 1352 122984 1358
rect 122932 1294 122984 1300
rect 123588 1290 123616 3062
rect 123760 1760 123812 1766
rect 123760 1702 123812 1708
rect 123772 1358 123800 1702
rect 123760 1352 123812 1358
rect 123760 1294 123812 1300
rect 123576 1284 123628 1290
rect 123576 1226 123628 1232
rect 123116 1216 123168 1222
rect 123116 1158 123168 1164
rect 123944 1216 123996 1222
rect 123944 1158 123996 1164
rect 123128 649 123156 1158
rect 123956 649 123984 1158
rect 121090 640 121146 649
rect 121090 575 121146 584
rect 121826 640 121882 649
rect 121826 575 121882 584
rect 122654 640 122710 649
rect 122654 575 122710 584
rect 123114 640 123170 649
rect 123114 575 123170 584
rect 123942 640 123998 649
rect 123942 575 123998 584
rect 124048 513 124076 3878
rect 124232 2802 124260 4134
rect 124312 4072 124364 4078
rect 124312 4014 124364 4020
rect 124324 2854 124352 4014
rect 124140 2774 124260 2802
rect 124312 2848 124364 2854
rect 124312 2790 124364 2796
rect 124140 1970 124168 2774
rect 124496 2440 124548 2446
rect 124496 2382 124548 2388
rect 124508 2106 124536 2382
rect 124772 2304 124824 2310
rect 124772 2246 124824 2252
rect 124496 2100 124548 2106
rect 124496 2042 124548 2048
rect 124128 1964 124180 1970
rect 124128 1906 124180 1912
rect 124784 649 124812 2246
rect 125060 1970 125088 8366
rect 125600 6724 125652 6730
rect 125600 6666 125652 6672
rect 125140 6316 125192 6322
rect 125140 6258 125192 6264
rect 125152 5574 125180 6258
rect 125612 6186 125640 6666
rect 125600 6180 125652 6186
rect 125600 6122 125652 6128
rect 125140 5568 125192 5574
rect 125140 5510 125192 5516
rect 125888 2774 125916 8502
rect 126164 8498 126192 8774
rect 126348 8634 126376 10231
rect 126704 10124 126756 10130
rect 126704 10066 126756 10072
rect 126716 8974 126744 10066
rect 126704 8968 126756 8974
rect 126704 8910 126756 8916
rect 126336 8628 126388 8634
rect 126336 8570 126388 8576
rect 126152 8492 126204 8498
rect 126152 8434 126204 8440
rect 125888 2746 126008 2774
rect 125980 1970 126008 2746
rect 126244 2440 126296 2446
rect 126244 2382 126296 2388
rect 126256 2106 126284 2382
rect 126336 2304 126388 2310
rect 126336 2246 126388 2252
rect 126244 2100 126296 2106
rect 126244 2042 126296 2048
rect 125048 1964 125100 1970
rect 125048 1906 125100 1912
rect 125968 1964 126020 1970
rect 125968 1906 126020 1912
rect 125416 1760 125468 1766
rect 125416 1702 125468 1708
rect 125428 1358 125456 1702
rect 125416 1352 125468 1358
rect 125416 1294 125468 1300
rect 125324 1216 125376 1222
rect 125324 1158 125376 1164
rect 125336 649 125364 1158
rect 126348 649 126376 2246
rect 126716 1970 126744 8910
rect 126808 8634 126836 10231
rect 127624 9920 127676 9926
rect 127624 9862 127676 9868
rect 127164 9036 127216 9042
rect 127164 8978 127216 8984
rect 127176 8838 127204 8978
rect 126888 8832 126940 8838
rect 126888 8774 126940 8780
rect 127164 8832 127216 8838
rect 127164 8774 127216 8780
rect 126796 8628 126848 8634
rect 126796 8570 126848 8576
rect 126900 8498 126928 8774
rect 127636 8498 127664 9862
rect 127820 9178 127848 10367
rect 127898 10296 127954 10305
rect 127898 10231 127954 10240
rect 128818 10296 128874 10305
rect 128818 10231 128874 10240
rect 127912 9722 127940 10231
rect 128832 9722 128860 10231
rect 127900 9716 127952 9722
rect 127900 9658 127952 9664
rect 128820 9716 128872 9722
rect 128820 9658 128872 9664
rect 129476 9586 129504 10542
rect 129646 10296 129702 10305
rect 129646 10231 129702 10240
rect 130474 10296 130530 10305
rect 130474 10231 130530 10240
rect 129660 9722 129688 10231
rect 129648 9716 129700 9722
rect 129648 9658 129700 9664
rect 127992 9580 128044 9586
rect 127992 9522 128044 9528
rect 128636 9580 128688 9586
rect 128636 9522 128688 9528
rect 129464 9580 129516 9586
rect 129464 9522 129516 9528
rect 130384 9580 130436 9586
rect 130384 9522 130436 9528
rect 127808 9172 127860 9178
rect 127808 9114 127860 9120
rect 127808 8900 127860 8906
rect 127808 8842 127860 8848
rect 127820 8498 127848 8842
rect 128004 8634 128032 9522
rect 128268 8968 128320 8974
rect 128268 8910 128320 8916
rect 128280 8838 128308 8910
rect 128268 8832 128320 8838
rect 128268 8774 128320 8780
rect 127992 8628 128044 8634
rect 127992 8570 128044 8576
rect 126888 8492 126940 8498
rect 126888 8434 126940 8440
rect 127624 8492 127676 8498
rect 127624 8434 127676 8440
rect 127808 8492 127860 8498
rect 127808 8434 127860 8440
rect 127636 1970 127664 8434
rect 127900 2440 127952 2446
rect 127900 2382 127952 2388
rect 127808 2304 127860 2310
rect 127808 2246 127860 2252
rect 126704 1964 126756 1970
rect 126704 1906 126756 1912
rect 127624 1964 127676 1970
rect 127624 1906 127676 1912
rect 127072 1760 127124 1766
rect 127072 1702 127124 1708
rect 127084 1358 127112 1702
rect 127072 1352 127124 1358
rect 127072 1294 127124 1300
rect 126796 1216 126848 1222
rect 126796 1158 126848 1164
rect 126808 649 126836 1158
rect 127820 649 127848 2246
rect 127912 2106 127940 2382
rect 127900 2100 127952 2106
rect 127900 2042 127952 2048
rect 128280 1358 128308 8774
rect 128648 8634 128676 9522
rect 129096 9444 129148 9450
rect 129096 9386 129148 9392
rect 128728 8900 128780 8906
rect 128728 8842 128780 8848
rect 128636 8628 128688 8634
rect 128636 8570 128688 8576
rect 128740 8566 128768 8842
rect 129004 8832 129056 8838
rect 129004 8774 129056 8780
rect 128728 8560 128780 8566
rect 128728 8502 128780 8508
rect 129016 8362 129044 8774
rect 129108 8498 129136 9386
rect 129280 9376 129332 9382
rect 129280 9318 129332 9324
rect 129292 9042 129320 9318
rect 129280 9036 129332 9042
rect 129280 8978 129332 8984
rect 129096 8492 129148 8498
rect 129096 8434 129148 8440
rect 129004 8356 129056 8362
rect 129004 8298 129056 8304
rect 129108 6914 129136 8434
rect 129476 6914 129504 9522
rect 130396 9042 130424 9522
rect 130384 9036 130436 9042
rect 130384 8978 130436 8984
rect 129556 8968 129608 8974
rect 129556 8910 129608 8916
rect 129568 8498 129596 8910
rect 130488 8634 130516 10231
rect 130476 8628 130528 8634
rect 130476 8570 130528 8576
rect 129556 8492 129608 8498
rect 129556 8434 129608 8440
rect 130580 8430 130608 10678
rect 131120 10532 131172 10538
rect 131120 10474 131172 10480
rect 131132 8974 131160 10474
rect 131856 10328 131908 10334
rect 131486 10296 131542 10305
rect 131856 10270 131908 10276
rect 132314 10296 132370 10305
rect 131486 10231 131542 10240
rect 131500 9722 131528 10231
rect 131488 9716 131540 9722
rect 131488 9658 131540 9664
rect 131396 9580 131448 9586
rect 131396 9522 131448 9528
rect 131408 9178 131436 9522
rect 131396 9172 131448 9178
rect 131396 9114 131448 9120
rect 131868 8974 131896 10270
rect 132314 10231 132370 10240
rect 131120 8968 131172 8974
rect 131120 8910 131172 8916
rect 131856 8968 131908 8974
rect 131856 8910 131908 8916
rect 130568 8424 130620 8430
rect 130568 8366 130620 8372
rect 130290 7440 130346 7449
rect 130290 7375 130346 7384
rect 129108 6886 129228 6914
rect 129476 6886 129596 6914
rect 128636 2440 128688 2446
rect 128636 2382 128688 2388
rect 128360 2304 128412 2310
rect 128360 2246 128412 2252
rect 128372 1465 128400 2246
rect 128452 1896 128504 1902
rect 128452 1838 128504 1844
rect 128358 1456 128414 1465
rect 128358 1391 128414 1400
rect 128464 1358 128492 1838
rect 128648 1358 128676 2382
rect 129200 2038 129228 6886
rect 129568 2038 129596 6886
rect 130304 6390 130332 7375
rect 130200 6384 130252 6390
rect 130200 6326 130252 6332
rect 130292 6384 130344 6390
rect 130292 6326 130344 6332
rect 129924 6316 129976 6322
rect 129924 6258 129976 6264
rect 129936 5710 129964 6258
rect 130212 5953 130240 6326
rect 130198 5944 130254 5953
rect 130198 5879 130254 5888
rect 130212 5778 130240 5879
rect 130200 5772 130252 5778
rect 130200 5714 130252 5720
rect 129924 5704 129976 5710
rect 129924 5646 129976 5652
rect 129936 4486 129964 5646
rect 129924 4480 129976 4486
rect 129924 4422 129976 4428
rect 129648 2440 129700 2446
rect 129648 2382 129700 2388
rect 129660 2106 129688 2382
rect 130016 2304 130068 2310
rect 130016 2246 130068 2252
rect 129648 2100 129700 2106
rect 129648 2042 129700 2048
rect 129188 2032 129240 2038
rect 129188 1974 129240 1980
rect 129556 2032 129608 2038
rect 129556 1974 129608 1980
rect 129556 1896 129608 1902
rect 129740 1896 129792 1902
rect 129608 1856 129740 1884
rect 129556 1838 129608 1844
rect 129740 1838 129792 1844
rect 129096 1760 129148 1766
rect 129096 1702 129148 1708
rect 129108 1358 129136 1702
rect 128268 1352 128320 1358
rect 128268 1294 128320 1300
rect 128452 1352 128504 1358
rect 128452 1294 128504 1300
rect 128636 1352 128688 1358
rect 128636 1294 128688 1300
rect 129096 1352 129148 1358
rect 129096 1294 129148 1300
rect 129280 1216 129332 1222
rect 129280 1158 129332 1164
rect 129292 649 129320 1158
rect 130028 649 130056 2246
rect 130580 1970 130608 8366
rect 131132 1970 131160 8910
rect 131672 2440 131724 2446
rect 131672 2382 131724 2388
rect 131580 2304 131632 2310
rect 131580 2246 131632 2252
rect 130568 1964 130620 1970
rect 130568 1906 130620 1912
rect 131120 1964 131172 1970
rect 131120 1906 131172 1912
rect 130660 1760 130712 1766
rect 130660 1702 130712 1708
rect 130672 1358 130700 1702
rect 130660 1352 130712 1358
rect 130660 1294 130712 1300
rect 130844 1216 130896 1222
rect 130844 1158 130896 1164
rect 124770 640 124826 649
rect 124770 575 124826 584
rect 125322 640 125378 649
rect 125322 575 125378 584
rect 126334 640 126390 649
rect 126334 575 126390 584
rect 126794 640 126850 649
rect 126794 575 126850 584
rect 127806 640 127862 649
rect 127806 575 127862 584
rect 129278 640 129334 649
rect 129278 575 129334 584
rect 130014 640 130070 649
rect 130014 575 130070 584
rect 120446 504 120502 513
rect 120446 439 120502 448
rect 124034 504 124090 513
rect 124034 439 124090 448
rect 130856 377 130884 1158
rect 131592 649 131620 2246
rect 131684 2106 131712 2382
rect 131672 2100 131724 2106
rect 131672 2042 131724 2048
rect 131868 1970 131896 8910
rect 132132 8832 132184 8838
rect 132132 8774 132184 8780
rect 132144 8498 132172 8774
rect 132328 8634 132356 10231
rect 132316 8628 132368 8634
rect 132316 8570 132368 8576
rect 132880 8498 132908 10746
rect 133708 10606 133736 10746
rect 133696 10600 133748 10606
rect 133696 10542 133748 10548
rect 133788 10532 133840 10538
rect 133788 10474 133840 10480
rect 133050 10296 133106 10305
rect 132960 10260 133012 10266
rect 133050 10231 133106 10240
rect 133510 10296 133566 10305
rect 133800 10266 133828 10474
rect 148414 10432 148470 10441
rect 133972 10396 134024 10402
rect 148414 10367 148470 10376
rect 151728 10396 151780 10402
rect 133972 10338 134024 10344
rect 133510 10231 133566 10240
rect 133788 10260 133840 10266
rect 132960 10202 133012 10208
rect 132972 8974 133000 10202
rect 132960 8968 133012 8974
rect 132960 8910 133012 8916
rect 132132 8492 132184 8498
rect 132868 8492 132920 8498
rect 132132 8434 132184 8440
rect 132788 8452 132868 8480
rect 131856 1964 131908 1970
rect 131856 1906 131908 1912
rect 132592 1760 132644 1766
rect 132592 1702 132644 1708
rect 132604 1358 132632 1702
rect 132788 1358 132816 8452
rect 132868 8434 132920 8440
rect 132868 8288 132920 8294
rect 132868 8230 132920 8236
rect 132880 7886 132908 8230
rect 132868 7880 132920 7886
rect 132868 7822 132920 7828
rect 132972 6914 133000 8910
rect 133064 8090 133092 10231
rect 133524 9722 133552 10231
rect 133788 10202 133840 10208
rect 133512 9716 133564 9722
rect 133512 9658 133564 9664
rect 133420 9580 133472 9586
rect 133420 9522 133472 9528
rect 133432 9110 133460 9522
rect 133984 9110 134012 10338
rect 134246 10296 134302 10305
rect 134246 10231 134302 10240
rect 134890 10296 134946 10305
rect 134890 10231 134946 10240
rect 138754 10296 138810 10305
rect 138754 10231 138810 10240
rect 143262 10296 143318 10305
rect 143262 10231 143318 10240
rect 134260 9722 134288 10231
rect 134248 9716 134300 9722
rect 134248 9658 134300 9664
rect 134248 9580 134300 9586
rect 134248 9522 134300 9528
rect 134260 9110 134288 9522
rect 134904 9110 134932 10231
rect 136143 9820 136451 9829
rect 136143 9818 136149 9820
rect 136205 9818 136229 9820
rect 136285 9818 136309 9820
rect 136365 9818 136389 9820
rect 136445 9818 136451 9820
rect 136205 9766 136207 9818
rect 136387 9766 136389 9818
rect 136143 9764 136149 9766
rect 136205 9764 136229 9766
rect 136285 9764 136309 9766
rect 136365 9764 136389 9766
rect 136445 9764 136451 9766
rect 136143 9755 136451 9764
rect 137284 9716 137336 9722
rect 137284 9658 137336 9664
rect 137296 9382 137324 9658
rect 137374 9616 137430 9625
rect 138768 9586 138796 10231
rect 138846 10160 138902 10169
rect 138846 10095 138902 10104
rect 140686 10160 140742 10169
rect 140686 10095 140742 10104
rect 141330 10160 141386 10169
rect 141330 10095 141386 10104
rect 141974 10160 142030 10169
rect 141974 10095 142030 10104
rect 138860 9586 138888 10095
rect 139766 9888 139822 9897
rect 139766 9823 139822 9832
rect 137374 9551 137376 9560
rect 137428 9551 137430 9560
rect 138756 9580 138808 9586
rect 137376 9522 137428 9528
rect 138756 9522 138808 9528
rect 138848 9580 138900 9586
rect 138848 9522 138900 9528
rect 137284 9376 137336 9382
rect 137284 9318 137336 9324
rect 137744 9376 137796 9382
rect 137744 9318 137796 9324
rect 138112 9376 138164 9382
rect 138112 9318 138164 9324
rect 133420 9104 133472 9110
rect 133420 9046 133472 9052
rect 133972 9104 134024 9110
rect 133972 9046 134024 9052
rect 134248 9104 134300 9110
rect 134248 9046 134300 9052
rect 134892 9104 134944 9110
rect 134892 9046 134944 9052
rect 133984 8974 134012 9046
rect 133144 8968 133196 8974
rect 133144 8910 133196 8916
rect 133972 8968 134024 8974
rect 133972 8910 134024 8916
rect 134524 8968 134576 8974
rect 134524 8910 134576 8916
rect 133156 8498 133184 8910
rect 133144 8492 133196 8498
rect 133144 8434 133196 8440
rect 133052 8084 133104 8090
rect 133052 8026 133104 8032
rect 133984 6914 134012 8910
rect 134248 8832 134300 8838
rect 134248 8774 134300 8780
rect 134260 8498 134288 8774
rect 134536 8634 134564 8910
rect 137284 8900 137336 8906
rect 137284 8842 137336 8848
rect 137376 8900 137428 8906
rect 137376 8842 137428 8848
rect 136143 8732 136451 8741
rect 136143 8730 136149 8732
rect 136205 8730 136229 8732
rect 136285 8730 136309 8732
rect 136365 8730 136389 8732
rect 136445 8730 136451 8732
rect 136205 8678 136207 8730
rect 136387 8678 136389 8730
rect 136143 8676 136149 8678
rect 136205 8676 136229 8678
rect 136285 8676 136309 8678
rect 136365 8676 136389 8678
rect 136445 8676 136451 8678
rect 136143 8667 136451 8676
rect 137296 8634 137324 8842
rect 134524 8628 134576 8634
rect 134524 8570 134576 8576
rect 137284 8628 137336 8634
rect 137284 8570 137336 8576
rect 134248 8492 134300 8498
rect 134248 8434 134300 8440
rect 137388 8362 137416 8842
rect 137376 8356 137428 8362
rect 137376 8298 137428 8304
rect 136143 7644 136451 7653
rect 136143 7642 136149 7644
rect 136205 7642 136229 7644
rect 136285 7642 136309 7644
rect 136365 7642 136389 7644
rect 136445 7642 136451 7644
rect 136205 7590 136207 7642
rect 136387 7590 136389 7642
rect 136143 7588 136149 7590
rect 136205 7588 136229 7590
rect 136285 7588 136309 7590
rect 136365 7588 136389 7590
rect 136445 7588 136451 7590
rect 136143 7579 136451 7588
rect 132972 6886 133092 6914
rect 132960 2304 133012 2310
rect 132960 2246 133012 2252
rect 132592 1352 132644 1358
rect 132592 1294 132644 1300
rect 132776 1352 132828 1358
rect 132776 1294 132828 1300
rect 132132 1216 132184 1222
rect 132132 1158 132184 1164
rect 132144 649 132172 1158
rect 132972 649 133000 2246
rect 133064 1970 133092 6886
rect 133892 6886 134012 6914
rect 133328 2440 133380 2446
rect 133328 2382 133380 2388
rect 133604 2440 133656 2446
rect 133604 2382 133656 2388
rect 133236 2372 133288 2378
rect 133236 2314 133288 2320
rect 133052 1964 133104 1970
rect 133052 1906 133104 1912
rect 133144 1896 133196 1902
rect 133144 1838 133196 1844
rect 133156 1358 133184 1838
rect 133248 1494 133276 2314
rect 133340 1494 133368 2382
rect 133616 2038 133644 2382
rect 133696 2304 133748 2310
rect 133696 2246 133748 2252
rect 133604 2032 133656 2038
rect 133604 1974 133656 1980
rect 133236 1488 133288 1494
rect 133236 1430 133288 1436
rect 133328 1488 133380 1494
rect 133328 1430 133380 1436
rect 133144 1352 133196 1358
rect 133144 1294 133196 1300
rect 133708 649 133736 2246
rect 133892 1358 133920 6886
rect 136143 6556 136451 6565
rect 136143 6554 136149 6556
rect 136205 6554 136229 6556
rect 136285 6554 136309 6556
rect 136365 6554 136389 6556
rect 136445 6554 136451 6556
rect 136205 6502 136207 6554
rect 136387 6502 136389 6554
rect 136143 6500 136149 6502
rect 136205 6500 136229 6502
rect 136285 6500 136309 6502
rect 136365 6500 136389 6502
rect 136445 6500 136451 6502
rect 136143 6491 136451 6500
rect 136143 5468 136451 5477
rect 136143 5466 136149 5468
rect 136205 5466 136229 5468
rect 136285 5466 136309 5468
rect 136365 5466 136389 5468
rect 136445 5466 136451 5468
rect 136205 5414 136207 5466
rect 136387 5414 136389 5466
rect 136143 5412 136149 5414
rect 136205 5412 136229 5414
rect 136285 5412 136309 5414
rect 136365 5412 136389 5414
rect 136445 5412 136451 5414
rect 136143 5403 136451 5412
rect 136143 4380 136451 4389
rect 136143 4378 136149 4380
rect 136205 4378 136229 4380
rect 136285 4378 136309 4380
rect 136365 4378 136389 4380
rect 136445 4378 136451 4380
rect 136205 4326 136207 4378
rect 136387 4326 136389 4378
rect 136143 4324 136149 4326
rect 136205 4324 136229 4326
rect 136285 4324 136309 4326
rect 136365 4324 136389 4326
rect 136445 4324 136451 4326
rect 136143 4315 136451 4324
rect 136143 3292 136451 3301
rect 136143 3290 136149 3292
rect 136205 3290 136229 3292
rect 136285 3290 136309 3292
rect 136365 3290 136389 3292
rect 136445 3290 136451 3292
rect 136205 3238 136207 3290
rect 136387 3238 136389 3290
rect 136143 3236 136149 3238
rect 136205 3236 136229 3238
rect 136285 3236 136309 3238
rect 136365 3236 136389 3238
rect 136445 3236 136451 3238
rect 136143 3227 136451 3236
rect 137756 3058 137784 9318
rect 137744 3052 137796 3058
rect 137744 2994 137796 3000
rect 137928 2984 137980 2990
rect 137928 2926 137980 2932
rect 134340 2440 134392 2446
rect 134340 2382 134392 2388
rect 134064 1896 134116 1902
rect 134064 1838 134116 1844
rect 134076 1358 134104 1838
rect 134352 1494 134380 2382
rect 134432 2304 134484 2310
rect 134432 2246 134484 2252
rect 134984 2304 135036 2310
rect 134984 2246 135036 2252
rect 134340 1488 134392 1494
rect 134340 1430 134392 1436
rect 133880 1352 133932 1358
rect 133880 1294 133932 1300
rect 134064 1352 134116 1358
rect 134064 1294 134116 1300
rect 134444 649 134472 2246
rect 134996 2038 135024 2246
rect 136143 2204 136451 2213
rect 136143 2202 136149 2204
rect 136205 2202 136229 2204
rect 136285 2202 136309 2204
rect 136365 2202 136389 2204
rect 136445 2202 136451 2204
rect 136205 2150 136207 2202
rect 136387 2150 136389 2202
rect 136143 2148 136149 2150
rect 136205 2148 136229 2150
rect 136285 2148 136309 2150
rect 136365 2148 136389 2150
rect 136445 2148 136451 2150
rect 136143 2139 136451 2148
rect 134984 2032 135036 2038
rect 134984 1974 135036 1980
rect 135260 1760 135312 1766
rect 135260 1702 135312 1708
rect 135272 1465 135300 1702
rect 135258 1456 135314 1465
rect 135258 1391 135314 1400
rect 137940 1222 137968 2926
rect 138124 1970 138152 9318
rect 139780 8974 139808 9823
rect 140700 9586 140728 10095
rect 141344 9586 141372 10095
rect 141988 9586 142016 10095
rect 143276 9586 143304 10231
rect 143354 10160 143410 10169
rect 143354 10095 143410 10104
rect 144550 10160 144606 10169
rect 144550 10095 144606 10104
rect 145838 10160 145894 10169
rect 145838 10095 145894 10104
rect 146206 10160 146262 10169
rect 146206 10095 146262 10104
rect 147126 10160 147182 10169
rect 147126 10095 147182 10104
rect 143368 9586 143396 10095
rect 144564 9586 144592 10095
rect 144734 9888 144790 9897
rect 144734 9823 144790 9832
rect 140688 9580 140740 9586
rect 140688 9522 140740 9528
rect 141332 9580 141384 9586
rect 141332 9522 141384 9528
rect 141976 9580 142028 9586
rect 141976 9522 142028 9528
rect 143264 9580 143316 9586
rect 143264 9522 143316 9528
rect 143356 9580 143408 9586
rect 143356 9522 143408 9528
rect 144552 9580 144604 9586
rect 144552 9522 144604 9528
rect 142712 9444 142764 9450
rect 142712 9386 142764 9392
rect 140504 9376 140556 9382
rect 140504 9318 140556 9324
rect 139768 8968 139820 8974
rect 139768 8910 139820 8916
rect 140412 8832 140464 8838
rect 140412 8774 140464 8780
rect 138664 7880 138716 7886
rect 138664 7822 138716 7828
rect 138572 3392 138624 3398
rect 138572 3334 138624 3340
rect 138388 2916 138440 2922
rect 138388 2858 138440 2864
rect 138112 1964 138164 1970
rect 138112 1906 138164 1912
rect 138400 1902 138428 2858
rect 138584 2417 138612 3334
rect 138676 3058 138704 7822
rect 139308 4820 139360 4826
rect 139308 4762 139360 4768
rect 139320 4078 139348 4762
rect 139308 4072 139360 4078
rect 139308 4014 139360 4020
rect 138940 3528 138992 3534
rect 138940 3470 138992 3476
rect 138952 3194 138980 3470
rect 139124 3460 139176 3466
rect 139124 3402 139176 3408
rect 138940 3188 138992 3194
rect 138940 3130 138992 3136
rect 138664 3052 138716 3058
rect 138664 2994 138716 3000
rect 139136 2990 139164 3402
rect 138756 2984 138808 2990
rect 138940 2984 138992 2990
rect 138756 2926 138808 2932
rect 138860 2944 138940 2972
rect 138768 2774 138796 2926
rect 138676 2746 138796 2774
rect 138570 2408 138626 2417
rect 138570 2343 138626 2352
rect 138296 1896 138348 1902
rect 138296 1838 138348 1844
rect 138388 1896 138440 1902
rect 138388 1838 138440 1844
rect 138308 1494 138336 1838
rect 138020 1488 138072 1494
rect 138018 1456 138020 1465
rect 138296 1488 138348 1494
rect 138072 1456 138074 1465
rect 138296 1430 138348 1436
rect 138018 1391 138074 1400
rect 137928 1216 137980 1222
rect 137928 1158 137980 1164
rect 136143 1116 136451 1125
rect 136143 1114 136149 1116
rect 136205 1114 136229 1116
rect 136285 1114 136309 1116
rect 136365 1114 136389 1116
rect 136445 1114 136451 1116
rect 136205 1062 136207 1114
rect 136387 1062 136389 1114
rect 136143 1060 136149 1062
rect 136205 1060 136229 1062
rect 136285 1060 136309 1062
rect 136365 1060 136389 1062
rect 136445 1060 136451 1062
rect 136143 1051 136451 1060
rect 131578 640 131634 649
rect 131578 575 131634 584
rect 132130 640 132186 649
rect 132130 575 132186 584
rect 132958 640 133014 649
rect 132958 575 133014 584
rect 133694 640 133750 649
rect 133694 575 133750 584
rect 134430 640 134486 649
rect 138676 610 138704 2746
rect 138860 2145 138888 2944
rect 138940 2926 138992 2932
rect 139124 2984 139176 2990
rect 139124 2926 139176 2932
rect 139136 2514 139164 2926
rect 139124 2508 139176 2514
rect 139124 2450 139176 2456
rect 139030 2408 139086 2417
rect 139030 2343 139086 2352
rect 139952 2372 140004 2378
rect 138846 2136 138902 2145
rect 138846 2071 138902 2080
rect 138860 1902 138888 2071
rect 139044 1970 139072 2343
rect 139952 2314 140004 2320
rect 139964 2038 139992 2314
rect 139952 2032 140004 2038
rect 139214 2000 139270 2009
rect 139032 1964 139084 1970
rect 139952 1974 140004 1980
rect 140424 1970 140452 8774
rect 140516 6866 140544 9318
rect 141700 7948 141752 7954
rect 141700 7890 141752 7896
rect 141608 7812 141660 7818
rect 141608 7754 141660 7760
rect 141620 6866 141648 7754
rect 141712 6866 141740 7890
rect 140504 6860 140556 6866
rect 140504 6802 140556 6808
rect 141332 6860 141384 6866
rect 141332 6802 141384 6808
rect 141608 6860 141660 6866
rect 141608 6802 141660 6808
rect 141700 6860 141752 6866
rect 141700 6802 141752 6808
rect 140872 6792 140924 6798
rect 140872 6734 140924 6740
rect 140688 3460 140740 3466
rect 140688 3402 140740 3408
rect 140700 2961 140728 3402
rect 140686 2952 140742 2961
rect 140686 2887 140742 2896
rect 140780 2916 140832 2922
rect 140780 2858 140832 2864
rect 139214 1935 139216 1944
rect 139032 1906 139084 1912
rect 139268 1935 139270 1944
rect 140412 1964 140464 1970
rect 139216 1906 139268 1912
rect 140412 1906 140464 1912
rect 138848 1896 138900 1902
rect 138848 1838 138900 1844
rect 140688 1896 140740 1902
rect 140688 1838 140740 1844
rect 140700 1494 140728 1838
rect 140792 1766 140820 2858
rect 140780 1760 140832 1766
rect 140780 1702 140832 1708
rect 140688 1488 140740 1494
rect 140688 1430 140740 1436
rect 138756 1352 138808 1358
rect 138756 1294 138808 1300
rect 138848 1352 138900 1358
rect 138848 1294 138900 1300
rect 140688 1352 140740 1358
rect 140780 1352 140832 1358
rect 140688 1294 140740 1300
rect 140778 1320 140780 1329
rect 140832 1320 140834 1329
rect 138768 649 138796 1294
rect 138860 785 138888 1294
rect 138846 776 138902 785
rect 138846 711 138902 720
rect 138754 640 138810 649
rect 134430 575 134486 584
rect 138664 604 138716 610
rect 138754 575 138810 584
rect 138664 546 138716 552
rect 140700 513 140728 1294
rect 140778 1255 140834 1264
rect 140884 1222 140912 6734
rect 141344 6390 141372 6802
rect 141712 6662 141740 6802
rect 141884 6792 141936 6798
rect 141884 6734 141936 6740
rect 141700 6656 141752 6662
rect 141700 6598 141752 6604
rect 141332 6384 141384 6390
rect 141332 6326 141384 6332
rect 141896 4162 141924 6734
rect 142620 6180 142672 6186
rect 142620 6122 142672 6128
rect 142632 5642 142660 6122
rect 142620 5636 142672 5642
rect 142620 5578 142672 5584
rect 142160 4548 142212 4554
rect 142160 4490 142212 4496
rect 141712 4134 141924 4162
rect 141424 3936 141476 3942
rect 141424 3878 141476 3884
rect 141436 3602 141464 3878
rect 141424 3596 141476 3602
rect 141424 3538 141476 3544
rect 141148 2508 141200 2514
rect 141148 2450 141200 2456
rect 141160 1834 141188 2450
rect 141332 2304 141384 2310
rect 141332 2246 141384 2252
rect 141148 1828 141200 1834
rect 141148 1770 141200 1776
rect 140872 1216 140924 1222
rect 140872 1158 140924 1164
rect 141344 882 141372 2246
rect 141712 2145 141740 4134
rect 142172 4078 142200 4490
rect 142436 4480 142488 4486
rect 142436 4422 142488 4428
rect 142448 4282 142476 4422
rect 142436 4276 142488 4282
rect 142436 4218 142488 4224
rect 141792 4072 141844 4078
rect 141792 4014 141844 4020
rect 142160 4072 142212 4078
rect 142160 4014 142212 4020
rect 141804 3194 141832 4014
rect 141792 3188 141844 3194
rect 141792 3130 141844 3136
rect 142172 3126 142200 4014
rect 142160 3120 142212 3126
rect 142160 3062 142212 3068
rect 141884 3052 141936 3058
rect 141884 2994 141936 3000
rect 141698 2136 141754 2145
rect 141698 2071 141754 2080
rect 141712 1970 141740 2071
rect 141424 1964 141476 1970
rect 141424 1906 141476 1912
rect 141700 1964 141752 1970
rect 141700 1906 141752 1912
rect 141436 1873 141464 1906
rect 141516 1896 141568 1902
rect 141422 1864 141478 1873
rect 141516 1838 141568 1844
rect 141422 1799 141478 1808
rect 141528 1018 141556 1838
rect 141896 1222 141924 2994
rect 142724 2990 142752 9386
rect 142988 9376 143040 9382
rect 142988 9318 143040 9324
rect 143264 9376 143316 9382
rect 143264 9318 143316 9324
rect 142804 5364 142856 5370
rect 142804 5306 142856 5312
rect 142816 4758 142844 5306
rect 142804 4752 142856 4758
rect 142804 4694 142856 4700
rect 143000 3602 143028 9318
rect 143080 6656 143132 6662
rect 143080 6598 143132 6604
rect 143092 5778 143120 6598
rect 143080 5772 143132 5778
rect 143080 5714 143132 5720
rect 142988 3596 143040 3602
rect 142988 3538 143040 3544
rect 143172 3528 143224 3534
rect 143172 3470 143224 3476
rect 143184 3108 143212 3470
rect 143092 3080 143212 3108
rect 142712 2984 142764 2990
rect 142712 2926 142764 2932
rect 142712 2848 142764 2854
rect 142712 2790 142764 2796
rect 141976 1352 142028 1358
rect 141976 1294 142028 1300
rect 142068 1352 142120 1358
rect 142068 1294 142120 1300
rect 141884 1216 141936 1222
rect 141884 1158 141936 1164
rect 141516 1012 141568 1018
rect 141516 954 141568 960
rect 141332 876 141384 882
rect 141332 818 141384 824
rect 141988 785 142016 1294
rect 141974 776 142030 785
rect 141974 711 142030 720
rect 142080 649 142108 1294
rect 142724 814 142752 2790
rect 142804 2440 142856 2446
rect 142804 2382 142856 2388
rect 142816 1834 142844 2382
rect 142988 1964 143040 1970
rect 142988 1906 143040 1912
rect 142804 1828 142856 1834
rect 142804 1770 142856 1776
rect 143000 1057 143028 1906
rect 143092 1222 143120 3080
rect 143276 2774 143304 9318
rect 144748 8974 144776 9823
rect 145852 9586 145880 10095
rect 146220 9586 146248 10095
rect 146392 9648 146444 9654
rect 146392 9590 146444 9596
rect 145840 9580 145892 9586
rect 145840 9522 145892 9528
rect 146208 9580 146260 9586
rect 146208 9522 146260 9528
rect 145380 9444 145432 9450
rect 145380 9386 145432 9392
rect 145840 9444 145892 9450
rect 145840 9386 145892 9392
rect 144736 8968 144788 8974
rect 144736 8910 144788 8916
rect 144000 7744 144052 7750
rect 144000 7686 144052 7692
rect 143448 6384 143500 6390
rect 143448 6326 143500 6332
rect 143356 6248 143408 6254
rect 143356 6190 143408 6196
rect 143368 5778 143396 6190
rect 143356 5772 143408 5778
rect 143356 5714 143408 5720
rect 143368 4554 143396 5714
rect 143356 4548 143408 4554
rect 143356 4490 143408 4496
rect 143460 3670 143488 6326
rect 143540 5772 143592 5778
rect 143540 5714 143592 5720
rect 143552 5681 143580 5714
rect 143538 5672 143594 5681
rect 143538 5607 143540 5616
rect 143592 5607 143594 5616
rect 143540 5578 143592 5584
rect 143448 3664 143500 3670
rect 143448 3606 143500 3612
rect 143460 2990 143488 3606
rect 144012 3602 144040 7686
rect 144550 7576 144606 7585
rect 144550 7511 144606 7520
rect 144460 6452 144512 6458
rect 144460 6394 144512 6400
rect 144472 5778 144500 6394
rect 144460 5772 144512 5778
rect 144460 5714 144512 5720
rect 144564 5114 144592 7511
rect 145196 5704 145248 5710
rect 145196 5646 145248 5652
rect 144472 5086 144592 5114
rect 144274 3632 144330 3641
rect 144000 3596 144052 3602
rect 144274 3567 144330 3576
rect 144000 3538 144052 3544
rect 144288 3534 144316 3567
rect 144276 3528 144328 3534
rect 144276 3470 144328 3476
rect 143816 3392 143868 3398
rect 143816 3334 143868 3340
rect 143722 3088 143778 3097
rect 143722 3023 143724 3032
rect 143776 3023 143778 3032
rect 143724 2994 143776 3000
rect 143448 2984 143500 2990
rect 143500 2944 143672 2972
rect 143448 2926 143500 2932
rect 143644 2802 143672 2944
rect 143644 2774 143764 2802
rect 143184 2746 143304 2774
rect 143184 2514 143212 2746
rect 143736 2582 143764 2774
rect 143724 2576 143776 2582
rect 143724 2518 143776 2524
rect 143172 2508 143224 2514
rect 143172 2450 143224 2456
rect 143172 1896 143224 1902
rect 143170 1864 143172 1873
rect 143224 1864 143226 1873
rect 143170 1799 143226 1808
rect 143540 1352 143592 1358
rect 143540 1294 143592 1300
rect 143080 1216 143132 1222
rect 143080 1158 143132 1164
rect 142986 1048 143042 1057
rect 142986 983 143042 992
rect 142712 808 142764 814
rect 143552 785 143580 1294
rect 143828 1222 143856 3334
rect 143908 2984 143960 2990
rect 143908 2926 143960 2932
rect 144000 2984 144052 2990
rect 144000 2926 144052 2932
rect 143816 1216 143868 1222
rect 143816 1158 143868 1164
rect 142712 750 142764 756
rect 143538 776 143594 785
rect 143538 711 143594 720
rect 143920 678 143948 2926
rect 144012 2530 144040 2926
rect 144288 2530 144316 3470
rect 144368 2984 144420 2990
rect 144368 2926 144420 2932
rect 144012 2502 144316 2530
rect 144012 2145 144040 2502
rect 144288 2446 144316 2502
rect 144184 2440 144236 2446
rect 144184 2382 144236 2388
rect 144276 2440 144328 2446
rect 144276 2382 144328 2388
rect 143998 2136 144054 2145
rect 143998 2071 144054 2080
rect 144196 1494 144224 2382
rect 144184 1488 144236 1494
rect 144184 1430 144236 1436
rect 144380 1222 144408 2926
rect 144472 2514 144500 5086
rect 144828 4684 144880 4690
rect 144828 4626 144880 4632
rect 144840 3670 144868 4626
rect 145208 4554 145236 5646
rect 145196 4548 145248 4554
rect 145196 4490 145248 4496
rect 144736 3664 144788 3670
rect 144734 3632 144736 3641
rect 144828 3664 144880 3670
rect 144788 3632 144790 3641
rect 144644 3596 144696 3602
rect 144828 3606 144880 3612
rect 145392 3602 145420 9386
rect 145564 9376 145616 9382
rect 145564 9318 145616 9324
rect 144734 3567 144790 3576
rect 145380 3596 145432 3602
rect 144644 3538 144696 3544
rect 145380 3538 145432 3544
rect 144460 2508 144512 2514
rect 144460 2450 144512 2456
rect 144656 2145 144684 3538
rect 144828 3460 144880 3466
rect 144828 3402 144880 3408
rect 144840 3194 144868 3402
rect 144828 3188 144880 3194
rect 144828 3130 144880 3136
rect 144840 2854 144868 3130
rect 145576 2990 145604 9318
rect 145852 6866 145880 9386
rect 146208 9376 146260 9382
rect 146208 9318 146260 9324
rect 146300 9376 146352 9382
rect 146300 9318 146352 9324
rect 146116 7268 146168 7274
rect 146116 7210 146168 7216
rect 145840 6860 145892 6866
rect 145840 6802 145892 6808
rect 145656 4072 145708 4078
rect 145656 4014 145708 4020
rect 145564 2984 145616 2990
rect 145564 2926 145616 2932
rect 144828 2848 144880 2854
rect 144828 2790 144880 2796
rect 145668 2582 145696 4014
rect 145656 2576 145708 2582
rect 145656 2518 145708 2524
rect 144642 2136 144698 2145
rect 144642 2071 144698 2080
rect 144920 1964 144972 1970
rect 144920 1906 144972 1912
rect 144932 1465 144960 1906
rect 144918 1456 144974 1465
rect 144918 1391 144974 1400
rect 144552 1352 144604 1358
rect 144552 1294 144604 1300
rect 145840 1352 145892 1358
rect 145840 1294 145892 1300
rect 144368 1216 144420 1222
rect 144368 1158 144420 1164
rect 144564 785 144592 1294
rect 145656 1216 145708 1222
rect 145656 1158 145708 1164
rect 145668 950 145696 1158
rect 145656 944 145708 950
rect 145656 886 145708 892
rect 145852 785 145880 1294
rect 146128 1222 146156 7210
rect 146220 2514 146248 9318
rect 146312 7546 146340 9318
rect 146404 7750 146432 9590
rect 147140 9586 147168 10095
rect 148428 9586 148456 10367
rect 151728 10338 151780 10344
rect 149060 10328 149112 10334
rect 149060 10270 149112 10276
rect 148506 10160 148562 10169
rect 148506 10095 148562 10104
rect 148520 9586 148548 10095
rect 147128 9580 147180 9586
rect 147128 9522 147180 9528
rect 148416 9580 148468 9586
rect 148416 9522 148468 9528
rect 148508 9580 148560 9586
rect 148508 9522 148560 9528
rect 148232 9376 148284 9382
rect 148232 9318 148284 9324
rect 147772 8832 147824 8838
rect 147772 8774 147824 8780
rect 146852 8288 146904 8294
rect 146852 8230 146904 8236
rect 146496 7818 146708 7834
rect 146484 7812 146720 7818
rect 146536 7806 146668 7812
rect 146484 7754 146536 7760
rect 146668 7754 146720 7760
rect 146392 7744 146444 7750
rect 146392 7686 146444 7692
rect 146574 7712 146630 7721
rect 146574 7647 146630 7656
rect 146300 7540 146352 7546
rect 146300 7482 146352 7488
rect 146300 7268 146352 7274
rect 146300 7210 146352 7216
rect 146312 6934 146340 7210
rect 146300 6928 146352 6934
rect 146300 6870 146352 6876
rect 146392 6860 146444 6866
rect 146392 6802 146444 6808
rect 146298 5400 146354 5409
rect 146298 5335 146354 5344
rect 146312 3534 146340 5335
rect 146300 3528 146352 3534
rect 146300 3470 146352 3476
rect 146208 2508 146260 2514
rect 146208 2450 146260 2456
rect 146208 1352 146260 1358
rect 146208 1294 146260 1300
rect 146116 1216 146168 1222
rect 146116 1158 146168 1164
rect 146220 785 146248 1294
rect 146404 1222 146432 6802
rect 146484 3528 146536 3534
rect 146484 3470 146536 3476
rect 146496 1766 146524 3470
rect 146588 3058 146616 7647
rect 146760 7540 146812 7546
rect 146760 7482 146812 7488
rect 146772 7410 146800 7482
rect 146760 7404 146812 7410
rect 146760 7346 146812 7352
rect 146864 7290 146892 8230
rect 146772 7262 146892 7290
rect 147036 7336 147088 7342
rect 147036 7278 147088 7284
rect 146772 6798 146800 7262
rect 147048 6798 147076 7278
rect 147496 7200 147548 7206
rect 147496 7142 147548 7148
rect 146760 6792 146812 6798
rect 146760 6734 146812 6740
rect 146944 6792 146996 6798
rect 146944 6734 146996 6740
rect 147036 6792 147088 6798
rect 147036 6734 147088 6740
rect 146852 6656 146904 6662
rect 146852 6598 146904 6604
rect 146864 3398 146892 6598
rect 146852 3392 146904 3398
rect 146852 3334 146904 3340
rect 146864 3058 146892 3334
rect 146576 3052 146628 3058
rect 146576 2994 146628 3000
rect 146852 3052 146904 3058
rect 146852 2994 146904 3000
rect 146760 2984 146812 2990
rect 146760 2926 146812 2932
rect 146484 1760 146536 1766
rect 146484 1702 146536 1708
rect 146392 1216 146444 1222
rect 146392 1158 146444 1164
rect 144550 776 144606 785
rect 144550 711 144606 720
rect 145838 776 145894 785
rect 145838 711 145894 720
rect 146206 776 146262 785
rect 146772 746 146800 2926
rect 146956 2774 146984 6734
rect 147048 6662 147076 6734
rect 147036 6656 147088 6662
rect 147036 6598 147088 6604
rect 147508 6390 147536 7142
rect 147588 6860 147640 6866
rect 147588 6802 147640 6808
rect 147600 6644 147628 6802
rect 147600 6616 147720 6644
rect 147692 6390 147720 6616
rect 147496 6384 147548 6390
rect 147496 6326 147548 6332
rect 147680 6384 147732 6390
rect 147680 6326 147732 6332
rect 147588 5772 147640 5778
rect 147588 5714 147640 5720
rect 147600 5574 147628 5714
rect 147588 5568 147640 5574
rect 147588 5510 147640 5516
rect 147496 4208 147548 4214
rect 147496 4150 147548 4156
rect 147508 3942 147536 4150
rect 147496 3936 147548 3942
rect 147496 3878 147548 3884
rect 147496 3528 147548 3534
rect 147496 3470 147548 3476
rect 147508 3194 147536 3470
rect 147496 3188 147548 3194
rect 147496 3130 147548 3136
rect 147784 3058 147812 8774
rect 148244 6866 148272 9318
rect 148692 8492 148744 8498
rect 148692 8434 148744 8440
rect 148232 6860 148284 6866
rect 148232 6802 148284 6808
rect 148324 6792 148376 6798
rect 148324 6734 148376 6740
rect 148232 6656 148284 6662
rect 148232 6598 148284 6604
rect 148048 6452 148100 6458
rect 148048 6394 148100 6400
rect 148060 5710 148088 6394
rect 148140 6248 148192 6254
rect 148138 6216 148140 6225
rect 148192 6216 148194 6225
rect 148138 6151 148194 6160
rect 148244 5778 148272 6598
rect 148232 5772 148284 5778
rect 148232 5714 148284 5720
rect 148048 5704 148100 5710
rect 148048 5646 148100 5652
rect 148140 5636 148192 5642
rect 148140 5578 148192 5584
rect 148152 4078 148180 5578
rect 147956 4072 148008 4078
rect 147956 4014 148008 4020
rect 148140 4072 148192 4078
rect 148140 4014 148192 4020
rect 147968 3670 147996 4014
rect 147956 3664 148008 3670
rect 147956 3606 148008 3612
rect 148048 3664 148100 3670
rect 148048 3606 148100 3612
rect 148060 3126 148088 3606
rect 148152 3194 148180 4014
rect 148140 3188 148192 3194
rect 148140 3130 148192 3136
rect 148048 3120 148100 3126
rect 148048 3062 148100 3068
rect 147772 3052 147824 3058
rect 147772 2994 147824 3000
rect 148140 2984 148192 2990
rect 148140 2926 148192 2932
rect 146956 2746 147076 2774
rect 147048 921 147076 2746
rect 147772 2440 147824 2446
rect 147772 2382 147824 2388
rect 147128 1352 147180 1358
rect 147128 1294 147180 1300
rect 147034 912 147090 921
rect 147034 847 147090 856
rect 147140 785 147168 1294
rect 147784 950 147812 2382
rect 148152 1834 148180 2926
rect 148336 2774 148364 6734
rect 148416 6248 148468 6254
rect 148416 6190 148468 6196
rect 148428 5642 148456 6190
rect 148416 5636 148468 5642
rect 148416 5578 148468 5584
rect 148416 4208 148468 4214
rect 148416 4150 148468 4156
rect 148428 3466 148456 4150
rect 148704 3466 148732 8434
rect 149072 7886 149100 10270
rect 149702 10160 149758 10169
rect 149702 10095 149758 10104
rect 150990 10160 151046 10169
rect 150990 10095 151046 10104
rect 151634 10160 151690 10169
rect 151634 10095 151690 10104
rect 149716 9586 149744 10095
rect 150070 9888 150126 9897
rect 150070 9823 150126 9832
rect 149704 9580 149756 9586
rect 149704 9522 149756 9528
rect 150084 8974 150112 9823
rect 151004 9586 151032 10095
rect 151648 9586 151676 10095
rect 150992 9580 151044 9586
rect 150992 9522 151044 9528
rect 151636 9580 151688 9586
rect 151636 9522 151688 9528
rect 150532 9444 150584 9450
rect 150532 9386 150584 9392
rect 150440 9376 150492 9382
rect 150440 9318 150492 9324
rect 150072 8968 150124 8974
rect 150072 8910 150124 8916
rect 149888 8832 149940 8838
rect 149888 8774 149940 8780
rect 149060 7880 149112 7886
rect 149060 7822 149112 7828
rect 149152 7880 149204 7886
rect 149152 7822 149204 7828
rect 149164 6866 149192 7822
rect 148968 6860 149020 6866
rect 148968 6802 149020 6808
rect 149152 6860 149204 6866
rect 149152 6802 149204 6808
rect 148980 6390 149008 6802
rect 149428 6792 149480 6798
rect 149428 6734 149480 6740
rect 149440 6662 149468 6734
rect 149428 6656 149480 6662
rect 149428 6598 149480 6604
rect 148784 6384 148836 6390
rect 148784 6326 148836 6332
rect 148968 6384 149020 6390
rect 148968 6326 149020 6332
rect 148416 3460 148468 3466
rect 148416 3402 148468 3408
rect 148692 3460 148744 3466
rect 148692 3402 148744 3408
rect 148692 2984 148744 2990
rect 148796 2972 148824 6326
rect 148876 6316 148928 6322
rect 148876 6258 148928 6264
rect 148888 4214 148916 6258
rect 149900 5234 149928 8774
rect 150256 6996 150308 7002
rect 150256 6938 150308 6944
rect 150072 6656 150124 6662
rect 150072 6598 150124 6604
rect 150084 6322 150112 6598
rect 150072 6316 150124 6322
rect 150072 6258 150124 6264
rect 150268 6089 150296 6938
rect 150348 6860 150400 6866
rect 150348 6802 150400 6808
rect 150254 6080 150310 6089
rect 150254 6015 150310 6024
rect 149888 5228 149940 5234
rect 149888 5170 149940 5176
rect 148968 4480 149020 4486
rect 148968 4422 149020 4428
rect 148876 4208 148928 4214
rect 148876 4150 148928 4156
rect 148980 3602 149008 4422
rect 150360 4162 150388 6802
rect 150452 4690 150480 9318
rect 150544 6866 150572 9386
rect 151268 9376 151320 9382
rect 151268 9318 151320 9324
rect 150900 8016 150952 8022
rect 150900 7958 150952 7964
rect 150912 7206 150940 7958
rect 150992 7336 151044 7342
rect 150992 7278 151044 7284
rect 150900 7200 150952 7206
rect 150900 7142 150952 7148
rect 150532 6860 150584 6866
rect 150532 6802 150584 6808
rect 150900 6860 150952 6866
rect 150900 6802 150952 6808
rect 150624 6792 150676 6798
rect 150624 6734 150676 6740
rect 150532 5296 150584 5302
rect 150530 5264 150532 5273
rect 150584 5264 150586 5273
rect 150530 5199 150586 5208
rect 150440 4684 150492 4690
rect 150440 4626 150492 4632
rect 150360 4134 150480 4162
rect 149060 4072 149112 4078
rect 149796 4072 149848 4078
rect 149060 4014 149112 4020
rect 149794 4040 149796 4049
rect 149848 4040 149850 4049
rect 148968 3596 149020 3602
rect 148968 3538 149020 3544
rect 148876 3460 148928 3466
rect 148876 3402 148928 3408
rect 148888 3058 148916 3402
rect 148876 3052 148928 3058
rect 148876 2994 148928 3000
rect 148744 2944 148824 2972
rect 148692 2926 148744 2932
rect 148244 2746 148364 2774
rect 148796 2774 148824 2944
rect 148968 2984 149020 2990
rect 148968 2926 149020 2932
rect 148796 2746 148916 2774
rect 148140 1828 148192 1834
rect 148140 1770 148192 1776
rect 148244 1222 148272 2746
rect 148888 2582 148916 2746
rect 148876 2576 148928 2582
rect 148876 2518 148928 2524
rect 148980 2310 149008 2926
rect 149072 2774 149100 4014
rect 149794 3975 149850 3984
rect 150070 3496 150126 3505
rect 150070 3431 150072 3440
rect 150124 3431 150126 3440
rect 150072 3402 150124 3408
rect 149152 3392 149204 3398
rect 149152 3334 149204 3340
rect 149164 3074 149192 3334
rect 149164 3058 149468 3074
rect 149152 3052 149468 3058
rect 149204 3046 149468 3052
rect 149152 2994 149204 3000
rect 149244 2848 149296 2854
rect 149244 2790 149296 2796
rect 149072 2746 149192 2774
rect 149164 2650 149192 2746
rect 149152 2644 149204 2650
rect 149152 2586 149204 2592
rect 149150 2544 149206 2553
rect 149150 2479 149152 2488
rect 149204 2479 149206 2488
rect 149152 2450 149204 2456
rect 148968 2304 149020 2310
rect 148968 2246 149020 2252
rect 149256 1426 149284 2790
rect 149440 2446 149468 3046
rect 149428 2440 149480 2446
rect 149428 2382 149480 2388
rect 150072 1964 150124 1970
rect 150072 1906 150124 1912
rect 149244 1420 149296 1426
rect 149244 1362 149296 1368
rect 148416 1352 148468 1358
rect 148416 1294 148468 1300
rect 148508 1352 148560 1358
rect 148508 1294 148560 1300
rect 149704 1352 149756 1358
rect 149704 1294 149756 1300
rect 148232 1216 148284 1222
rect 148232 1158 148284 1164
rect 147772 944 147824 950
rect 147772 886 147824 892
rect 147126 776 147182 785
rect 146206 711 146262 720
rect 146760 740 146812 746
rect 147126 711 147182 720
rect 146760 682 146812 688
rect 143908 672 143960 678
rect 142066 640 142122 649
rect 148428 649 148456 1294
rect 148520 785 148548 1294
rect 148784 1284 148836 1290
rect 148784 1226 148836 1232
rect 148506 776 148562 785
rect 148506 711 148562 720
rect 143908 614 143960 620
rect 148414 640 148470 649
rect 142066 575 142122 584
rect 148414 575 148470 584
rect 140686 504 140742 513
rect 148796 474 148824 1226
rect 149716 785 149744 1294
rect 150084 1057 150112 1906
rect 150452 1873 150480 4134
rect 150438 1864 150494 1873
rect 150438 1799 150494 1808
rect 150636 1290 150664 6734
rect 150716 6384 150768 6390
rect 150912 6372 150940 6802
rect 150768 6344 150940 6372
rect 150716 6326 150768 6332
rect 150912 5166 150940 6344
rect 151004 6254 151032 7278
rect 151084 6656 151136 6662
rect 151084 6598 151136 6604
rect 150992 6248 151044 6254
rect 150992 6190 151044 6196
rect 150808 5160 150860 5166
rect 150808 5102 150860 5108
rect 150900 5160 150952 5166
rect 150900 5102 150952 5108
rect 150716 4616 150768 4622
rect 150716 4558 150768 4564
rect 150624 1284 150676 1290
rect 150624 1226 150676 1232
rect 150728 1222 150756 4558
rect 150820 2106 150848 5102
rect 150912 4690 150940 5102
rect 150900 4684 150952 4690
rect 150900 4626 150952 4632
rect 151004 4162 151032 6190
rect 151096 4758 151124 6598
rect 151084 4752 151136 4758
rect 151084 4694 151136 4700
rect 151096 4282 151124 4694
rect 151176 4684 151228 4690
rect 151176 4626 151228 4632
rect 151084 4276 151136 4282
rect 151084 4218 151136 4224
rect 150900 4140 150952 4146
rect 151004 4134 151124 4162
rect 150900 4082 150952 4088
rect 150808 2100 150860 2106
rect 150808 2042 150860 2048
rect 150912 1222 150940 4082
rect 150992 3936 151044 3942
rect 150992 3878 151044 3884
rect 151004 3194 151032 3878
rect 150992 3188 151044 3194
rect 150992 3130 151044 3136
rect 151096 2774 151124 4134
rect 151188 3466 151216 4626
rect 151280 4078 151308 9318
rect 151740 8294 151768 10338
rect 152278 10160 152334 10169
rect 152278 10095 152334 10104
rect 152292 9586 152320 10095
rect 152280 9580 152332 9586
rect 152280 9522 152332 9528
rect 152384 9518 152412 10814
rect 152464 10804 152516 10810
rect 152464 10746 152516 10752
rect 152476 9722 152504 10746
rect 162308 10464 162360 10470
rect 162308 10406 162360 10412
rect 154210 10296 154266 10305
rect 154210 10231 154266 10240
rect 157246 10296 157302 10305
rect 157246 10231 157302 10240
rect 153198 10160 153254 10169
rect 153198 10095 153254 10104
rect 152464 9716 152516 9722
rect 152464 9658 152516 9664
rect 153212 9586 153240 10095
rect 154224 9586 154252 10231
rect 156512 10192 156564 10198
rect 154578 10160 154634 10169
rect 156512 10134 156564 10140
rect 154578 10095 154634 10104
rect 154592 9586 154620 10095
rect 155130 9888 155186 9897
rect 155130 9823 155186 9832
rect 153200 9580 153252 9586
rect 153200 9522 153252 9528
rect 154212 9580 154264 9586
rect 154212 9522 154264 9528
rect 154580 9580 154632 9586
rect 154580 9522 154632 9528
rect 152372 9512 152424 9518
rect 152372 9454 152424 9460
rect 151912 9376 151964 9382
rect 151912 9318 151964 9324
rect 154580 9376 154632 9382
rect 154580 9318 154632 9324
rect 151728 8288 151780 8294
rect 151728 8230 151780 8236
rect 151358 7984 151414 7993
rect 151358 7919 151414 7928
rect 151372 6338 151400 7919
rect 151452 7744 151504 7750
rect 151452 7686 151504 7692
rect 151464 6866 151492 7686
rect 151452 6860 151504 6866
rect 151452 6802 151504 6808
rect 151544 6792 151596 6798
rect 151544 6734 151596 6740
rect 151728 6792 151780 6798
rect 151728 6734 151780 6740
rect 151372 6310 151492 6338
rect 151358 5264 151414 5273
rect 151358 5199 151414 5208
rect 151372 5166 151400 5199
rect 151360 5160 151412 5166
rect 151360 5102 151412 5108
rect 151464 4622 151492 6310
rect 151452 4616 151504 4622
rect 151452 4558 151504 4564
rect 151268 4072 151320 4078
rect 151268 4014 151320 4020
rect 151176 3460 151228 3466
rect 151176 3402 151228 3408
rect 151004 2746 151124 2774
rect 151004 2514 151032 2746
rect 150992 2508 151044 2514
rect 150992 2450 151044 2456
rect 150992 1352 151044 1358
rect 150992 1294 151044 1300
rect 150716 1216 150768 1222
rect 150716 1158 150768 1164
rect 150900 1216 150952 1222
rect 150900 1158 150952 1164
rect 150070 1048 150126 1057
rect 150070 983 150126 992
rect 151004 785 151032 1294
rect 149702 776 149758 785
rect 149702 711 149758 720
rect 150990 776 151046 785
rect 150990 711 151046 720
rect 140686 439 140742 448
rect 148784 468 148836 474
rect 148784 410 148836 416
rect 151556 406 151584 6734
rect 151740 6662 151768 6734
rect 151728 6656 151780 6662
rect 151728 6598 151780 6604
rect 151728 5160 151780 5166
rect 151728 5102 151780 5108
rect 151820 5160 151872 5166
rect 151820 5102 151872 5108
rect 151636 4616 151688 4622
rect 151636 4558 151688 4564
rect 151648 4457 151676 4558
rect 151634 4448 151690 4457
rect 151634 4383 151690 4392
rect 151636 1352 151688 1358
rect 151636 1294 151688 1300
rect 151648 785 151676 1294
rect 151740 1057 151768 5102
rect 151832 4486 151860 5102
rect 151924 4690 151952 9318
rect 152832 8016 152884 8022
rect 152832 7958 152884 7964
rect 152556 7948 152608 7954
rect 152556 7890 152608 7896
rect 152568 7478 152596 7890
rect 152372 7472 152424 7478
rect 152372 7414 152424 7420
rect 152556 7472 152608 7478
rect 152556 7414 152608 7420
rect 152384 6866 152412 7414
rect 152372 6860 152424 6866
rect 152372 6802 152424 6808
rect 152372 6656 152424 6662
rect 152372 6598 152424 6604
rect 152646 6624 152702 6633
rect 152004 5568 152056 5574
rect 152004 5510 152056 5516
rect 151912 4684 151964 4690
rect 151912 4626 151964 4632
rect 152016 4593 152044 5510
rect 152384 5370 152412 6598
rect 152646 6559 152702 6568
rect 152660 6390 152688 6559
rect 152648 6384 152700 6390
rect 152646 6352 152648 6361
rect 152740 6384 152792 6390
rect 152700 6352 152702 6361
rect 152740 6326 152792 6332
rect 152646 6287 152702 6296
rect 152752 5778 152780 6326
rect 152740 5772 152792 5778
rect 152740 5714 152792 5720
rect 152844 5658 152872 7958
rect 154118 7848 154174 7857
rect 154118 7783 154174 7792
rect 153292 6248 153344 6254
rect 153292 6190 153344 6196
rect 152660 5630 152872 5658
rect 153304 5642 153332 6190
rect 153384 5704 153436 5710
rect 153384 5646 153436 5652
rect 153292 5636 153344 5642
rect 152372 5364 152424 5370
rect 152372 5306 152424 5312
rect 152372 5160 152424 5166
rect 152372 5102 152424 5108
rect 152384 4622 152412 5102
rect 152464 4752 152516 4758
rect 152464 4694 152516 4700
rect 152372 4616 152424 4622
rect 152002 4584 152058 4593
rect 152372 4558 152424 4564
rect 152002 4519 152058 4528
rect 152280 4548 152332 4554
rect 152280 4490 152332 4496
rect 151820 4480 151872 4486
rect 152292 4434 152320 4490
rect 151820 4422 151872 4428
rect 151924 4406 152320 4434
rect 151924 4298 151952 4406
rect 151832 4270 151952 4298
rect 151832 4214 151860 4270
rect 151820 4208 151872 4214
rect 151820 4150 151872 4156
rect 152476 4078 152504 4694
rect 152660 4146 152688 5630
rect 153292 5578 153344 5584
rect 153304 5302 153332 5578
rect 153396 5370 153424 5646
rect 153384 5364 153436 5370
rect 153384 5306 153436 5312
rect 153292 5296 153344 5302
rect 153292 5238 153344 5244
rect 153752 5024 153804 5030
rect 153752 4966 153804 4972
rect 153764 4826 153792 4966
rect 153752 4820 153804 4826
rect 153752 4762 153804 4768
rect 154132 4622 154160 7783
rect 153384 4616 153436 4622
rect 153384 4558 153436 4564
rect 154120 4616 154172 4622
rect 154120 4558 154172 4564
rect 154304 4616 154356 4622
rect 154304 4558 154356 4564
rect 154396 4616 154448 4622
rect 154396 4558 154448 4564
rect 152648 4140 152700 4146
rect 152648 4082 152700 4088
rect 152464 4072 152516 4078
rect 152464 4014 152516 4020
rect 152832 4072 152884 4078
rect 152832 4014 152884 4020
rect 152924 4072 152976 4078
rect 152924 4014 152976 4020
rect 152844 3738 152872 4014
rect 152372 3732 152424 3738
rect 152372 3674 152424 3680
rect 152832 3732 152884 3738
rect 152832 3674 152884 3680
rect 152384 3534 152412 3674
rect 152372 3528 152424 3534
rect 152372 3470 152424 3476
rect 152384 2514 152412 3470
rect 152936 3126 152964 4014
rect 152924 3120 152976 3126
rect 152924 3062 152976 3068
rect 153108 2848 153160 2854
rect 153108 2790 153160 2796
rect 152372 2508 152424 2514
rect 152372 2450 152424 2456
rect 153120 1737 153148 2790
rect 153396 2774 153424 4558
rect 153304 2746 153424 2774
rect 153106 1728 153162 1737
rect 153106 1663 153162 1672
rect 152280 1352 152332 1358
rect 152280 1294 152332 1300
rect 153200 1352 153252 1358
rect 153200 1294 153252 1300
rect 152096 1216 152148 1222
rect 152096 1158 152148 1164
rect 151726 1048 151782 1057
rect 151726 983 151782 992
rect 152108 950 152136 1158
rect 152096 944 152148 950
rect 152096 886 152148 892
rect 152292 785 152320 1294
rect 152464 876 152516 882
rect 152464 818 152516 824
rect 152556 876 152608 882
rect 152556 818 152608 824
rect 151634 776 151690 785
rect 151634 711 151690 720
rect 152278 776 152334 785
rect 152278 711 152334 720
rect 152476 542 152504 818
rect 152464 536 152516 542
rect 152464 478 152516 484
rect 152568 406 152596 818
rect 153212 785 153240 1294
rect 153304 1290 153332 2746
rect 154212 1352 154264 1358
rect 154212 1294 154264 1300
rect 153292 1284 153344 1290
rect 153292 1226 153344 1232
rect 153198 776 153254 785
rect 153198 711 153254 720
rect 154224 649 154252 1294
rect 154210 640 154266 649
rect 154210 575 154266 584
rect 154316 406 154344 4558
rect 154408 4282 154436 4558
rect 154396 4276 154448 4282
rect 154396 4218 154448 4224
rect 154408 3398 154436 4218
rect 154488 4140 154540 4146
rect 154488 4082 154540 4088
rect 154500 3670 154528 4082
rect 154488 3664 154540 3670
rect 154488 3606 154540 3612
rect 154592 3602 154620 9318
rect 155144 8974 155172 9823
rect 155958 9752 156014 9761
rect 155868 9716 155920 9722
rect 155958 9687 155960 9696
rect 155868 9658 155920 9664
rect 156012 9687 156014 9696
rect 155960 9658 156012 9664
rect 155880 9602 155908 9658
rect 155776 9580 155828 9586
rect 155604 9540 155776 9568
rect 155604 9382 155632 9540
rect 155880 9574 156000 9602
rect 155776 9522 155828 9528
rect 155776 9444 155828 9450
rect 155776 9386 155828 9392
rect 155592 9376 155644 9382
rect 155592 9318 155644 9324
rect 155500 9172 155552 9178
rect 155500 9114 155552 9120
rect 155132 8968 155184 8974
rect 155132 8910 155184 8916
rect 155512 8838 155540 9114
rect 155684 8968 155736 8974
rect 155788 8956 155816 9386
rect 155736 8928 155816 8956
rect 155684 8910 155736 8916
rect 155500 8832 155552 8838
rect 155500 8774 155552 8780
rect 155776 8832 155828 8838
rect 155776 8774 155828 8780
rect 155592 7540 155644 7546
rect 155592 7482 155644 7488
rect 155604 6730 155632 7482
rect 155592 6724 155644 6730
rect 155592 6666 155644 6672
rect 155040 6112 155092 6118
rect 155040 6054 155092 6060
rect 155052 5778 155080 6054
rect 155040 5772 155092 5778
rect 155040 5714 155092 5720
rect 155684 5704 155736 5710
rect 155684 5646 155736 5652
rect 155224 4480 155276 4486
rect 155224 4422 155276 4428
rect 154672 4208 154724 4214
rect 154672 4150 154724 4156
rect 154580 3596 154632 3602
rect 154580 3538 154632 3544
rect 154684 3534 154712 4150
rect 154856 4072 154908 4078
rect 154856 4014 154908 4020
rect 154672 3528 154724 3534
rect 154672 3470 154724 3476
rect 154868 3466 154896 4014
rect 155236 3534 155264 4422
rect 155696 4146 155724 5646
rect 155684 4140 155736 4146
rect 155684 4082 155736 4088
rect 155684 3732 155736 3738
rect 155684 3674 155736 3680
rect 155224 3528 155276 3534
rect 155224 3470 155276 3476
rect 154856 3460 154908 3466
rect 154856 3402 154908 3408
rect 154396 3392 154448 3398
rect 154396 3334 154448 3340
rect 155038 3360 155094 3369
rect 155038 3295 155094 3304
rect 155052 1902 155080 3295
rect 155130 2680 155186 2689
rect 155130 2615 155186 2624
rect 155144 2582 155172 2615
rect 155132 2576 155184 2582
rect 155132 2518 155184 2524
rect 155224 2440 155276 2446
rect 155224 2382 155276 2388
rect 155040 1896 155092 1902
rect 155040 1838 155092 1844
rect 154580 1352 154632 1358
rect 155236 1329 155264 2382
rect 155696 2281 155724 3674
rect 155788 2378 155816 8774
rect 155868 5636 155920 5642
rect 155868 5578 155920 5584
rect 155880 5166 155908 5578
rect 155868 5160 155920 5166
rect 155868 5102 155920 5108
rect 155880 4554 155908 5102
rect 155868 4548 155920 4554
rect 155868 4490 155920 4496
rect 155868 3528 155920 3534
rect 155868 3470 155920 3476
rect 155776 2372 155828 2378
rect 155776 2314 155828 2320
rect 155682 2272 155738 2281
rect 155682 2207 155738 2216
rect 155776 1828 155828 1834
rect 155776 1770 155828 1776
rect 155788 1601 155816 1770
rect 155774 1592 155830 1601
rect 155774 1527 155830 1536
rect 154580 1294 154632 1300
rect 155222 1320 155278 1329
rect 154592 785 154620 1294
rect 155222 1255 155278 1264
rect 155880 950 155908 3470
rect 155972 3058 156000 9574
rect 156144 9580 156196 9586
rect 156144 9522 156196 9528
rect 156156 9178 156184 9522
rect 156144 9172 156196 9178
rect 156144 9114 156196 9120
rect 156524 8430 156552 10134
rect 156878 9752 156934 9761
rect 157260 9722 157288 10231
rect 162216 10192 162268 10198
rect 162216 10134 162268 10140
rect 158628 10124 158680 10130
rect 158628 10066 158680 10072
rect 157982 9752 158038 9761
rect 156878 9687 156880 9696
rect 156932 9687 156934 9696
rect 157248 9716 157300 9722
rect 156880 9658 156932 9664
rect 157982 9687 157984 9696
rect 157248 9658 157300 9664
rect 158036 9687 158038 9696
rect 157984 9658 158036 9664
rect 156972 9580 157024 9586
rect 156972 9522 157024 9528
rect 157432 9580 157484 9586
rect 157432 9522 157484 9528
rect 157800 9580 157852 9586
rect 157800 9522 157852 9528
rect 156984 9178 157012 9522
rect 156972 9172 157024 9178
rect 156972 9114 157024 9120
rect 156696 8968 156748 8974
rect 156696 8910 156748 8916
rect 156708 8838 156736 8910
rect 156696 8832 156748 8838
rect 156696 8774 156748 8780
rect 157156 8832 157208 8838
rect 157156 8774 157208 8780
rect 157248 8832 157300 8838
rect 157248 8774 157300 8780
rect 156512 8424 156564 8430
rect 156512 8366 156564 8372
rect 156052 7200 156104 7206
rect 156052 7142 156104 7148
rect 156064 6769 156092 7142
rect 156050 6760 156106 6769
rect 156050 6695 156106 6704
rect 156144 6316 156196 6322
rect 156144 6258 156196 6264
rect 156052 5024 156104 5030
rect 156052 4966 156104 4972
rect 156064 4758 156092 4966
rect 156052 4752 156104 4758
rect 156052 4694 156104 4700
rect 156052 3664 156104 3670
rect 156052 3606 156104 3612
rect 156064 3233 156092 3606
rect 156050 3224 156106 3233
rect 156050 3159 156106 3168
rect 156156 3126 156184 6258
rect 156328 6112 156380 6118
rect 156328 6054 156380 6060
rect 156340 4486 156368 6054
rect 156420 4548 156472 4554
rect 156420 4490 156472 4496
rect 156328 4480 156380 4486
rect 156328 4422 156380 4428
rect 156328 4140 156380 4146
rect 156328 4082 156380 4088
rect 156236 4072 156288 4078
rect 156236 4014 156288 4020
rect 156144 3120 156196 3126
rect 156144 3062 156196 3068
rect 155960 3052 156012 3058
rect 155960 2994 156012 3000
rect 156144 2984 156196 2990
rect 156144 2926 156196 2932
rect 156052 2848 156104 2854
rect 156052 2790 156104 2796
rect 155960 1760 156012 1766
rect 155960 1702 156012 1708
rect 155972 1465 156000 1702
rect 155958 1456 156014 1465
rect 155958 1391 156014 1400
rect 156064 1222 156092 2790
rect 156156 1358 156184 2926
rect 156144 1352 156196 1358
rect 156144 1294 156196 1300
rect 156248 1290 156276 4014
rect 156340 3602 156368 4082
rect 156328 3596 156380 3602
rect 156328 3538 156380 3544
rect 156432 2553 156460 4490
rect 156418 2544 156474 2553
rect 156418 2479 156474 2488
rect 156524 2310 156552 8366
rect 156788 6316 156840 6322
rect 156788 6258 156840 6264
rect 156972 6316 157024 6322
rect 156972 6258 157024 6264
rect 156800 5030 156828 6258
rect 156984 5846 157012 6258
rect 157064 6248 157116 6254
rect 157064 6190 157116 6196
rect 156972 5840 157024 5846
rect 156972 5782 157024 5788
rect 156788 5024 156840 5030
rect 156788 4966 156840 4972
rect 156604 4820 156656 4826
rect 156604 4762 156656 4768
rect 156616 3602 156644 4762
rect 156972 3936 157024 3942
rect 156972 3878 157024 3884
rect 156694 3632 156750 3641
rect 156604 3596 156656 3602
rect 156694 3567 156696 3576
rect 156604 3538 156656 3544
rect 156748 3567 156750 3576
rect 156880 3596 156932 3602
rect 156696 3538 156748 3544
rect 156880 3538 156932 3544
rect 156892 3398 156920 3538
rect 156984 3398 157012 3878
rect 156880 3392 156932 3398
rect 156880 3334 156932 3340
rect 156972 3392 157024 3398
rect 156972 3334 157024 3340
rect 156602 3224 156658 3233
rect 156602 3159 156658 3168
rect 156616 2922 156644 3159
rect 156984 3058 157012 3334
rect 157076 3233 157104 6190
rect 157062 3224 157118 3233
rect 157062 3159 157118 3168
rect 156880 3052 156932 3058
rect 156800 3012 156880 3040
rect 156604 2916 156656 2922
rect 156604 2858 156656 2864
rect 156800 2553 156828 3012
rect 156880 2994 156932 3000
rect 156972 3052 157024 3058
rect 156972 2994 157024 3000
rect 157168 2650 157196 8774
rect 157260 8430 157288 8774
rect 157444 8634 157472 9522
rect 157708 9376 157760 9382
rect 157708 9318 157760 9324
rect 157524 8968 157576 8974
rect 157524 8910 157576 8916
rect 157616 8968 157668 8974
rect 157616 8910 157668 8916
rect 157432 8628 157484 8634
rect 157432 8570 157484 8576
rect 157248 8424 157300 8430
rect 157248 8366 157300 8372
rect 157248 6248 157300 6254
rect 157248 6190 157300 6196
rect 157260 4826 157288 6190
rect 157248 4820 157300 4826
rect 157248 4762 157300 4768
rect 157246 2816 157302 2825
rect 157302 2774 157380 2802
rect 157246 2751 157302 2760
rect 157352 2650 157380 2774
rect 156880 2644 156932 2650
rect 156880 2586 156932 2592
rect 156972 2644 157024 2650
rect 156972 2586 157024 2592
rect 157156 2644 157208 2650
rect 157156 2586 157208 2592
rect 157340 2644 157392 2650
rect 157340 2586 157392 2592
rect 156786 2544 156842 2553
rect 156892 2514 156920 2586
rect 156786 2479 156842 2488
rect 156880 2508 156932 2514
rect 156880 2450 156932 2456
rect 156604 2440 156656 2446
rect 156604 2382 156656 2388
rect 156328 2304 156380 2310
rect 156328 2246 156380 2252
rect 156512 2304 156564 2310
rect 156512 2246 156564 2252
rect 156340 1884 156368 2246
rect 156512 1896 156564 1902
rect 156340 1856 156512 1884
rect 156512 1838 156564 1844
rect 156512 1556 156564 1562
rect 156512 1498 156564 1504
rect 156524 1426 156552 1498
rect 156512 1420 156564 1426
rect 156512 1362 156564 1368
rect 156616 1329 156644 2382
rect 156880 2372 156932 2378
rect 156880 2314 156932 2320
rect 156892 2122 156920 2314
rect 156984 2258 157012 2586
rect 157536 2530 157564 8910
rect 157628 8498 157656 8910
rect 157616 8492 157668 8498
rect 157616 8434 157668 8440
rect 157720 4078 157748 9318
rect 157812 9178 157840 9522
rect 157984 9512 158036 9518
rect 157984 9454 158036 9460
rect 157800 9172 157852 9178
rect 157800 9114 157852 9120
rect 157800 5364 157852 5370
rect 157800 5306 157852 5312
rect 157812 4214 157840 5306
rect 157892 4616 157944 4622
rect 157892 4558 157944 4564
rect 157800 4208 157852 4214
rect 157800 4150 157852 4156
rect 157708 4072 157760 4078
rect 157708 4014 157760 4020
rect 157904 3126 157932 4558
rect 157892 3120 157944 3126
rect 157892 3062 157944 3068
rect 157996 2990 158024 9454
rect 158352 9104 158404 9110
rect 158352 9046 158404 9052
rect 158168 6316 158220 6322
rect 158168 6258 158220 6264
rect 158076 5568 158128 5574
rect 158076 5510 158128 5516
rect 158088 5098 158116 5510
rect 158076 5092 158128 5098
rect 158076 5034 158128 5040
rect 158088 4554 158116 5034
rect 158076 4548 158128 4554
rect 158076 4490 158128 4496
rect 158180 4486 158208 6258
rect 158260 5160 158312 5166
rect 158260 5102 158312 5108
rect 158168 4480 158220 4486
rect 158168 4422 158220 4428
rect 158272 3738 158300 5102
rect 158260 3732 158312 3738
rect 158260 3674 158312 3680
rect 158364 3602 158392 9046
rect 158640 7886 158668 10066
rect 160928 10056 160980 10062
rect 160928 9998 160980 10004
rect 158720 9988 158772 9994
rect 158720 9930 158772 9936
rect 158732 8906 158760 9930
rect 159454 9752 159510 9761
rect 159454 9687 159456 9696
rect 159508 9687 159510 9696
rect 159456 9658 159508 9664
rect 159272 9580 159324 9586
rect 159272 9522 159324 9528
rect 159364 9580 159416 9586
rect 159364 9522 159416 9528
rect 158720 8900 158772 8906
rect 158720 8842 158772 8848
rect 158732 8430 158760 8842
rect 159284 8634 159312 9522
rect 159376 8634 159404 9522
rect 160940 9518 160968 9998
rect 161388 9920 161440 9926
rect 161388 9862 161440 9868
rect 160928 9512 160980 9518
rect 159454 9480 159510 9489
rect 160928 9454 160980 9460
rect 159454 9415 159456 9424
rect 159508 9415 159510 9424
rect 159456 9386 159508 9392
rect 159824 9172 159876 9178
rect 159824 9114 159876 9120
rect 159836 8974 159864 9114
rect 160008 9104 160060 9110
rect 160008 9046 160060 9052
rect 159824 8968 159876 8974
rect 159824 8910 159876 8916
rect 159916 8968 159968 8974
rect 159916 8910 159968 8916
rect 159640 8900 159692 8906
rect 159640 8842 159692 8848
rect 159272 8628 159324 8634
rect 159272 8570 159324 8576
rect 159364 8628 159416 8634
rect 159364 8570 159416 8576
rect 158720 8424 158772 8430
rect 158720 8366 158772 8372
rect 159088 8424 159140 8430
rect 159088 8366 159140 8372
rect 158628 7880 158680 7886
rect 158628 7822 158680 7828
rect 158628 7336 158680 7342
rect 158628 7278 158680 7284
rect 158640 5273 158668 7278
rect 158812 6112 158864 6118
rect 158812 6054 158864 6060
rect 158626 5264 158682 5273
rect 158626 5199 158682 5208
rect 158536 5160 158588 5166
rect 158536 5102 158588 5108
rect 158548 4826 158576 5102
rect 158628 5024 158680 5030
rect 158628 4966 158680 4972
rect 158536 4820 158588 4826
rect 158536 4762 158588 4768
rect 158548 4554 158576 4762
rect 158536 4548 158588 4554
rect 158536 4490 158588 4496
rect 158640 4078 158668 4966
rect 158628 4072 158680 4078
rect 158628 4014 158680 4020
rect 158640 3738 158668 4014
rect 158628 3732 158680 3738
rect 158628 3674 158680 3680
rect 158352 3596 158404 3602
rect 158352 3538 158404 3544
rect 158536 3528 158588 3534
rect 158536 3470 158588 3476
rect 157984 2984 158036 2990
rect 157984 2926 158036 2932
rect 158352 2848 158404 2854
rect 158352 2790 158404 2796
rect 157168 2502 157840 2530
rect 156984 2230 157104 2258
rect 156892 2094 157012 2122
rect 156696 1964 156748 1970
rect 156696 1906 156748 1912
rect 156788 1964 156840 1970
rect 156788 1906 156840 1912
rect 156708 1562 156736 1906
rect 156696 1556 156748 1562
rect 156696 1498 156748 1504
rect 156602 1320 156658 1329
rect 156236 1284 156288 1290
rect 156602 1255 156658 1264
rect 156236 1226 156288 1232
rect 156052 1216 156104 1222
rect 156052 1158 156104 1164
rect 155868 944 155920 950
rect 155868 886 155920 892
rect 156800 785 156828 1906
rect 156880 1828 156932 1834
rect 156880 1770 156932 1776
rect 156892 1601 156920 1770
rect 156878 1592 156934 1601
rect 156878 1527 156934 1536
rect 156984 1222 157012 2094
rect 157076 1902 157104 2230
rect 157168 2038 157196 2502
rect 157812 2446 157840 2502
rect 157340 2440 157392 2446
rect 157340 2382 157392 2388
rect 157708 2440 157760 2446
rect 157708 2382 157760 2388
rect 157800 2440 157852 2446
rect 157800 2382 157852 2388
rect 157156 2032 157208 2038
rect 157156 1974 157208 1980
rect 157064 1896 157116 1902
rect 157064 1838 157116 1844
rect 157076 1426 157104 1838
rect 157352 1562 157380 2382
rect 157432 2304 157484 2310
rect 157432 2246 157484 2252
rect 157340 1556 157392 1562
rect 157340 1498 157392 1504
rect 157444 1465 157472 2246
rect 157430 1456 157486 1465
rect 157064 1420 157116 1426
rect 157430 1391 157486 1400
rect 157064 1362 157116 1368
rect 157720 1222 157748 2382
rect 158168 2372 158220 2378
rect 158168 2314 158220 2320
rect 157892 2100 157944 2106
rect 157892 2042 157944 2048
rect 157984 2100 158036 2106
rect 157984 2042 158036 2048
rect 157904 1465 157932 2042
rect 157996 1970 158024 2042
rect 157984 1964 158036 1970
rect 157984 1906 158036 1912
rect 158180 1902 158208 2314
rect 158168 1896 158220 1902
rect 158168 1838 158220 1844
rect 157890 1456 157946 1465
rect 158180 1426 158208 1838
rect 157890 1391 157946 1400
rect 158168 1420 158220 1426
rect 158168 1362 158220 1368
rect 156972 1216 157024 1222
rect 156972 1158 157024 1164
rect 157708 1216 157760 1222
rect 157708 1158 157760 1164
rect 154578 776 154634 785
rect 154578 711 154634 720
rect 156786 776 156842 785
rect 156786 711 156842 720
rect 158364 542 158392 2790
rect 158548 2689 158576 3470
rect 158640 2922 158668 3674
rect 158824 3058 158852 6054
rect 158812 3052 158864 3058
rect 158812 2994 158864 3000
rect 158904 3052 158956 3058
rect 158904 2994 158956 3000
rect 158628 2916 158680 2922
rect 158628 2858 158680 2864
rect 158534 2680 158590 2689
rect 158534 2615 158590 2624
rect 158628 2440 158680 2446
rect 158628 2382 158680 2388
rect 158536 2372 158588 2378
rect 158536 2314 158588 2320
rect 158548 1902 158576 2314
rect 158536 1896 158588 1902
rect 158536 1838 158588 1844
rect 158352 536 158404 542
rect 158640 513 158668 2382
rect 158812 1284 158864 1290
rect 158812 1226 158864 1232
rect 158824 649 158852 1226
rect 158916 882 158944 2994
rect 159100 1426 159128 8366
rect 159272 7200 159324 7206
rect 159272 7142 159324 7148
rect 159180 6928 159232 6934
rect 159180 6870 159232 6876
rect 159192 4146 159220 6870
rect 159180 4140 159232 4146
rect 159180 4082 159232 4088
rect 159284 3602 159312 7142
rect 159456 5296 159508 5302
rect 159456 5238 159508 5244
rect 159468 4146 159496 5238
rect 159456 4140 159508 4146
rect 159456 4082 159508 4088
rect 159468 4026 159496 4082
rect 159468 3998 159588 4026
rect 159560 3602 159588 3998
rect 159272 3596 159324 3602
rect 159272 3538 159324 3544
rect 159548 3596 159600 3602
rect 159548 3538 159600 3544
rect 159456 3528 159508 3534
rect 159456 3470 159508 3476
rect 159468 2582 159496 3470
rect 159560 2922 159588 3538
rect 159548 2916 159600 2922
rect 159548 2858 159600 2864
rect 159456 2576 159508 2582
rect 159456 2518 159508 2524
rect 159652 1970 159680 8842
rect 159824 8628 159876 8634
rect 159824 8570 159876 8576
rect 159836 8430 159864 8570
rect 159824 8424 159876 8430
rect 159824 8366 159876 8372
rect 159836 2774 159864 8366
rect 159928 8362 159956 8910
rect 159916 8356 159968 8362
rect 159916 8298 159968 8304
rect 160020 7750 160048 9046
rect 160836 8968 160888 8974
rect 160836 8910 160888 8916
rect 160848 8566 160876 8910
rect 160836 8560 160888 8566
rect 160836 8502 160888 8508
rect 160282 8392 160338 8401
rect 160940 8362 160968 9454
rect 161112 9376 161164 9382
rect 161112 9318 161164 9324
rect 160282 8327 160338 8336
rect 160928 8356 160980 8362
rect 160100 8288 160152 8294
rect 160100 8230 160152 8236
rect 160112 7886 160140 8230
rect 160296 8090 160324 8327
rect 160928 8298 160980 8304
rect 160284 8084 160336 8090
rect 160284 8026 160336 8032
rect 160100 7880 160152 7886
rect 160100 7822 160152 7828
rect 160008 7744 160060 7750
rect 160008 7686 160060 7692
rect 160652 5704 160704 5710
rect 160652 5646 160704 5652
rect 160664 5574 160692 5646
rect 160560 5568 160612 5574
rect 160560 5510 160612 5516
rect 160652 5568 160704 5574
rect 160652 5510 160704 5516
rect 160572 5273 160600 5510
rect 160558 5264 160614 5273
rect 160558 5199 160614 5208
rect 160008 5160 160060 5166
rect 160008 5102 160060 5108
rect 160020 5030 160048 5102
rect 160008 5024 160060 5030
rect 159928 4972 160008 4978
rect 159928 4966 160060 4972
rect 159928 4950 160048 4966
rect 159928 3913 159956 4950
rect 160008 4820 160060 4826
rect 160008 4762 160060 4768
rect 159914 3904 159970 3913
rect 159914 3839 159970 3848
rect 160020 3097 160048 4762
rect 160834 4584 160890 4593
rect 160834 4519 160836 4528
rect 160888 4519 160890 4528
rect 160836 4490 160888 4496
rect 160744 4140 160796 4146
rect 160744 4082 160796 4088
rect 160468 3936 160520 3942
rect 160468 3878 160520 3884
rect 160006 3088 160062 3097
rect 160006 3023 160062 3032
rect 160192 3052 160244 3058
rect 160192 2994 160244 3000
rect 160006 2816 160062 2825
rect 159836 2746 159956 2774
rect 160062 2760 160140 2774
rect 160006 2751 160140 2760
rect 160020 2746 160140 2751
rect 159928 2446 159956 2746
rect 160112 2650 160140 2746
rect 160100 2644 160152 2650
rect 160100 2586 160152 2592
rect 160204 2530 160232 2994
rect 160112 2502 160232 2530
rect 159916 2440 159968 2446
rect 159916 2382 159968 2388
rect 160008 2440 160060 2446
rect 160008 2382 160060 2388
rect 159272 1964 159324 1970
rect 159272 1906 159324 1912
rect 159640 1964 159692 1970
rect 159640 1906 159692 1912
rect 159088 1420 159140 1426
rect 159088 1362 159140 1368
rect 159284 1358 159312 1906
rect 160020 1902 160048 2382
rect 160008 1896 160060 1902
rect 160008 1838 160060 1844
rect 159272 1352 159324 1358
rect 159272 1294 159324 1300
rect 158904 876 158956 882
rect 158904 818 158956 824
rect 158810 640 158866 649
rect 158810 575 158866 584
rect 158352 478 158404 484
rect 158626 504 158682 513
rect 158626 439 158682 448
rect 151544 400 151596 406
rect 90822 368 90878 377
rect 90822 303 90878 312
rect 91742 368 91798 377
rect 91742 303 91798 312
rect 93030 368 93086 377
rect 93030 303 93086 312
rect 98734 368 98790 377
rect 98734 303 98790 312
rect 113546 368 113602 377
rect 113546 303 113602 312
rect 130842 368 130898 377
rect 151544 342 151596 348
rect 152556 400 152608 406
rect 152556 342 152608 348
rect 154304 400 154356 406
rect 160112 377 160140 2502
rect 160376 2440 160428 2446
rect 160376 2382 160428 2388
rect 160192 1760 160244 1766
rect 160192 1702 160244 1708
rect 160204 1358 160232 1702
rect 160388 1426 160416 2382
rect 160376 1420 160428 1426
rect 160376 1362 160428 1368
rect 160192 1352 160244 1358
rect 160192 1294 160244 1300
rect 160480 474 160508 3878
rect 160560 3392 160612 3398
rect 160560 3334 160612 3340
rect 160652 3392 160704 3398
rect 160652 3334 160704 3340
rect 160572 3058 160600 3334
rect 160560 3052 160612 3058
rect 160560 2994 160612 3000
rect 160664 2854 160692 3334
rect 160652 2848 160704 2854
rect 160652 2790 160704 2796
rect 160756 2650 160784 4082
rect 160836 3528 160888 3534
rect 160836 3470 160888 3476
rect 160848 3126 160876 3470
rect 160836 3120 160888 3126
rect 160836 3062 160888 3068
rect 160940 2774 160968 8298
rect 161124 7410 161152 9318
rect 161204 8968 161256 8974
rect 161204 8910 161256 8916
rect 161216 8634 161244 8910
rect 161204 8628 161256 8634
rect 161204 8570 161256 8576
rect 161294 8392 161350 8401
rect 161294 8327 161350 8336
rect 161308 7546 161336 8327
rect 161400 7954 161428 9862
rect 161664 9580 161716 9586
rect 161664 9522 161716 9528
rect 161572 8424 161624 8430
rect 161676 8412 161704 9522
rect 161756 9444 161808 9450
rect 161756 9386 161808 9392
rect 161768 8430 161796 9386
rect 161848 9376 161900 9382
rect 161848 9318 161900 9324
rect 161624 8384 161704 8412
rect 161572 8366 161624 8372
rect 161676 7954 161704 8384
rect 161756 8424 161808 8430
rect 161756 8366 161808 8372
rect 161388 7948 161440 7954
rect 161388 7890 161440 7896
rect 161664 7948 161716 7954
rect 161664 7890 161716 7896
rect 161296 7540 161348 7546
rect 161296 7482 161348 7488
rect 161112 7404 161164 7410
rect 161112 7346 161164 7352
rect 161400 6984 161428 7890
rect 161400 6956 161520 6984
rect 161112 6656 161164 6662
rect 161112 6598 161164 6604
rect 161124 5234 161152 6598
rect 161296 5772 161348 5778
rect 161296 5714 161348 5720
rect 161308 5574 161336 5714
rect 161296 5568 161348 5574
rect 161296 5510 161348 5516
rect 161112 5228 161164 5234
rect 161112 5170 161164 5176
rect 161388 5228 161440 5234
rect 161388 5170 161440 5176
rect 161204 5092 161256 5098
rect 161204 5034 161256 5040
rect 161020 4616 161072 4622
rect 161020 4558 161072 4564
rect 161032 3738 161060 4558
rect 161216 4554 161244 5034
rect 161400 4554 161428 5170
rect 161204 4548 161256 4554
rect 161204 4490 161256 4496
rect 161388 4548 161440 4554
rect 161388 4490 161440 4496
rect 161216 4298 161244 4490
rect 161216 4270 161336 4298
rect 161308 4214 161336 4270
rect 161296 4208 161348 4214
rect 161296 4150 161348 4156
rect 161020 3732 161072 3738
rect 161020 3674 161072 3680
rect 161308 3466 161336 4150
rect 161388 4072 161440 4078
rect 161388 4014 161440 4020
rect 161400 3942 161428 4014
rect 161388 3936 161440 3942
rect 161388 3878 161440 3884
rect 161296 3460 161348 3466
rect 161296 3402 161348 3408
rect 161308 2990 161336 3402
rect 161296 2984 161348 2990
rect 161296 2926 161348 2932
rect 161492 2774 161520 6956
rect 161860 6934 161888 9318
rect 162228 8974 162256 10134
rect 162320 9722 162348 10406
rect 163688 10056 163740 10062
rect 163688 9998 163740 10004
rect 162584 9988 162636 9994
rect 162584 9930 162636 9936
rect 162308 9716 162360 9722
rect 162308 9658 162360 9664
rect 162320 9586 162348 9658
rect 162400 9648 162452 9654
rect 162400 9590 162452 9596
rect 162308 9580 162360 9586
rect 162308 9522 162360 9528
rect 162216 8968 162268 8974
rect 162216 8910 162268 8916
rect 162412 8838 162440 9590
rect 162596 8974 162624 9930
rect 163596 9920 163648 9926
rect 163596 9862 163648 9868
rect 162768 9512 162820 9518
rect 162768 9454 162820 9460
rect 162584 8968 162636 8974
rect 162584 8910 162636 8916
rect 162400 8832 162452 8838
rect 162400 8774 162452 8780
rect 162306 8528 162362 8537
rect 161940 8492 161992 8498
rect 162306 8463 162362 8472
rect 162676 8492 162728 8498
rect 161940 8434 161992 8440
rect 161952 8362 161980 8434
rect 162216 8424 162268 8430
rect 162216 8366 162268 8372
rect 161940 8356 161992 8362
rect 161940 8298 161992 8304
rect 161848 6928 161900 6934
rect 161848 6870 161900 6876
rect 161572 6248 161624 6254
rect 161572 6190 161624 6196
rect 161584 5234 161612 6190
rect 162032 5636 162084 5642
rect 162032 5578 162084 5584
rect 161572 5228 161624 5234
rect 161572 5170 161624 5176
rect 161584 5030 161612 5170
rect 161572 5024 161624 5030
rect 161572 4966 161624 4972
rect 162044 4486 162072 5578
rect 162122 5128 162178 5137
rect 162122 5063 162124 5072
rect 162176 5063 162178 5072
rect 162124 5034 162176 5040
rect 162032 4480 162084 4486
rect 162032 4422 162084 4428
rect 161940 3732 161992 3738
rect 161940 3674 161992 3680
rect 161662 3632 161718 3641
rect 161662 3567 161718 3576
rect 160940 2746 161244 2774
rect 161492 2746 161612 2774
rect 160744 2644 160796 2650
rect 160744 2586 160796 2592
rect 160928 2304 160980 2310
rect 160928 2246 160980 2252
rect 160940 1193 160968 2246
rect 161216 1970 161244 2746
rect 161388 2644 161440 2650
rect 161388 2586 161440 2592
rect 161204 1964 161256 1970
rect 161204 1906 161256 1912
rect 161400 1290 161428 2586
rect 161584 1970 161612 2746
rect 161676 2378 161704 3567
rect 161952 2417 161980 3674
rect 162044 3058 162072 4422
rect 162032 3052 162084 3058
rect 162032 2994 162084 3000
rect 161938 2408 161994 2417
rect 161664 2372 161716 2378
rect 161938 2343 161994 2352
rect 161664 2314 161716 2320
rect 161756 2304 161808 2310
rect 161756 2246 161808 2252
rect 162124 2304 162176 2310
rect 162124 2246 162176 2252
rect 161572 1964 161624 1970
rect 161572 1906 161624 1912
rect 161480 1760 161532 1766
rect 161480 1702 161532 1708
rect 161492 1358 161520 1702
rect 161480 1352 161532 1358
rect 161480 1294 161532 1300
rect 161388 1284 161440 1290
rect 161388 1226 161440 1232
rect 161296 1216 161348 1222
rect 160926 1184 160982 1193
rect 161768 1193 161796 2246
rect 162136 2106 162164 2246
rect 162124 2100 162176 2106
rect 162124 2042 162176 2048
rect 162228 1970 162256 8366
rect 162320 8090 162348 8463
rect 162676 8434 162728 8440
rect 162582 8392 162638 8401
rect 162582 8327 162638 8336
rect 162400 8288 162452 8294
rect 162400 8230 162452 8236
rect 162308 8084 162360 8090
rect 162308 8026 162360 8032
rect 162412 7410 162440 8230
rect 162596 7546 162624 8327
rect 162688 7954 162716 8434
rect 162780 8430 162808 9454
rect 163412 9172 163464 9178
rect 163412 9114 163464 9120
rect 162768 8424 162820 8430
rect 162768 8366 162820 8372
rect 162860 8356 162912 8362
rect 162860 8298 162912 8304
rect 162872 8022 162900 8298
rect 163320 8288 163372 8294
rect 163320 8230 163372 8236
rect 162860 8016 162912 8022
rect 162860 7958 162912 7964
rect 162952 8016 163004 8022
rect 162952 7958 163004 7964
rect 162676 7948 162728 7954
rect 162676 7890 162728 7896
rect 162688 7546 162716 7890
rect 162584 7540 162636 7546
rect 162584 7482 162636 7488
rect 162676 7540 162728 7546
rect 162676 7482 162728 7488
rect 162400 7404 162452 7410
rect 162400 7346 162452 7352
rect 162964 7342 162992 7958
rect 162952 7336 163004 7342
rect 162952 7278 163004 7284
rect 162676 6656 162728 6662
rect 162676 6598 162728 6604
rect 162492 6452 162544 6458
rect 162492 6394 162544 6400
rect 162584 6452 162636 6458
rect 162584 6394 162636 6400
rect 162504 4146 162532 6394
rect 162596 6254 162624 6394
rect 162584 6248 162636 6254
rect 162584 6190 162636 6196
rect 162584 5568 162636 5574
rect 162584 5510 162636 5516
rect 162596 5302 162624 5510
rect 162584 5296 162636 5302
rect 162584 5238 162636 5244
rect 162688 5166 162716 6598
rect 162860 6384 162912 6390
rect 162766 6352 162822 6361
rect 162860 6326 162912 6332
rect 162766 6287 162822 6296
rect 162780 5914 162808 6287
rect 162872 6254 162900 6326
rect 162860 6248 162912 6254
rect 162860 6190 162912 6196
rect 162768 5908 162820 5914
rect 162768 5850 162820 5856
rect 163044 5908 163096 5914
rect 163044 5850 163096 5856
rect 162780 5642 162808 5850
rect 162768 5636 162820 5642
rect 162768 5578 162820 5584
rect 163056 5370 163084 5850
rect 163044 5364 163096 5370
rect 163044 5306 163096 5312
rect 163228 5364 163280 5370
rect 163228 5306 163280 5312
rect 162676 5160 162728 5166
rect 162676 5102 162728 5108
rect 163134 5128 163190 5137
rect 162492 4140 162544 4146
rect 162492 4082 162544 4088
rect 162688 3670 162716 5102
rect 163134 5063 163190 5072
rect 162952 5024 163004 5030
rect 162952 4966 163004 4972
rect 162676 3664 162728 3670
rect 162676 3606 162728 3612
rect 162492 3528 162544 3534
rect 162492 3470 162544 3476
rect 162308 2440 162360 2446
rect 162308 2382 162360 2388
rect 162320 2106 162348 2382
rect 162504 2310 162532 3470
rect 162676 3460 162728 3466
rect 162676 3402 162728 3408
rect 162688 3126 162716 3402
rect 162676 3120 162728 3126
rect 162676 3062 162728 3068
rect 162964 3058 162992 4966
rect 163148 4554 163176 5063
rect 163240 4826 163268 5306
rect 163228 4820 163280 4826
rect 163228 4762 163280 4768
rect 163136 4548 163188 4554
rect 163136 4490 163188 4496
rect 162952 3052 163004 3058
rect 162952 2994 163004 3000
rect 163136 2848 163188 2854
rect 163136 2790 163188 2796
rect 162492 2304 162544 2310
rect 162492 2246 162544 2252
rect 162308 2100 162360 2106
rect 162308 2042 162360 2048
rect 162216 1964 162268 1970
rect 162216 1906 162268 1912
rect 163148 1902 163176 2790
rect 163136 1896 163188 1902
rect 163136 1838 163188 1844
rect 163136 1760 163188 1766
rect 163136 1702 163188 1708
rect 163148 1358 163176 1702
rect 163136 1352 163188 1358
rect 163136 1294 163188 1300
rect 162492 1216 162544 1222
rect 161296 1158 161348 1164
rect 161754 1184 161810 1193
rect 160926 1119 160982 1128
rect 161308 649 161336 1158
rect 162492 1158 162544 1164
rect 161754 1119 161810 1128
rect 162504 649 162532 1158
rect 161294 640 161350 649
rect 161294 575 161350 584
rect 162490 640 162546 649
rect 162490 575 162546 584
rect 160468 468 160520 474
rect 160468 410 160520 416
rect 163332 377 163360 8230
rect 163424 3466 163452 9114
rect 163504 6724 163556 6730
rect 163504 6666 163556 6672
rect 163516 5234 163544 6666
rect 163504 5228 163556 5234
rect 163504 5170 163556 5176
rect 163412 3460 163464 3466
rect 163412 3402 163464 3408
rect 163608 2553 163636 9862
rect 163700 8498 163728 9998
rect 163870 9752 163926 9761
rect 163870 9687 163872 9696
rect 163924 9687 163926 9696
rect 163872 9658 163924 9664
rect 163872 8900 163924 8906
rect 163792 8860 163872 8888
rect 163688 8492 163740 8498
rect 163688 8434 163740 8440
rect 163792 7886 163820 8860
rect 163872 8842 163924 8848
rect 163976 8430 164004 10814
rect 164148 10804 164200 10810
rect 164148 10746 164200 10752
rect 164332 10804 164384 10810
rect 164332 10746 164384 10752
rect 164160 8906 164188 10746
rect 164344 9586 164372 10746
rect 164608 10736 164660 10742
rect 164608 10678 164660 10684
rect 164792 10736 164844 10742
rect 164792 10678 164844 10684
rect 164332 9580 164384 9586
rect 164332 9522 164384 9528
rect 164620 9518 164648 10678
rect 164608 9512 164660 9518
rect 164608 9454 164660 9460
rect 164148 8900 164200 8906
rect 164148 8842 164200 8848
rect 164240 8832 164292 8838
rect 164240 8774 164292 8780
rect 163964 8424 164016 8430
rect 164148 8424 164200 8430
rect 163964 8366 164016 8372
rect 164054 8392 164110 8401
rect 164148 8366 164200 8372
rect 164054 8327 164110 8336
rect 163780 7880 163832 7886
rect 163780 7822 163832 7828
rect 163686 7304 163742 7313
rect 163686 7239 163742 7248
rect 163700 4078 163728 7239
rect 163688 4072 163740 4078
rect 163688 4014 163740 4020
rect 163792 2774 163820 7822
rect 163872 7744 163924 7750
rect 163872 7686 163924 7692
rect 163884 7410 163912 7686
rect 164068 7546 164096 8327
rect 164056 7540 164108 7546
rect 164056 7482 164108 7488
rect 163872 7404 163924 7410
rect 163872 7346 163924 7352
rect 163700 2746 163820 2774
rect 163594 2544 163650 2553
rect 163594 2479 163650 2488
rect 163410 2408 163466 2417
rect 163410 2343 163466 2352
rect 163424 2009 163452 2343
rect 163410 2000 163466 2009
rect 163700 1970 163728 2746
rect 163964 2440 164016 2446
rect 163964 2382 164016 2388
rect 163872 2304 163924 2310
rect 163872 2246 163924 2252
rect 163410 1935 163466 1944
rect 163688 1964 163740 1970
rect 163688 1906 163740 1912
rect 163780 1964 163832 1970
rect 163780 1906 163832 1912
rect 163792 1358 163820 1906
rect 163780 1352 163832 1358
rect 163780 1294 163832 1300
rect 163884 1193 163912 2246
rect 163976 2106 164004 2382
rect 163964 2100 164016 2106
rect 163964 2042 164016 2048
rect 164160 1426 164188 8366
rect 164252 5098 164280 8774
rect 164620 7886 164648 9454
rect 164804 9178 164832 10678
rect 165344 10668 165396 10674
rect 165344 10610 165396 10616
rect 165252 9988 165304 9994
rect 165252 9930 165304 9936
rect 165160 9580 165212 9586
rect 165160 9522 165212 9528
rect 164792 9172 164844 9178
rect 164712 9132 164792 9160
rect 164712 8974 164740 9132
rect 164792 9114 164844 9120
rect 164700 8968 164752 8974
rect 164700 8910 164752 8916
rect 165172 8634 165200 9522
rect 165264 8974 165292 9930
rect 165356 9042 165384 10610
rect 167092 10600 167144 10606
rect 167092 10542 167144 10548
rect 196716 10600 196768 10606
rect 196716 10542 196768 10548
rect 208306 10568 208362 10577
rect 166264 10260 166316 10266
rect 166264 10202 166316 10208
rect 165804 9648 165856 9654
rect 165804 9590 165856 9596
rect 165528 9580 165580 9586
rect 165528 9522 165580 9528
rect 165344 9036 165396 9042
rect 165344 8978 165396 8984
rect 165252 8968 165304 8974
rect 165252 8910 165304 8916
rect 165160 8628 165212 8634
rect 165160 8570 165212 8576
rect 164790 8392 164846 8401
rect 164790 8327 164846 8336
rect 164332 7880 164384 7886
rect 164332 7822 164384 7828
rect 164608 7880 164660 7886
rect 164608 7822 164660 7828
rect 164240 5092 164292 5098
rect 164240 5034 164292 5040
rect 164240 2304 164292 2310
rect 164240 2246 164292 2252
rect 164252 1465 164280 2246
rect 164344 1970 164372 7822
rect 164608 7744 164660 7750
rect 164608 7686 164660 7692
rect 164620 7410 164648 7686
rect 164804 7546 164832 8327
rect 165356 7886 165384 8978
rect 165540 8498 165568 9522
rect 165816 9382 165844 9590
rect 166276 9518 166304 10202
rect 167104 9518 167132 10542
rect 167736 10532 167788 10538
rect 167736 10474 167788 10480
rect 192484 10532 192536 10538
rect 192484 10474 192536 10480
rect 166264 9512 166316 9518
rect 166264 9454 166316 9460
rect 167092 9512 167144 9518
rect 167092 9454 167144 9460
rect 167552 9512 167604 9518
rect 167552 9454 167604 9460
rect 165804 9376 165856 9382
rect 165804 9318 165856 9324
rect 166172 9376 166224 9382
rect 166172 9318 166224 9324
rect 165528 8492 165580 8498
rect 165448 8452 165528 8480
rect 165448 7886 165476 8452
rect 165528 8434 165580 8440
rect 165526 8392 165582 8401
rect 165526 8327 165582 8336
rect 165344 7880 165396 7886
rect 165264 7828 165344 7834
rect 165264 7822 165396 7828
rect 165436 7880 165488 7886
rect 165436 7822 165488 7828
rect 165264 7806 165384 7822
rect 164792 7540 164844 7546
rect 164792 7482 164844 7488
rect 164608 7404 164660 7410
rect 164608 7346 164660 7352
rect 165160 7336 165212 7342
rect 165160 7278 165212 7284
rect 165172 7002 165200 7278
rect 165160 6996 165212 7002
rect 165160 6938 165212 6944
rect 164424 2440 164476 2446
rect 164424 2382 164476 2388
rect 164332 1964 164384 1970
rect 164332 1906 164384 1912
rect 164238 1456 164294 1465
rect 164148 1420 164200 1426
rect 164238 1391 164294 1400
rect 164148 1362 164200 1368
rect 164436 1358 164464 2382
rect 165264 1970 165292 7806
rect 165344 7744 165396 7750
rect 165344 7686 165396 7692
rect 165356 7410 165384 7686
rect 165540 7546 165568 8327
rect 165620 7948 165672 7954
rect 165620 7890 165672 7896
rect 165528 7540 165580 7546
rect 165528 7482 165580 7488
rect 165344 7404 165396 7410
rect 165344 7346 165396 7352
rect 165632 7206 165660 7890
rect 166184 7886 166212 9318
rect 166276 8906 166304 9454
rect 166264 8900 166316 8906
rect 166264 8842 166316 8848
rect 166172 7880 166224 7886
rect 166172 7822 166224 7828
rect 165620 7200 165672 7206
rect 165620 7142 165672 7148
rect 165620 2440 165672 2446
rect 165620 2382 165672 2388
rect 165896 2440 165948 2446
rect 165896 2382 165948 2388
rect 165344 2304 165396 2310
rect 165344 2246 165396 2252
rect 165252 1964 165304 1970
rect 165252 1906 165304 1912
rect 164516 1760 164568 1766
rect 164516 1702 164568 1708
rect 164528 1358 164556 1702
rect 164424 1352 164476 1358
rect 164424 1294 164476 1300
rect 164516 1352 164568 1358
rect 164516 1294 164568 1300
rect 164700 1216 164752 1222
rect 163870 1184 163926 1193
rect 165356 1193 165384 2246
rect 165632 2106 165660 2382
rect 165908 2106 165936 2382
rect 166080 2304 166132 2310
rect 166080 2246 166132 2252
rect 165620 2100 165672 2106
rect 165620 2042 165672 2048
rect 165896 2100 165948 2106
rect 165896 2042 165948 2048
rect 166092 1193 166120 2246
rect 166276 1970 166304 8842
rect 167104 8430 167132 9454
rect 167460 9376 167512 9382
rect 167460 9318 167512 9324
rect 167368 8900 167420 8906
rect 167368 8842 167420 8848
rect 167380 8498 167408 8842
rect 167368 8492 167420 8498
rect 167368 8434 167420 8440
rect 167092 8424 167144 8430
rect 166354 8392 166410 8401
rect 167092 8366 167144 8372
rect 166354 8327 166410 8336
rect 166368 8090 166396 8327
rect 166814 8256 166870 8265
rect 166814 8191 166870 8200
rect 166828 8090 166856 8191
rect 166356 8084 166408 8090
rect 166356 8026 166408 8032
rect 166816 8084 166868 8090
rect 166816 8026 166868 8032
rect 166816 2304 166868 2310
rect 166816 2246 166868 2252
rect 166264 1964 166316 1970
rect 166264 1906 166316 1912
rect 166828 1193 166856 2246
rect 167104 1970 167132 8366
rect 167472 7886 167500 9318
rect 167564 8838 167592 9454
rect 167748 8974 167776 10474
rect 181810 10432 181866 10441
rect 191286 10432 191342 10441
rect 181810 10367 181866 10376
rect 181996 10396 182048 10402
rect 172520 10328 172572 10334
rect 171690 10296 171746 10305
rect 170312 10260 170364 10266
rect 171690 10231 171746 10240
rect 172334 10296 172390 10305
rect 172520 10270 172572 10276
rect 173070 10296 173126 10305
rect 172334 10231 172390 10240
rect 170312 10202 170364 10208
rect 168104 9580 168156 9586
rect 168104 9522 168156 9528
rect 169300 9580 169352 9586
rect 169300 9522 169352 9528
rect 167920 9512 167972 9518
rect 167920 9454 167972 9460
rect 167736 8968 167788 8974
rect 167736 8910 167788 8916
rect 167552 8832 167604 8838
rect 167552 8774 167604 8780
rect 167644 8832 167696 8838
rect 167644 8774 167696 8780
rect 167656 7886 167684 8774
rect 167748 8430 167776 8910
rect 167736 8424 167788 8430
rect 167736 8366 167788 8372
rect 167826 8392 167882 8401
rect 167826 8327 167882 8336
rect 167840 8090 167868 8327
rect 167828 8084 167880 8090
rect 167828 8026 167880 8032
rect 167460 7880 167512 7886
rect 167460 7822 167512 7828
rect 167644 7880 167696 7886
rect 167644 7822 167696 7828
rect 167736 2984 167788 2990
rect 167736 2926 167788 2932
rect 167748 2446 167776 2926
rect 167460 2440 167512 2446
rect 167460 2382 167512 2388
rect 167736 2440 167788 2446
rect 167736 2382 167788 2388
rect 167828 2440 167880 2446
rect 167828 2382 167880 2388
rect 167472 2106 167500 2382
rect 167552 2372 167604 2378
rect 167552 2314 167604 2320
rect 167564 2106 167592 2314
rect 167460 2100 167512 2106
rect 167460 2042 167512 2048
rect 167552 2100 167604 2106
rect 167552 2042 167604 2048
rect 167092 1964 167144 1970
rect 167092 1906 167144 1912
rect 167840 1902 167868 2382
rect 167932 1970 167960 9454
rect 168116 8974 168144 9522
rect 168288 9512 168340 9518
rect 168288 9454 168340 9460
rect 169116 9512 169168 9518
rect 169116 9454 169168 9460
rect 168300 8974 168328 9454
rect 168840 9376 168892 9382
rect 168840 9318 168892 9324
rect 168104 8968 168156 8974
rect 168104 8910 168156 8916
rect 168288 8968 168340 8974
rect 168288 8910 168340 8916
rect 168104 8424 168156 8430
rect 168104 8366 168156 8372
rect 168012 2304 168064 2310
rect 168012 2246 168064 2252
rect 167920 1964 167972 1970
rect 167920 1906 167972 1912
rect 167184 1896 167236 1902
rect 167184 1838 167236 1844
rect 167828 1896 167880 1902
rect 167828 1838 167880 1844
rect 167196 1358 167224 1838
rect 168024 1358 168052 2246
rect 168116 1426 168144 8366
rect 168378 8120 168434 8129
rect 168378 8055 168380 8064
rect 168432 8055 168434 8064
rect 168380 8026 168432 8032
rect 168852 7886 168880 9318
rect 169022 9208 169078 9217
rect 169022 9143 169024 9152
rect 169076 9143 169078 9152
rect 169024 9114 169076 9120
rect 168840 7880 168892 7886
rect 168840 7822 168892 7828
rect 168288 7540 168340 7546
rect 168288 7482 168340 7488
rect 168196 7472 168248 7478
rect 168196 7414 168248 7420
rect 168208 2378 168236 7414
rect 168300 6458 168328 7482
rect 169128 7206 169156 9454
rect 169116 7200 169168 7206
rect 169116 7142 169168 7148
rect 169128 7002 169156 7142
rect 169116 6996 169168 7002
rect 169116 6938 169168 6944
rect 169208 6792 169260 6798
rect 169208 6734 169260 6740
rect 168288 6452 168340 6458
rect 168288 6394 168340 6400
rect 169220 6186 169248 6734
rect 169208 6180 169260 6186
rect 169208 6122 169260 6128
rect 169312 6118 169340 9522
rect 169760 9512 169812 9518
rect 169760 9454 169812 9460
rect 169772 8498 169800 9454
rect 169942 9276 170250 9285
rect 169942 9274 169948 9276
rect 170004 9274 170028 9276
rect 170084 9274 170108 9276
rect 170164 9274 170188 9276
rect 170244 9274 170250 9276
rect 170004 9222 170006 9274
rect 170186 9222 170188 9274
rect 169942 9220 169948 9222
rect 170004 9220 170028 9222
rect 170084 9220 170108 9222
rect 170164 9220 170188 9222
rect 170244 9220 170250 9222
rect 169942 9211 170250 9220
rect 169852 8968 169904 8974
rect 169852 8910 169904 8916
rect 169944 8968 169996 8974
rect 169944 8910 169996 8916
rect 169864 8838 169892 8910
rect 169852 8832 169904 8838
rect 169852 8774 169904 8780
rect 169956 8634 169984 8910
rect 170324 8838 170352 10202
rect 170588 9648 170640 9654
rect 170588 9590 170640 9596
rect 170600 9178 170628 9590
rect 171704 9586 171732 10231
rect 172348 9654 172376 10231
rect 172532 9654 172560 10270
rect 173070 10231 173126 10240
rect 173714 10296 173770 10305
rect 173714 10231 173770 10240
rect 174450 10296 174506 10305
rect 174450 10231 174506 10240
rect 175186 10296 175242 10305
rect 175186 10231 175242 10240
rect 175922 10296 175978 10305
rect 175922 10231 175978 10240
rect 176750 10296 176806 10305
rect 176750 10231 176806 10240
rect 177486 10296 177542 10305
rect 177486 10231 177542 10240
rect 177946 10296 178002 10305
rect 177946 10231 178002 10240
rect 179142 10296 179198 10305
rect 179142 10231 179198 10240
rect 179602 10296 179658 10305
rect 179602 10231 179658 10240
rect 180338 10296 180394 10305
rect 180338 10231 180394 10240
rect 181718 10296 181774 10305
rect 181718 10231 181774 10240
rect 173084 9654 173112 10231
rect 172336 9648 172388 9654
rect 172336 9590 172388 9596
rect 172520 9648 172572 9654
rect 172520 9590 172572 9596
rect 173072 9648 173124 9654
rect 173072 9590 173124 9596
rect 171692 9580 171744 9586
rect 171692 9522 171744 9528
rect 173164 9376 173216 9382
rect 173164 9318 173216 9324
rect 170588 9172 170640 9178
rect 170588 9114 170640 9120
rect 170312 8832 170364 8838
rect 170312 8774 170364 8780
rect 169944 8628 169996 8634
rect 169944 8570 169996 8576
rect 170036 8628 170088 8634
rect 170036 8570 170088 8576
rect 169760 8492 169812 8498
rect 169760 8434 169812 8440
rect 169576 8424 169628 8430
rect 169576 8366 169628 8372
rect 169588 7954 169616 8366
rect 170048 8362 170076 8570
rect 170036 8356 170088 8362
rect 170036 8298 170088 8304
rect 169942 8188 170250 8197
rect 169942 8186 169948 8188
rect 170004 8186 170028 8188
rect 170084 8186 170108 8188
rect 170164 8186 170188 8188
rect 170244 8186 170250 8188
rect 170004 8134 170006 8186
rect 170186 8134 170188 8186
rect 169942 8132 169948 8134
rect 170004 8132 170028 8134
rect 170084 8132 170108 8134
rect 170164 8132 170188 8134
rect 170244 8132 170250 8134
rect 169942 8123 170250 8132
rect 169576 7948 169628 7954
rect 169576 7890 169628 7896
rect 169760 7404 169812 7410
rect 169760 7346 169812 7352
rect 169772 6934 169800 7346
rect 172520 7336 172572 7342
rect 172520 7278 172572 7284
rect 169942 7100 170250 7109
rect 169942 7098 169948 7100
rect 170004 7098 170028 7100
rect 170084 7098 170108 7100
rect 170164 7098 170188 7100
rect 170244 7098 170250 7100
rect 170004 7046 170006 7098
rect 170186 7046 170188 7098
rect 169942 7044 169948 7046
rect 170004 7044 170028 7046
rect 170084 7044 170108 7046
rect 170164 7044 170188 7046
rect 170244 7044 170250 7046
rect 169942 7035 170250 7044
rect 169760 6928 169812 6934
rect 169760 6870 169812 6876
rect 172532 6798 172560 7278
rect 172520 6792 172572 6798
rect 172520 6734 172572 6740
rect 170586 6352 170642 6361
rect 170586 6287 170642 6296
rect 169300 6112 169352 6118
rect 169300 6054 169352 6060
rect 169942 6012 170250 6021
rect 169942 6010 169948 6012
rect 170004 6010 170028 6012
rect 170084 6010 170108 6012
rect 170164 6010 170188 6012
rect 170244 6010 170250 6012
rect 170004 5958 170006 6010
rect 170186 5958 170188 6010
rect 169942 5956 169948 5958
rect 170004 5956 170028 5958
rect 170084 5956 170108 5958
rect 170164 5956 170188 5958
rect 170244 5956 170250 5958
rect 169942 5947 170250 5956
rect 170600 5817 170628 6287
rect 170586 5808 170642 5817
rect 170586 5743 170642 5752
rect 169942 4924 170250 4933
rect 169942 4922 169948 4924
rect 170004 4922 170028 4924
rect 170084 4922 170108 4924
rect 170164 4922 170188 4924
rect 170244 4922 170250 4924
rect 170004 4870 170006 4922
rect 170186 4870 170188 4922
rect 169942 4868 169948 4870
rect 170004 4868 170028 4870
rect 170084 4868 170108 4870
rect 170164 4868 170188 4870
rect 170244 4868 170250 4870
rect 169942 4859 170250 4868
rect 169942 3836 170250 3845
rect 169942 3834 169948 3836
rect 170004 3834 170028 3836
rect 170084 3834 170108 3836
rect 170164 3834 170188 3836
rect 170244 3834 170250 3836
rect 170004 3782 170006 3834
rect 170186 3782 170188 3834
rect 169942 3780 169948 3782
rect 170004 3780 170028 3782
rect 170084 3780 170108 3782
rect 170164 3780 170188 3782
rect 170244 3780 170250 3782
rect 169942 3771 170250 3780
rect 173176 3738 173204 9318
rect 173728 8974 173756 10231
rect 174464 9586 174492 10231
rect 175200 9654 175228 10231
rect 175936 9654 175964 10231
rect 175188 9648 175240 9654
rect 175188 9590 175240 9596
rect 175924 9648 175976 9654
rect 175924 9590 175976 9596
rect 174452 9580 174504 9586
rect 174452 9522 174504 9528
rect 174728 9512 174780 9518
rect 174728 9454 174780 9460
rect 173716 8968 173768 8974
rect 173716 8910 173768 8916
rect 174176 8832 174228 8838
rect 174176 8774 174228 8780
rect 173440 8492 173492 8498
rect 173440 8434 173492 8440
rect 173452 7993 173480 8434
rect 173438 7984 173494 7993
rect 173438 7919 173494 7928
rect 173806 4448 173862 4457
rect 173806 4383 173862 4392
rect 173164 3732 173216 3738
rect 173164 3674 173216 3680
rect 169942 2748 170250 2757
rect 169942 2746 169948 2748
rect 170004 2746 170028 2748
rect 170084 2746 170108 2748
rect 170164 2746 170188 2748
rect 170244 2746 170250 2748
rect 170004 2694 170006 2746
rect 170186 2694 170188 2746
rect 169942 2692 169948 2694
rect 170004 2692 170028 2694
rect 170084 2692 170108 2694
rect 170164 2692 170188 2694
rect 170244 2692 170250 2694
rect 169942 2683 170250 2692
rect 173254 2408 173310 2417
rect 168196 2372 168248 2378
rect 173254 2343 173310 2352
rect 168196 2314 168248 2320
rect 173268 1970 173296 2343
rect 173820 2310 173848 4383
rect 174188 3369 174216 8774
rect 174740 7818 174768 9454
rect 175924 9376 175976 9382
rect 175924 9318 175976 9324
rect 174728 7812 174780 7818
rect 174728 7754 174780 7760
rect 175936 5370 175964 9318
rect 176764 8906 176792 10231
rect 177212 9036 177264 9042
rect 177212 8978 177264 8984
rect 176752 8900 176804 8906
rect 176752 8842 176804 8848
rect 176844 8832 176896 8838
rect 176844 8774 176896 8780
rect 176856 7585 176884 8774
rect 177224 7886 177252 8978
rect 177500 8974 177528 10231
rect 177960 9586 177988 10231
rect 179156 9586 179184 10231
rect 177948 9580 178000 9586
rect 177948 9522 178000 9528
rect 179144 9580 179196 9586
rect 179144 9522 179196 9528
rect 178040 9512 178092 9518
rect 178040 9454 178092 9460
rect 177948 9376 178000 9382
rect 177948 9318 178000 9324
rect 177488 8968 177540 8974
rect 177488 8910 177540 8916
rect 177580 8832 177632 8838
rect 177580 8774 177632 8780
rect 177856 8832 177908 8838
rect 177856 8774 177908 8780
rect 177212 7880 177264 7886
rect 177212 7822 177264 7828
rect 176842 7576 176898 7585
rect 176842 7511 176898 7520
rect 177026 6352 177082 6361
rect 177026 6287 177082 6296
rect 177040 5574 177068 6287
rect 177028 5568 177080 5574
rect 177028 5510 177080 5516
rect 177592 5409 177620 8774
rect 177868 6390 177896 8774
rect 177960 7857 177988 9318
rect 177946 7848 178002 7857
rect 177946 7783 178002 7792
rect 178052 7721 178080 9454
rect 179616 9042 179644 10231
rect 179972 9716 180024 9722
rect 179972 9658 180024 9664
rect 179604 9036 179656 9042
rect 179604 8978 179656 8984
rect 179880 8968 179932 8974
rect 179880 8910 179932 8916
rect 178038 7712 178094 7721
rect 178038 7647 178094 7656
rect 177946 7168 178002 7177
rect 177946 7103 178002 7112
rect 177960 6633 177988 7103
rect 177946 6624 178002 6633
rect 177946 6559 178002 6568
rect 177856 6384 177908 6390
rect 177856 6326 177908 6332
rect 177948 5568 178000 5574
rect 177948 5510 178000 5516
rect 177578 5400 177634 5409
rect 175924 5364 175976 5370
rect 177578 5335 177634 5344
rect 175924 5306 175976 5312
rect 177960 5166 177988 5510
rect 177948 5160 178000 5166
rect 177948 5102 178000 5108
rect 175832 5092 175884 5098
rect 175832 5034 175884 5040
rect 174174 3360 174230 3369
rect 174174 3295 174230 3304
rect 174728 2372 174780 2378
rect 174728 2314 174780 2320
rect 173808 2304 173860 2310
rect 173808 2246 173860 2252
rect 174740 1970 174768 2314
rect 173256 1964 173308 1970
rect 173256 1906 173308 1912
rect 174728 1964 174780 1970
rect 174728 1906 174780 1912
rect 172980 1896 173032 1902
rect 172980 1838 173032 1844
rect 174452 1896 174504 1902
rect 174452 1838 174504 1844
rect 168380 1760 168432 1766
rect 168380 1702 168432 1708
rect 168392 1465 168420 1702
rect 169942 1660 170250 1669
rect 169942 1658 169948 1660
rect 170004 1658 170028 1660
rect 170084 1658 170108 1660
rect 170164 1658 170188 1660
rect 170244 1658 170250 1660
rect 170004 1606 170006 1658
rect 170186 1606 170188 1658
rect 169942 1604 169948 1606
rect 170004 1604 170028 1606
rect 170084 1604 170108 1606
rect 170164 1604 170188 1606
rect 170244 1604 170250 1606
rect 169942 1595 170250 1604
rect 168378 1456 168434 1465
rect 168104 1420 168156 1426
rect 168378 1391 168434 1400
rect 171692 1420 171744 1426
rect 168104 1362 168156 1368
rect 171692 1362 171744 1368
rect 167184 1352 167236 1358
rect 167184 1294 167236 1300
rect 168012 1352 168064 1358
rect 168012 1294 168064 1300
rect 169298 1320 169354 1329
rect 169298 1255 169354 1264
rect 168012 1216 168064 1222
rect 164700 1158 164752 1164
rect 165342 1184 165398 1193
rect 163870 1119 163926 1128
rect 164712 649 164740 1158
rect 165342 1119 165398 1128
rect 166078 1184 166134 1193
rect 166078 1119 166134 1128
rect 166814 1184 166870 1193
rect 168012 1158 168064 1164
rect 169024 1216 169076 1222
rect 169024 1158 169076 1164
rect 166814 1119 166870 1128
rect 168024 649 168052 1158
rect 169036 649 169064 1158
rect 169312 785 169340 1255
rect 171414 1184 171470 1193
rect 171414 1119 171470 1128
rect 171428 921 171456 1119
rect 171704 921 171732 1362
rect 172244 1352 172296 1358
rect 172244 1294 172296 1300
rect 172520 1352 172572 1358
rect 172520 1294 172572 1300
rect 172256 921 172284 1294
rect 171414 912 171470 921
rect 171414 847 171470 856
rect 171690 912 171746 921
rect 171690 847 171746 856
rect 172242 912 172298 921
rect 172242 847 172298 856
rect 169298 776 169354 785
rect 169298 711 169354 720
rect 164698 640 164754 649
rect 164698 575 164754 584
rect 168010 640 168066 649
rect 168010 575 168066 584
rect 169022 640 169078 649
rect 172532 610 172560 1294
rect 172992 921 173020 1838
rect 173808 1352 173860 1358
rect 173808 1294 173860 1300
rect 174268 1352 174320 1358
rect 174268 1294 174320 1300
rect 173820 921 173848 1294
rect 174280 1018 174308 1294
rect 174268 1012 174320 1018
rect 174268 954 174320 960
rect 174464 921 174492 1838
rect 175844 1562 175872 5034
rect 179892 4826 179920 8910
rect 179984 8430 180012 9658
rect 180352 9042 180380 10231
rect 181732 9586 181760 10231
rect 181720 9580 181772 9586
rect 181720 9522 181772 9528
rect 181824 9042 181852 10367
rect 191286 10367 191342 10376
rect 181996 10338 182048 10344
rect 182008 9586 182036 10338
rect 182546 10296 182602 10305
rect 182546 10231 182602 10240
rect 183282 10296 183338 10305
rect 183282 10231 183338 10240
rect 184294 10296 184350 10305
rect 184294 10231 184350 10240
rect 184754 10296 184810 10305
rect 184754 10231 184810 10240
rect 185490 10296 185546 10305
rect 185490 10231 185546 10240
rect 186226 10296 186282 10305
rect 186226 10231 186282 10240
rect 186962 10296 187018 10305
rect 186962 10231 187018 10240
rect 187698 10296 187754 10305
rect 187698 10231 187754 10240
rect 188434 10296 188490 10305
rect 188434 10231 188490 10240
rect 189446 10296 189502 10305
rect 189446 10231 189502 10240
rect 189906 10296 189962 10305
rect 189906 10231 189962 10240
rect 182456 10124 182508 10130
rect 182456 10066 182508 10072
rect 181996 9580 182048 9586
rect 181996 9522 182048 9528
rect 182468 9042 182496 10066
rect 182560 9586 182588 10231
rect 182548 9580 182600 9586
rect 182548 9522 182600 9528
rect 180340 9036 180392 9042
rect 180340 8978 180392 8984
rect 181812 9036 181864 9042
rect 181812 8978 181864 8984
rect 182456 9036 182508 9042
rect 182456 8978 182508 8984
rect 181168 8968 181220 8974
rect 181168 8910 181220 8916
rect 179972 8424 180024 8430
rect 179972 8366 180024 8372
rect 181180 7274 181208 8910
rect 183296 8498 183324 10231
rect 184308 9042 184336 10231
rect 184572 9512 184624 9518
rect 184572 9454 184624 9460
rect 184584 9110 184612 9454
rect 184572 9104 184624 9110
rect 184572 9046 184624 9052
rect 184768 9042 184796 10231
rect 185504 9586 185532 10231
rect 185492 9580 185544 9586
rect 185492 9522 185544 9528
rect 185952 9444 186004 9450
rect 185952 9386 186004 9392
rect 184296 9036 184348 9042
rect 184296 8978 184348 8984
rect 184756 9036 184808 9042
rect 184756 8978 184808 8984
rect 184572 8968 184624 8974
rect 184572 8910 184624 8916
rect 185860 8968 185912 8974
rect 185860 8910 185912 8916
rect 183284 8492 183336 8498
rect 183284 8434 183336 8440
rect 184584 8022 184612 8910
rect 185872 8634 185900 8910
rect 185964 8634 185992 9386
rect 186240 9042 186268 10231
rect 186228 9036 186280 9042
rect 186228 8978 186280 8984
rect 185860 8628 185912 8634
rect 185860 8570 185912 8576
rect 185952 8628 186004 8634
rect 185952 8570 186004 8576
rect 186976 8498 187004 10231
rect 187056 9920 187108 9926
rect 187056 9862 187108 9868
rect 187068 8498 187096 9862
rect 187712 9586 187740 10231
rect 187700 9580 187752 9586
rect 187700 9522 187752 9528
rect 187240 8968 187292 8974
rect 187240 8910 187292 8916
rect 186964 8492 187016 8498
rect 186964 8434 187016 8440
rect 187056 8492 187108 8498
rect 187056 8434 187108 8440
rect 184572 8016 184624 8022
rect 184572 7958 184624 7964
rect 187252 7954 187280 8910
rect 187700 8560 187752 8566
rect 187700 8502 187752 8508
rect 187712 8129 187740 8502
rect 188448 8498 188476 10231
rect 189460 9042 189488 10231
rect 189724 9512 189776 9518
rect 189724 9454 189776 9460
rect 189736 9178 189764 9454
rect 189724 9172 189776 9178
rect 189724 9114 189776 9120
rect 189448 9036 189500 9042
rect 189448 8978 189500 8984
rect 189920 8634 189948 10231
rect 190000 9580 190052 9586
rect 190000 9522 190052 9528
rect 190828 9580 190880 9586
rect 190828 9522 190880 9528
rect 189908 8628 189960 8634
rect 189908 8570 189960 8576
rect 188436 8492 188488 8498
rect 188436 8434 188488 8440
rect 187698 8120 187754 8129
rect 187698 8055 187754 8064
rect 187240 7948 187292 7954
rect 187240 7890 187292 7896
rect 189264 7812 189316 7818
rect 189264 7754 189316 7760
rect 181168 7268 181220 7274
rect 181168 7210 181220 7216
rect 180064 6996 180116 7002
rect 180064 6938 180116 6944
rect 180076 6497 180104 6938
rect 180984 6928 181036 6934
rect 180984 6870 181036 6876
rect 180062 6488 180118 6497
rect 180062 6423 180118 6432
rect 180996 6390 181024 6870
rect 189080 6860 189132 6866
rect 189080 6802 189132 6808
rect 181812 6452 181864 6458
rect 181812 6394 181864 6400
rect 180984 6384 181036 6390
rect 180984 6326 181036 6332
rect 180996 5914 181024 6326
rect 180984 5908 181036 5914
rect 180984 5850 181036 5856
rect 181824 5846 181852 6394
rect 182180 6384 182232 6390
rect 182180 6326 182232 6332
rect 188436 6384 188488 6390
rect 188436 6326 188488 6332
rect 182088 6248 182140 6254
rect 182088 6190 182140 6196
rect 182100 6089 182128 6190
rect 182086 6080 182142 6089
rect 182086 6015 182142 6024
rect 181812 5840 181864 5846
rect 181812 5782 181864 5788
rect 182100 5710 182128 6015
rect 182192 5778 182220 6326
rect 182548 6316 182600 6322
rect 182548 6258 182600 6264
rect 182180 5772 182232 5778
rect 182180 5714 182232 5720
rect 182088 5704 182140 5710
rect 182088 5646 182140 5652
rect 182100 5234 182128 5646
rect 182192 5234 182220 5714
rect 182560 5710 182588 6258
rect 182914 6216 182970 6225
rect 182914 6151 182970 6160
rect 182928 5914 182956 6151
rect 188448 5953 188476 6326
rect 189092 6118 189120 6802
rect 189172 6452 189224 6458
rect 189172 6394 189224 6400
rect 189080 6112 189132 6118
rect 189080 6054 189132 6060
rect 188434 5944 188490 5953
rect 182916 5908 182968 5914
rect 188434 5879 188490 5888
rect 182916 5850 182968 5856
rect 182548 5704 182600 5710
rect 182548 5646 182600 5652
rect 182560 5234 182588 5646
rect 186320 5568 186372 5574
rect 186320 5510 186372 5516
rect 180616 5228 180668 5234
rect 180616 5170 180668 5176
rect 182088 5228 182140 5234
rect 182088 5170 182140 5176
rect 182180 5228 182232 5234
rect 182180 5170 182232 5176
rect 182548 5228 182600 5234
rect 182548 5170 182600 5176
rect 179880 4820 179932 4826
rect 179880 4762 179932 4768
rect 175922 4176 175978 4185
rect 175922 4111 175978 4120
rect 175936 3126 175964 4111
rect 176660 3596 176712 3602
rect 176660 3538 176712 3544
rect 175924 3120 175976 3126
rect 175924 3062 175976 3068
rect 176672 2650 176700 3538
rect 176660 2644 176712 2650
rect 176660 2586 176712 2592
rect 176660 2440 176712 2446
rect 176660 2382 176712 2388
rect 176936 2440 176988 2446
rect 176936 2382 176988 2388
rect 179604 2440 179656 2446
rect 179604 2382 179656 2388
rect 176568 1896 176620 1902
rect 176568 1838 176620 1844
rect 175832 1556 175884 1562
rect 175832 1498 175884 1504
rect 175188 1352 175240 1358
rect 175188 1294 175240 1300
rect 175200 921 175228 1294
rect 176580 921 176608 1838
rect 176672 1329 176700 2382
rect 176842 2136 176898 2145
rect 176842 2071 176898 2080
rect 176856 1970 176884 2071
rect 176844 1964 176896 1970
rect 176844 1906 176896 1912
rect 176948 1494 176976 2382
rect 177856 1896 177908 1902
rect 177856 1838 177908 1844
rect 179144 1896 179196 1902
rect 179144 1838 179196 1844
rect 176936 1488 176988 1494
rect 176936 1430 176988 1436
rect 176844 1352 176896 1358
rect 176658 1320 176714 1329
rect 176844 1294 176896 1300
rect 176658 1255 176714 1264
rect 172978 912 173034 921
rect 172978 847 173034 856
rect 173806 912 173862 921
rect 173806 847 173862 856
rect 174450 912 174506 921
rect 174450 847 174506 856
rect 175186 912 175242 921
rect 175186 847 175242 856
rect 176566 912 176622 921
rect 176566 847 176622 856
rect 176856 678 176884 1294
rect 177868 921 177896 1838
rect 178408 1352 178460 1358
rect 178408 1294 178460 1300
rect 178420 921 178448 1294
rect 179156 921 179184 1838
rect 179512 1828 179564 1834
rect 179512 1770 179564 1776
rect 179420 1352 179472 1358
rect 179420 1294 179472 1300
rect 177854 912 177910 921
rect 177854 847 177910 856
rect 178406 912 178462 921
rect 178406 847 178462 856
rect 179142 912 179198 921
rect 179142 847 179198 856
rect 179432 746 179460 1294
rect 179524 1290 179552 1770
rect 179616 1329 179644 2382
rect 180628 1562 180656 5170
rect 182548 5092 182600 5098
rect 182548 5034 182600 5040
rect 182560 4729 182588 5034
rect 182546 4720 182602 4729
rect 182546 4655 182602 4664
rect 180892 3460 180944 3466
rect 180892 3402 180944 3408
rect 180616 1556 180668 1562
rect 180616 1498 180668 1504
rect 179602 1320 179658 1329
rect 179512 1284 179564 1290
rect 179602 1255 179658 1264
rect 180524 1284 180576 1290
rect 179512 1226 179564 1232
rect 180524 1226 180576 1232
rect 180536 921 180564 1226
rect 180522 912 180578 921
rect 180522 847 180578 856
rect 179420 740 179472 746
rect 179420 682 179472 688
rect 176844 672 176896 678
rect 176844 614 176896 620
rect 169022 575 169078 584
rect 172520 604 172572 610
rect 172520 546 172572 552
rect 154304 342 154356 348
rect 160098 368 160154 377
rect 130842 303 130898 312
rect 160098 303 160154 312
rect 163318 368 163374 377
rect 163318 303 163374 312
rect 87050 232 87106 241
rect 87050 167 87106 176
rect 180904 105 180932 3402
rect 186332 2553 186360 5510
rect 188448 5302 188476 5879
rect 189184 5302 189212 6394
rect 188436 5296 188488 5302
rect 188436 5238 188488 5244
rect 189172 5296 189224 5302
rect 189172 5238 189224 5244
rect 189276 5030 189304 7754
rect 190012 6934 190040 9522
rect 190840 9042 190868 9522
rect 190920 9376 190972 9382
rect 190920 9318 190972 9324
rect 190828 9036 190880 9042
rect 190828 8978 190880 8984
rect 190932 8974 190960 9318
rect 190920 8968 190972 8974
rect 191196 8968 191248 8974
rect 190920 8910 190972 8916
rect 191116 8928 191196 8956
rect 190828 8900 190880 8906
rect 190828 8842 190880 8848
rect 190368 8832 190420 8838
rect 190368 8774 190420 8780
rect 190380 8498 190408 8774
rect 190368 8492 190420 8498
rect 190368 8434 190420 8440
rect 190000 6928 190052 6934
rect 190000 6870 190052 6876
rect 189356 6792 189408 6798
rect 189356 6734 189408 6740
rect 189368 6458 189396 6734
rect 189356 6452 189408 6458
rect 189356 6394 189408 6400
rect 189264 5024 189316 5030
rect 189264 4966 189316 4972
rect 190000 5024 190052 5030
rect 190000 4966 190052 4972
rect 190012 4214 190040 4966
rect 190000 4208 190052 4214
rect 190000 4150 190052 4156
rect 190366 2816 190422 2825
rect 190422 2774 190500 2802
rect 190366 2751 190422 2760
rect 190472 2650 190500 2774
rect 190460 2644 190512 2650
rect 190460 2586 190512 2592
rect 186318 2544 186374 2553
rect 186318 2479 186374 2488
rect 186964 2440 187016 2446
rect 186964 2382 187016 2388
rect 189724 2440 189776 2446
rect 189724 2382 189776 2388
rect 190368 2440 190420 2446
rect 190840 2417 190868 8842
rect 191116 8838 191144 8928
rect 191196 8910 191248 8916
rect 191104 8832 191156 8838
rect 191104 8774 191156 8780
rect 190920 4140 190972 4146
rect 190920 4082 190972 4088
rect 190368 2382 190420 2388
rect 190826 2408 190882 2417
rect 183560 2304 183612 2310
rect 183560 2246 183612 2252
rect 185030 2272 185086 2281
rect 183572 1970 183600 2246
rect 185030 2207 185086 2216
rect 185044 1970 185072 2207
rect 181904 1964 181956 1970
rect 181904 1906 181956 1912
rect 183560 1964 183612 1970
rect 183560 1906 183612 1912
rect 185032 1964 185084 1970
rect 185032 1906 185084 1912
rect 181916 1329 181944 1906
rect 183284 1896 183336 1902
rect 181994 1864 182050 1873
rect 183284 1838 183336 1844
rect 184756 1896 184808 1902
rect 184756 1838 184808 1844
rect 186320 1896 186372 1902
rect 186320 1838 186372 1844
rect 181994 1799 182050 1808
rect 182008 1766 182036 1799
rect 181996 1760 182048 1766
rect 181996 1702 182048 1708
rect 182548 1352 182600 1358
rect 181902 1320 181958 1329
rect 181812 1284 181864 1290
rect 182548 1294 182600 1300
rect 182824 1352 182876 1358
rect 182824 1294 182876 1300
rect 181902 1255 181958 1264
rect 181812 1226 181864 1232
rect 181824 921 181852 1226
rect 181904 1216 181956 1222
rect 181902 1184 181904 1193
rect 181956 1184 181958 1193
rect 181902 1119 181958 1128
rect 182560 921 182588 1294
rect 182836 950 182864 1294
rect 183296 1057 183324 1838
rect 184296 1352 184348 1358
rect 184296 1294 184348 1300
rect 184572 1352 184624 1358
rect 184572 1294 184624 1300
rect 183282 1048 183338 1057
rect 183282 983 183338 992
rect 182824 944 182876 950
rect 181810 912 181866 921
rect 181810 847 181866 856
rect 182546 912 182602 921
rect 184308 921 184336 1294
rect 184584 1193 184612 1294
rect 184570 1184 184626 1193
rect 184570 1119 184626 1128
rect 184768 1057 184796 1838
rect 186332 1465 186360 1838
rect 186318 1456 186374 1465
rect 186318 1391 186374 1400
rect 185584 1352 185636 1358
rect 186976 1329 187004 2382
rect 189736 1970 189764 2382
rect 190380 2106 190408 2382
rect 190826 2343 190882 2352
rect 190368 2100 190420 2106
rect 190368 2042 190420 2048
rect 190840 1970 190868 2343
rect 190932 1970 190960 4082
rect 189724 1964 189776 1970
rect 189724 1906 189776 1912
rect 190828 1964 190880 1970
rect 190828 1906 190880 1912
rect 190920 1964 190972 1970
rect 190920 1906 190972 1912
rect 188160 1896 188212 1902
rect 188160 1838 188212 1844
rect 189448 1896 189500 1902
rect 189448 1838 189500 1844
rect 187148 1352 187200 1358
rect 185584 1294 185636 1300
rect 186962 1320 187018 1329
rect 184754 1048 184810 1057
rect 184754 983 184810 992
rect 185596 921 185624 1294
rect 187148 1294 187200 1300
rect 186962 1255 187018 1264
rect 182824 886 182876 892
rect 184294 912 184350 921
rect 182546 847 182602 856
rect 184294 847 184350 856
rect 185582 912 185638 921
rect 185582 847 185638 856
rect 187160 542 187188 1294
rect 188172 1057 188200 1838
rect 188528 1352 188580 1358
rect 188528 1294 188580 1300
rect 188158 1048 188214 1057
rect 188158 983 188214 992
rect 188540 921 188568 1294
rect 189460 1057 189488 1838
rect 190932 1426 190960 1906
rect 191116 1601 191144 8774
rect 191300 8634 191328 10367
rect 191378 10296 191434 10305
rect 191378 10231 191434 10240
rect 191392 8634 191420 10231
rect 192392 9580 192444 9586
rect 192392 9522 192444 9528
rect 192404 9178 192432 9522
rect 192392 9172 192444 9178
rect 192392 9114 192444 9120
rect 192496 8974 192524 10474
rect 194230 10432 194286 10441
rect 194230 10367 194286 10376
rect 193220 10328 193272 10334
rect 192574 10296 192630 10305
rect 192574 10231 192630 10240
rect 192850 10296 192906 10305
rect 193220 10270 193272 10276
rect 192850 10231 192906 10240
rect 192588 9722 192616 10231
rect 192864 9722 192892 10231
rect 192576 9716 192628 9722
rect 192576 9658 192628 9664
rect 192852 9716 192904 9722
rect 192852 9658 192904 9664
rect 192484 8968 192536 8974
rect 192484 8910 192536 8916
rect 191932 8832 191984 8838
rect 191932 8774 191984 8780
rect 192024 8832 192076 8838
rect 192024 8774 192076 8780
rect 191288 8628 191340 8634
rect 191288 8570 191340 8576
rect 191380 8628 191432 8634
rect 191380 8570 191432 8576
rect 191944 8498 191972 8774
rect 192036 8498 192064 8774
rect 191932 8492 191984 8498
rect 191932 8434 191984 8440
rect 192024 8492 192076 8498
rect 192024 8434 192076 8440
rect 192496 6914 192524 8910
rect 193232 8498 193260 10270
rect 193588 9580 193640 9586
rect 193588 9522 193640 9528
rect 193310 9072 193366 9081
rect 193310 9007 193366 9016
rect 193324 8974 193352 9007
rect 193312 8968 193364 8974
rect 193312 8910 193364 8916
rect 193220 8492 193272 8498
rect 193220 8434 193272 8440
rect 192312 6886 192524 6914
rect 191746 2816 191802 2825
rect 191802 2774 191880 2802
rect 191746 2751 191802 2760
rect 191852 2650 191880 2774
rect 191840 2644 191892 2650
rect 191840 2586 191892 2592
rect 191380 2440 191432 2446
rect 191380 2382 191432 2388
rect 191288 2304 191340 2310
rect 191288 2246 191340 2252
rect 191102 1592 191158 1601
rect 191102 1527 191158 1536
rect 190920 1420 190972 1426
rect 190920 1362 190972 1368
rect 191116 1358 191144 1527
rect 189724 1352 189776 1358
rect 189724 1294 189776 1300
rect 191104 1352 191156 1358
rect 191104 1294 191156 1300
rect 189446 1048 189502 1057
rect 189446 983 189502 992
rect 188526 912 188582 921
rect 189736 882 189764 1294
rect 191300 1193 191328 2246
rect 191392 1494 191420 2382
rect 192312 2038 192340 6886
rect 192392 2440 192444 2446
rect 192392 2382 192444 2388
rect 192404 2106 192432 2382
rect 192392 2100 192444 2106
rect 192392 2042 192444 2048
rect 192300 2032 192352 2038
rect 192300 1974 192352 1980
rect 193232 1970 193260 8434
rect 193324 2038 193352 8910
rect 193496 8900 193548 8906
rect 193496 8842 193548 8848
rect 193508 8498 193536 8842
rect 193600 8634 193628 9522
rect 194048 8832 194100 8838
rect 194048 8774 194100 8780
rect 193588 8628 193640 8634
rect 193588 8570 193640 8576
rect 194060 8498 194088 8774
rect 194244 8634 194272 10367
rect 194322 10296 194378 10305
rect 194322 10231 194378 10240
rect 195610 10296 195666 10305
rect 195610 10231 195666 10240
rect 195794 10296 195850 10305
rect 195794 10231 195850 10240
rect 196530 10296 196586 10305
rect 196530 10231 196586 10240
rect 194336 9722 194364 10231
rect 194324 9716 194376 9722
rect 194324 9658 194376 9664
rect 194416 9512 194468 9518
rect 194416 9454 194468 9460
rect 194600 9512 194652 9518
rect 194600 9454 194652 9460
rect 194232 8628 194284 8634
rect 194232 8570 194284 8576
rect 193496 8492 193548 8498
rect 193496 8434 193548 8440
rect 194048 8492 194100 8498
rect 194048 8434 194100 8440
rect 194428 7993 194456 9454
rect 194612 8974 194640 9454
rect 195520 9376 195572 9382
rect 195520 9318 195572 9324
rect 195532 8974 195560 9318
rect 194600 8968 194652 8974
rect 194600 8910 194652 8916
rect 195520 8968 195572 8974
rect 195520 8910 195572 8916
rect 194414 7984 194470 7993
rect 194414 7919 194470 7928
rect 193312 2032 193364 2038
rect 193312 1974 193364 1980
rect 194612 1970 194640 8910
rect 195532 6914 195560 8910
rect 195624 8634 195652 10231
rect 195808 9722 195836 10231
rect 196544 9722 196572 10231
rect 195796 9716 195848 9722
rect 195796 9658 195848 9664
rect 196532 9716 196584 9722
rect 196532 9658 196584 9664
rect 195796 9580 195848 9586
rect 195796 9522 195848 9528
rect 196624 9580 196676 9586
rect 196624 9522 196676 9528
rect 195808 9178 195836 9522
rect 195796 9172 195848 9178
rect 195796 9114 195848 9120
rect 196256 8968 196308 8974
rect 196256 8910 196308 8916
rect 196532 8968 196584 8974
rect 196532 8910 196584 8916
rect 195612 8628 195664 8634
rect 195612 8570 195664 8576
rect 195440 6886 195560 6914
rect 196268 8378 196296 8910
rect 196348 8832 196400 8838
rect 196348 8774 196400 8780
rect 196360 8498 196388 8774
rect 196544 8566 196572 8910
rect 196636 8634 196664 9522
rect 196624 8628 196676 8634
rect 196624 8570 196676 8576
rect 196532 8560 196584 8566
rect 196532 8502 196584 8508
rect 196348 8492 196400 8498
rect 196348 8434 196400 8440
rect 196728 8430 196756 10542
rect 208306 10503 208362 10512
rect 199474 10432 199530 10441
rect 199474 10367 199530 10376
rect 200946 10432 201002 10441
rect 200946 10367 201002 10376
rect 202602 10432 202658 10441
rect 202602 10367 202658 10376
rect 202788 10396 202840 10402
rect 197266 10296 197322 10305
rect 197266 10231 197322 10240
rect 198002 10296 198058 10305
rect 198002 10231 198058 10240
rect 197280 9450 197308 10231
rect 198016 9722 198044 10231
rect 198648 10124 198700 10130
rect 198648 10066 198700 10072
rect 198004 9716 198056 9722
rect 198004 9658 198056 9664
rect 197544 9580 197596 9586
rect 197544 9522 197596 9528
rect 197912 9580 197964 9586
rect 197912 9522 197964 9528
rect 197268 9444 197320 9450
rect 197268 9386 197320 9392
rect 197176 9104 197228 9110
rect 197176 9046 197228 9052
rect 196532 8424 196584 8430
rect 196268 8362 196388 8378
rect 196532 8366 196584 8372
rect 196716 8424 196768 8430
rect 196716 8366 196768 8372
rect 196268 8356 196400 8362
rect 196268 8350 196348 8356
rect 194692 2304 194744 2310
rect 194692 2246 194744 2252
rect 193220 1964 193272 1970
rect 193220 1906 193272 1912
rect 194600 1964 194652 1970
rect 194600 1906 194652 1912
rect 193220 1760 193272 1766
rect 193220 1702 193272 1708
rect 193312 1760 193364 1766
rect 193312 1702 193364 1708
rect 194600 1760 194652 1766
rect 194600 1702 194652 1708
rect 191380 1488 191432 1494
rect 191380 1430 191432 1436
rect 193232 1358 193260 1702
rect 193324 1358 193352 1702
rect 194612 1358 194640 1702
rect 194704 1465 194732 2246
rect 195440 1970 195468 6886
rect 196268 2774 196296 8350
rect 196348 8298 196400 8304
rect 196544 2774 196572 8366
rect 197188 7857 197216 9046
rect 197360 8968 197412 8974
rect 197360 8910 197412 8916
rect 197372 8498 197400 8910
rect 197556 8634 197584 9522
rect 197924 9178 197952 9522
rect 198188 9444 198240 9450
rect 198188 9386 198240 9392
rect 197912 9172 197964 9178
rect 197912 9114 197964 9120
rect 198096 9104 198148 9110
rect 198200 9081 198228 9386
rect 198096 9046 198148 9052
rect 198186 9072 198242 9081
rect 198004 8968 198056 8974
rect 198004 8910 198056 8916
rect 197544 8628 197596 8634
rect 197544 8570 197596 8576
rect 197360 8492 197412 8498
rect 197360 8434 197412 8440
rect 197268 8424 197320 8430
rect 197268 8366 197320 8372
rect 197174 7848 197230 7857
rect 197174 7783 197230 7792
rect 197280 2774 197308 8366
rect 196176 2746 196296 2774
rect 196452 2746 196572 2774
rect 197188 2746 197308 2774
rect 195704 2440 195756 2446
rect 195704 2382 195756 2388
rect 195716 2106 195744 2382
rect 195980 2304 196032 2310
rect 195980 2246 196032 2252
rect 195704 2100 195756 2106
rect 195704 2042 195756 2048
rect 195428 1964 195480 1970
rect 195428 1906 195480 1912
rect 195992 1465 196020 2246
rect 196176 1970 196204 2746
rect 196256 2440 196308 2446
rect 196256 2382 196308 2388
rect 196268 2106 196296 2382
rect 196256 2100 196308 2106
rect 196256 2042 196308 2048
rect 196452 1970 196480 2746
rect 197188 2446 197216 2746
rect 197176 2440 197228 2446
rect 197176 2382 197228 2388
rect 197268 2440 197320 2446
rect 197268 2382 197320 2388
rect 197280 1970 197308 2382
rect 197452 2304 197504 2310
rect 197452 2246 197504 2252
rect 196164 1964 196216 1970
rect 196164 1906 196216 1912
rect 196440 1964 196492 1970
rect 196440 1906 196492 1912
rect 197268 1964 197320 1970
rect 197268 1906 197320 1912
rect 196532 1760 196584 1766
rect 196532 1702 196584 1708
rect 194690 1456 194746 1465
rect 194690 1391 194746 1400
rect 195978 1456 196034 1465
rect 195978 1391 196034 1400
rect 196544 1358 196572 1702
rect 197464 1358 197492 2246
rect 198016 1970 198044 8910
rect 198108 8634 198136 9046
rect 198186 9007 198242 9016
rect 198660 8974 198688 10066
rect 198832 9580 198884 9586
rect 198832 9522 198884 9528
rect 198648 8968 198700 8974
rect 198648 8910 198700 8916
rect 198844 8634 198872 9522
rect 199292 8832 199344 8838
rect 199292 8774 199344 8780
rect 198096 8628 198148 8634
rect 198096 8570 198148 8576
rect 198832 8628 198884 8634
rect 198832 8570 198884 8576
rect 198108 8430 198136 8570
rect 199304 8498 199332 8774
rect 199488 8634 199516 10367
rect 200026 10296 200082 10305
rect 200026 10231 200082 10240
rect 200854 10296 200910 10305
rect 200854 10231 200910 10240
rect 199660 9920 199712 9926
rect 199660 9862 199712 9868
rect 199672 8974 199700 9862
rect 200040 9722 200068 10231
rect 200028 9716 200080 9722
rect 200028 9658 200080 9664
rect 200120 9716 200172 9722
rect 200120 9658 200172 9664
rect 199844 9580 199896 9586
rect 199844 9522 199896 9528
rect 199856 9178 199884 9522
rect 199844 9172 199896 9178
rect 199844 9114 199896 9120
rect 200132 9110 200160 9658
rect 200672 9376 200724 9382
rect 200672 9318 200724 9324
rect 200120 9104 200172 9110
rect 200120 9046 200172 9052
rect 200684 9042 200712 9318
rect 200672 9036 200724 9042
rect 200672 8978 200724 8984
rect 199660 8968 199712 8974
rect 199660 8910 199712 8916
rect 200488 8968 200540 8974
rect 200488 8910 200540 8916
rect 199476 8628 199528 8634
rect 199476 8570 199528 8576
rect 199292 8492 199344 8498
rect 199292 8434 199344 8440
rect 198096 8424 198148 8430
rect 198096 8366 198148 8372
rect 198832 8424 198884 8430
rect 198832 8366 198884 8372
rect 198844 6662 198872 8366
rect 198832 6656 198884 6662
rect 198832 6598 198884 6604
rect 198556 2304 198608 2310
rect 198556 2246 198608 2252
rect 198004 1964 198056 1970
rect 198004 1906 198056 1912
rect 197912 1760 197964 1766
rect 197912 1702 197964 1708
rect 197924 1358 197952 1702
rect 193220 1352 193272 1358
rect 193220 1294 193272 1300
rect 193312 1352 193364 1358
rect 193312 1294 193364 1300
rect 194600 1352 194652 1358
rect 194600 1294 194652 1300
rect 196532 1352 196584 1358
rect 196532 1294 196584 1300
rect 197452 1352 197504 1358
rect 197452 1294 197504 1300
rect 197912 1352 197964 1358
rect 197912 1294 197964 1300
rect 197268 1284 197320 1290
rect 197268 1226 197320 1232
rect 192668 1216 192720 1222
rect 191286 1184 191342 1193
rect 192668 1158 192720 1164
rect 192944 1216 192996 1222
rect 192944 1158 192996 1164
rect 193680 1216 193732 1222
rect 193680 1158 193732 1164
rect 195796 1216 195848 1222
rect 195796 1158 195848 1164
rect 196624 1216 196676 1222
rect 196624 1158 196676 1164
rect 191286 1119 191342 1128
rect 192680 921 192708 1158
rect 192956 921 192984 1158
rect 193692 921 193720 1158
rect 195808 921 195836 1158
rect 196636 921 196664 1158
rect 197280 921 197308 1226
rect 198568 1193 198596 2246
rect 198844 1970 198872 6598
rect 199200 2440 199252 2446
rect 199200 2382 199252 2388
rect 199212 2106 199240 2382
rect 199200 2100 199252 2106
rect 199200 2042 199252 2048
rect 199672 1970 199700 8910
rect 199936 2304 199988 2310
rect 199936 2246 199988 2252
rect 198832 1964 198884 1970
rect 198832 1906 198884 1912
rect 199660 1964 199712 1970
rect 199660 1906 199712 1912
rect 199752 1760 199804 1766
rect 199752 1702 199804 1708
rect 199764 1358 199792 1702
rect 199752 1352 199804 1358
rect 199948 1329 199976 2246
rect 200500 1970 200528 8910
rect 200868 8634 200896 10231
rect 200960 8634 200988 10367
rect 202510 10296 202566 10305
rect 202510 10231 202566 10240
rect 202524 9722 202552 10231
rect 202616 9722 202644 10367
rect 202788 10338 202840 10344
rect 202512 9716 202564 9722
rect 202512 9658 202564 9664
rect 202604 9716 202656 9722
rect 202604 9658 202656 9664
rect 202696 9580 202748 9586
rect 202696 9522 202748 9528
rect 202052 9104 202104 9110
rect 202052 9046 202104 9052
rect 202064 8974 202092 9046
rect 201132 8968 201184 8974
rect 201132 8910 201184 8916
rect 202052 8968 202104 8974
rect 202052 8910 202104 8916
rect 202604 8968 202656 8974
rect 202604 8910 202656 8916
rect 201040 8832 201092 8838
rect 201040 8774 201092 8780
rect 200856 8628 200908 8634
rect 200856 8570 200908 8576
rect 200948 8628 201000 8634
rect 200948 8570 201000 8576
rect 201052 8498 201080 8774
rect 201040 8492 201092 8498
rect 201040 8434 201092 8440
rect 201144 8362 201172 8910
rect 201132 8356 201184 8362
rect 201132 8298 201184 8304
rect 200764 6316 200816 6322
rect 200764 6258 200816 6264
rect 200776 5846 200804 6258
rect 200764 5840 200816 5846
rect 200764 5782 200816 5788
rect 200856 2440 200908 2446
rect 200856 2382 200908 2388
rect 200868 2106 200896 2382
rect 200856 2100 200908 2106
rect 200856 2042 200908 2048
rect 201144 1970 201172 8298
rect 201224 2440 201276 2446
rect 201224 2382 201276 2388
rect 201316 2440 201368 2446
rect 201316 2382 201368 2388
rect 200488 1964 200540 1970
rect 200488 1906 200540 1912
rect 201132 1964 201184 1970
rect 201132 1906 201184 1912
rect 199752 1294 199804 1300
rect 199934 1320 199990 1329
rect 199934 1255 199990 1264
rect 201236 1222 201264 2382
rect 201328 2106 201356 2382
rect 201408 2304 201460 2310
rect 201408 2246 201460 2252
rect 201316 2100 201368 2106
rect 201316 2042 201368 2048
rect 201328 1358 201356 2042
rect 201316 1352 201368 1358
rect 201316 1294 201368 1300
rect 199936 1216 199988 1222
rect 198554 1184 198610 1193
rect 199936 1158 199988 1164
rect 200672 1216 200724 1222
rect 200672 1158 200724 1164
rect 201224 1216 201276 1222
rect 201420 1193 201448 2246
rect 201684 1760 201736 1766
rect 201684 1702 201736 1708
rect 201696 1290 201724 1702
rect 202064 1426 202092 8910
rect 202512 8900 202564 8906
rect 202512 8842 202564 8848
rect 202420 8832 202472 8838
rect 202420 8774 202472 8780
rect 202432 8498 202460 8774
rect 202524 8498 202552 8842
rect 202616 8838 202644 8910
rect 202604 8832 202656 8838
rect 202604 8774 202656 8780
rect 202420 8492 202472 8498
rect 202420 8434 202472 8440
rect 202512 8492 202564 8498
rect 202512 8434 202564 8440
rect 202236 8424 202288 8430
rect 202236 8366 202288 8372
rect 202248 1970 202276 8366
rect 202328 2984 202380 2990
rect 202328 2926 202380 2932
rect 202236 1964 202288 1970
rect 202236 1906 202288 1912
rect 202340 1426 202368 2926
rect 202616 2514 202644 8774
rect 202708 8634 202736 9522
rect 202696 8628 202748 8634
rect 202696 8570 202748 8576
rect 202800 8430 202828 10338
rect 204074 10296 204130 10305
rect 204074 10231 204130 10240
rect 203740 9820 204048 9829
rect 203740 9818 203746 9820
rect 203802 9818 203826 9820
rect 203882 9818 203906 9820
rect 203962 9818 203986 9820
rect 204042 9818 204048 9820
rect 203802 9766 203804 9818
rect 203984 9766 203986 9818
rect 203740 9764 203746 9766
rect 203802 9764 203826 9766
rect 203882 9764 203906 9766
rect 203962 9764 203986 9766
rect 204042 9764 204048 9766
rect 203740 9755 204048 9764
rect 203432 9580 203484 9586
rect 203432 9522 203484 9528
rect 203444 8974 203472 9522
rect 204088 9178 204116 10231
rect 206558 10160 206614 10169
rect 206558 10095 206614 10104
rect 207662 10160 207718 10169
rect 207662 10095 207718 10104
rect 205822 9616 205878 9625
rect 206572 9586 206600 10095
rect 207676 9586 207704 10095
rect 208320 9586 208348 10503
rect 210882 10432 210938 10441
rect 210882 10367 210938 10376
rect 211710 10432 211766 10441
rect 211710 10367 211766 10376
rect 208400 10260 208452 10266
rect 208400 10202 208452 10208
rect 205822 9551 205824 9560
rect 205876 9551 205878 9560
rect 206560 9580 206612 9586
rect 205824 9522 205876 9528
rect 206560 9522 206612 9528
rect 207664 9580 207716 9586
rect 207664 9522 207716 9528
rect 208308 9580 208360 9586
rect 208308 9522 208360 9528
rect 207388 9376 207440 9382
rect 207388 9318 207440 9324
rect 208124 9376 208176 9382
rect 208124 9318 208176 9324
rect 204076 9172 204128 9178
rect 204076 9114 204128 9120
rect 203616 9104 203668 9110
rect 203616 9046 203668 9052
rect 203432 8968 203484 8974
rect 203432 8910 203484 8916
rect 203524 8968 203576 8974
rect 203524 8910 203576 8916
rect 203536 8634 203564 8910
rect 203628 8838 203656 9046
rect 203616 8832 203668 8838
rect 203616 8774 203668 8780
rect 203740 8732 204048 8741
rect 203740 8730 203746 8732
rect 203802 8730 203826 8732
rect 203882 8730 203906 8732
rect 203962 8730 203986 8732
rect 204042 8730 204048 8732
rect 203802 8678 203804 8730
rect 203984 8678 203986 8730
rect 203740 8676 203746 8678
rect 203802 8676 203826 8678
rect 203882 8676 203906 8678
rect 203962 8676 203986 8678
rect 204042 8676 204048 8678
rect 203740 8667 204048 8676
rect 203524 8628 203576 8634
rect 203524 8570 203576 8576
rect 202788 8424 202840 8430
rect 202788 8366 202840 8372
rect 203156 8424 203208 8430
rect 203156 8366 203208 8372
rect 203168 7954 203196 8366
rect 203156 7948 203208 7954
rect 203156 7890 203208 7896
rect 203740 7644 204048 7653
rect 203740 7642 203746 7644
rect 203802 7642 203826 7644
rect 203882 7642 203906 7644
rect 203962 7642 203986 7644
rect 204042 7642 204048 7644
rect 203802 7590 203804 7642
rect 203984 7590 203986 7642
rect 203740 7588 203746 7590
rect 203802 7588 203826 7590
rect 203882 7588 203906 7590
rect 203962 7588 203986 7590
rect 204042 7588 204048 7590
rect 203740 7579 204048 7588
rect 206928 7200 206980 7206
rect 206928 7142 206980 7148
rect 203740 6556 204048 6565
rect 203740 6554 203746 6556
rect 203802 6554 203826 6556
rect 203882 6554 203906 6556
rect 203962 6554 203986 6556
rect 204042 6554 204048 6556
rect 203802 6502 203804 6554
rect 203984 6502 203986 6554
rect 203740 6500 203746 6502
rect 203802 6500 203826 6502
rect 203882 6500 203906 6502
rect 203962 6500 203986 6502
rect 204042 6500 204048 6502
rect 203740 6491 204048 6500
rect 206940 6118 206968 7142
rect 206928 6112 206980 6118
rect 206928 6054 206980 6060
rect 203740 5468 204048 5477
rect 203740 5466 203746 5468
rect 203802 5466 203826 5468
rect 203882 5466 203906 5468
rect 203962 5466 203986 5468
rect 204042 5466 204048 5468
rect 203802 5414 203804 5466
rect 203984 5414 203986 5466
rect 203740 5412 203746 5414
rect 203802 5412 203826 5414
rect 203882 5412 203906 5414
rect 203962 5412 203986 5414
rect 204042 5412 204048 5414
rect 203740 5403 204048 5412
rect 204258 4992 204314 5001
rect 204258 4927 204314 4936
rect 203740 4380 204048 4389
rect 203740 4378 203746 4380
rect 203802 4378 203826 4380
rect 203882 4378 203906 4380
rect 203962 4378 203986 4380
rect 204042 4378 204048 4380
rect 203802 4326 203804 4378
rect 203984 4326 203986 4378
rect 203740 4324 203746 4326
rect 203802 4324 203826 4326
rect 203882 4324 203906 4326
rect 203962 4324 203986 4326
rect 204042 4324 204048 4326
rect 203740 4315 204048 4324
rect 204272 3534 204300 4927
rect 207202 3768 207258 3777
rect 207202 3703 207258 3712
rect 207216 3602 207244 3703
rect 205088 3596 205140 3602
rect 205088 3538 205140 3544
rect 207204 3596 207256 3602
rect 207204 3538 207256 3544
rect 204260 3528 204312 3534
rect 204260 3470 204312 3476
rect 204904 3528 204956 3534
rect 204904 3470 204956 3476
rect 203740 3292 204048 3301
rect 203740 3290 203746 3292
rect 203802 3290 203826 3292
rect 203882 3290 203906 3292
rect 203962 3290 203986 3292
rect 204042 3290 204048 3292
rect 203802 3238 203804 3290
rect 203984 3238 203986 3290
rect 203740 3236 203746 3238
rect 203802 3236 203826 3238
rect 203882 3236 203906 3238
rect 203962 3236 203986 3238
rect 204042 3236 204048 3238
rect 203740 3227 204048 3236
rect 204916 3194 204944 3470
rect 205100 3466 205128 3538
rect 205088 3460 205140 3466
rect 205088 3402 205140 3408
rect 207112 3460 207164 3466
rect 207112 3402 207164 3408
rect 204904 3188 204956 3194
rect 204904 3130 204956 3136
rect 205100 2990 205128 3402
rect 205088 2984 205140 2990
rect 203798 2952 203854 2961
rect 203798 2887 203800 2896
rect 203852 2887 203854 2896
rect 204442 2952 204498 2961
rect 205088 2926 205140 2932
rect 206376 2984 206428 2990
rect 206376 2926 206428 2932
rect 204442 2887 204444 2896
rect 203800 2858 203852 2864
rect 204496 2887 204498 2896
rect 204444 2858 204496 2864
rect 202786 2816 202842 2825
rect 202842 2774 202920 2802
rect 202786 2751 202842 2760
rect 202892 2650 202920 2774
rect 202880 2644 202932 2650
rect 202880 2586 202932 2592
rect 205100 2514 205128 2926
rect 202604 2508 202656 2514
rect 202604 2450 202656 2456
rect 205088 2508 205140 2514
rect 205088 2450 205140 2456
rect 205364 2508 205416 2514
rect 205364 2450 205416 2456
rect 205376 2310 205404 2450
rect 204260 2304 204312 2310
rect 204260 2246 204312 2252
rect 205364 2304 205416 2310
rect 205364 2246 205416 2252
rect 203740 2204 204048 2213
rect 203740 2202 203746 2204
rect 203802 2202 203826 2204
rect 203882 2202 203906 2204
rect 203962 2202 203986 2204
rect 204042 2202 204048 2204
rect 203802 2150 203804 2202
rect 203984 2150 203986 2202
rect 203740 2148 203746 2150
rect 203802 2148 203826 2150
rect 203882 2148 203906 2150
rect 203962 2148 203986 2150
rect 204042 2148 204048 2150
rect 203740 2139 204048 2148
rect 202880 1760 202932 1766
rect 202880 1702 202932 1708
rect 202892 1601 202920 1702
rect 202878 1592 202934 1601
rect 202878 1527 202934 1536
rect 202052 1420 202104 1426
rect 202052 1362 202104 1368
rect 202328 1420 202380 1426
rect 202328 1362 202380 1368
rect 201684 1284 201736 1290
rect 201684 1226 201736 1232
rect 203340 1216 203392 1222
rect 201224 1158 201276 1164
rect 201406 1184 201462 1193
rect 198554 1119 198610 1128
rect 199948 921 199976 1158
rect 200684 921 200712 1158
rect 203340 1158 203392 1164
rect 201406 1119 201462 1128
rect 203352 921 203380 1158
rect 203740 1116 204048 1125
rect 203740 1114 203746 1116
rect 203802 1114 203826 1116
rect 203882 1114 203906 1116
rect 203962 1114 203986 1116
rect 204042 1114 204048 1116
rect 203802 1062 203804 1114
rect 203984 1062 203986 1114
rect 203740 1060 203746 1062
rect 203802 1060 203826 1062
rect 203882 1060 203906 1062
rect 203962 1060 203986 1062
rect 204042 1060 204048 1062
rect 203740 1051 204048 1060
rect 192666 912 192722 921
rect 188526 847 188582 856
rect 189724 876 189776 882
rect 192666 847 192722 856
rect 192942 912 192998 921
rect 192942 847 192998 856
rect 193678 912 193734 921
rect 193678 847 193734 856
rect 195794 912 195850 921
rect 195794 847 195850 856
rect 196622 912 196678 921
rect 196622 847 196678 856
rect 197266 912 197322 921
rect 197266 847 197322 856
rect 199934 912 199990 921
rect 199934 847 199990 856
rect 200670 912 200726 921
rect 200670 847 200726 856
rect 203338 912 203394 921
rect 203338 847 203394 856
rect 189724 818 189776 824
rect 204272 814 204300 2246
rect 205824 1420 205876 1426
rect 205824 1362 205876 1368
rect 205836 921 205864 1362
rect 206388 1222 206416 2926
rect 207124 2310 207152 3402
rect 207400 3058 207428 9318
rect 207756 6248 207808 6254
rect 207756 6190 207808 6196
rect 207768 4078 207796 6190
rect 207480 4072 207532 4078
rect 207480 4014 207532 4020
rect 207756 4072 207808 4078
rect 207756 4014 207808 4020
rect 207492 3738 207520 4014
rect 207664 3936 207716 3942
rect 207664 3878 207716 3884
rect 207480 3732 207532 3738
rect 207480 3674 207532 3680
rect 207676 3602 207704 3878
rect 207664 3596 207716 3602
rect 207664 3538 207716 3544
rect 207768 3466 207796 4014
rect 208032 4004 208084 4010
rect 208032 3946 208084 3952
rect 207756 3460 207808 3466
rect 207756 3402 207808 3408
rect 208044 3210 208072 3946
rect 207952 3182 208072 3210
rect 207952 3126 207980 3182
rect 207940 3120 207992 3126
rect 207940 3062 207992 3068
rect 207204 3052 207256 3058
rect 207204 2994 207256 3000
rect 207388 3052 207440 3058
rect 207388 2994 207440 3000
rect 207020 2304 207072 2310
rect 207020 2246 207072 2252
rect 207112 2304 207164 2310
rect 207112 2246 207164 2252
rect 207032 2106 207060 2246
rect 207020 2100 207072 2106
rect 207020 2042 207072 2048
rect 206560 1352 206612 1358
rect 206560 1294 206612 1300
rect 206376 1216 206428 1222
rect 206376 1158 206428 1164
rect 206572 921 206600 1294
rect 205822 912 205878 921
rect 205822 847 205878 856
rect 206558 912 206614 921
rect 206558 847 206614 856
rect 204260 808 204312 814
rect 204260 750 204312 756
rect 207216 746 207244 2994
rect 208136 2514 208164 9318
rect 208412 8090 208440 10202
rect 208950 10160 209006 10169
rect 208950 10095 209006 10104
rect 209318 10160 209374 10169
rect 209318 10095 209374 10104
rect 210790 10160 210846 10169
rect 210790 10095 210846 10104
rect 208964 9586 208992 10095
rect 209332 9586 209360 10095
rect 209596 9716 209648 9722
rect 209596 9658 209648 9664
rect 208952 9580 209004 9586
rect 208952 9522 209004 9528
rect 209320 9580 209372 9586
rect 209320 9522 209372 9528
rect 208768 9376 208820 9382
rect 208768 9318 208820 9324
rect 208400 8084 208452 8090
rect 208400 8026 208452 8032
rect 208780 6866 208808 9318
rect 208768 6860 208820 6866
rect 208768 6802 208820 6808
rect 208400 6248 208452 6254
rect 208400 6190 208452 6196
rect 208412 5681 208440 6190
rect 208398 5672 208454 5681
rect 208398 5607 208454 5616
rect 209320 4140 209372 4146
rect 209320 4082 209372 4088
rect 209332 3942 209360 4082
rect 209320 3936 209372 3942
rect 209320 3878 209372 3884
rect 208674 3632 208730 3641
rect 208674 3567 208730 3576
rect 208400 3392 208452 3398
rect 208400 3334 208452 3340
rect 208412 2990 208440 3334
rect 208688 3058 208716 3567
rect 208676 3052 208728 3058
rect 208676 2994 208728 3000
rect 209608 2990 209636 9658
rect 210804 9654 210832 10095
rect 210792 9648 210844 9654
rect 210792 9590 210844 9596
rect 210896 9586 210924 10367
rect 210884 9580 210936 9586
rect 210884 9522 210936 9528
rect 210056 9376 210108 9382
rect 210056 9318 210108 9324
rect 211252 9376 211304 9382
rect 211252 9318 211304 9324
rect 210068 9110 210096 9318
rect 210056 9104 210108 9110
rect 210056 9046 210108 9052
rect 211068 8832 211120 8838
rect 211068 8774 211120 8780
rect 211080 8294 211108 8774
rect 211068 8288 211120 8294
rect 211068 8230 211120 8236
rect 210792 6860 210844 6866
rect 210792 6802 210844 6808
rect 209872 6792 209924 6798
rect 209872 6734 209924 6740
rect 209688 4208 209740 4214
rect 209688 4150 209740 4156
rect 209700 3466 209728 4150
rect 209688 3460 209740 3466
rect 209688 3402 209740 3408
rect 208400 2984 208452 2990
rect 208400 2926 208452 2932
rect 208860 2984 208912 2990
rect 208860 2926 208912 2932
rect 209596 2984 209648 2990
rect 209596 2926 209648 2932
rect 208124 2508 208176 2514
rect 208124 2450 208176 2456
rect 207664 1352 207716 1358
rect 207664 1294 207716 1300
rect 208308 1352 208360 1358
rect 208308 1294 208360 1300
rect 207480 1216 207532 1222
rect 207480 1158 207532 1164
rect 207492 1018 207520 1158
rect 207480 1012 207532 1018
rect 207480 954 207532 960
rect 207676 921 207704 1294
rect 208320 921 208348 1294
rect 207662 912 207718 921
rect 207662 847 207718 856
rect 208306 912 208362 921
rect 208306 847 208362 856
rect 207204 740 207256 746
rect 207204 682 207256 688
rect 208872 678 208900 2926
rect 208952 1352 209004 1358
rect 208952 1294 209004 1300
rect 209780 1352 209832 1358
rect 209780 1294 209832 1300
rect 208964 921 208992 1294
rect 209792 921 209820 1294
rect 209884 1222 209912 6734
rect 209964 5636 210016 5642
rect 209964 5578 210016 5584
rect 209976 4078 210004 5578
rect 210056 5024 210108 5030
rect 210056 4966 210108 4972
rect 209964 4072 210016 4078
rect 209964 4014 210016 4020
rect 210068 3670 210096 4966
rect 210700 4684 210752 4690
rect 210700 4626 210752 4632
rect 210056 3664 210108 3670
rect 210608 3664 210660 3670
rect 210056 3606 210108 3612
rect 210344 3612 210608 3618
rect 210344 3606 210660 3612
rect 210344 3590 210648 3606
rect 210712 3602 210740 4626
rect 210700 3596 210752 3602
rect 210344 3466 210372 3590
rect 210700 3538 210752 3544
rect 210332 3460 210384 3466
rect 210332 3402 210384 3408
rect 210148 3392 210200 3398
rect 210148 3334 210200 3340
rect 210160 2582 210188 3334
rect 210240 2984 210292 2990
rect 210240 2926 210292 2932
rect 210148 2576 210200 2582
rect 210148 2518 210200 2524
rect 209964 2440 210016 2446
rect 209964 2382 210016 2388
rect 209976 1290 210004 2382
rect 209964 1284 210016 1290
rect 209964 1226 210016 1232
rect 209872 1216 209924 1222
rect 209872 1158 209924 1164
rect 210252 1018 210280 2926
rect 210804 2854 210832 6802
rect 211160 6792 211212 6798
rect 211160 6734 211212 6740
rect 211172 5953 211200 6734
rect 211158 5944 211214 5953
rect 211158 5879 211214 5888
rect 210884 3936 210936 3942
rect 210884 3878 210936 3884
rect 210792 2848 210844 2854
rect 210896 2825 210924 3878
rect 211264 3602 211292 9318
rect 211724 8974 211752 10367
rect 213458 10160 213514 10169
rect 213458 10095 213514 10104
rect 213918 10160 213974 10169
rect 213918 10095 213974 10104
rect 212552 9722 212764 9738
rect 212540 9716 212776 9722
rect 212592 9710 212724 9716
rect 212540 9658 212592 9664
rect 212724 9658 212776 9664
rect 213472 9586 213500 10095
rect 213932 9586 213960 10095
rect 212540 9580 212592 9586
rect 212540 9522 212592 9528
rect 213460 9580 213512 9586
rect 213460 9522 213512 9528
rect 213920 9580 213972 9586
rect 213920 9522 213972 9528
rect 212172 9104 212224 9110
rect 212172 9046 212224 9052
rect 212356 9104 212408 9110
rect 212356 9046 212408 9052
rect 211712 8968 211764 8974
rect 211712 8910 211764 8916
rect 211344 6792 211396 6798
rect 211344 6734 211396 6740
rect 211436 6792 211488 6798
rect 211436 6734 211488 6740
rect 211252 3596 211304 3602
rect 211252 3538 211304 3544
rect 210974 3224 211030 3233
rect 210974 3159 211030 3168
rect 210988 3058 211016 3159
rect 210976 3052 211028 3058
rect 210976 2994 211028 3000
rect 211068 3052 211120 3058
rect 211068 2994 211120 3000
rect 210792 2790 210844 2796
rect 210882 2816 210938 2825
rect 210804 2582 210832 2790
rect 211080 2774 211108 2994
rect 211252 2984 211304 2990
rect 211252 2926 211304 2932
rect 210882 2751 210938 2760
rect 210988 2746 211108 2774
rect 210792 2576 210844 2582
rect 210422 2544 210478 2553
rect 210792 2518 210844 2524
rect 210422 2479 210478 2488
rect 210436 2281 210464 2479
rect 210422 2272 210478 2281
rect 210422 2207 210478 2216
rect 210884 1352 210936 1358
rect 210884 1294 210936 1300
rect 210332 1216 210384 1222
rect 210332 1158 210384 1164
rect 210344 1018 210372 1158
rect 210896 1057 210924 1294
rect 210882 1048 210938 1057
rect 210240 1012 210292 1018
rect 210240 954 210292 960
rect 210332 1012 210384 1018
rect 210882 983 210938 992
rect 210332 954 210384 960
rect 210988 950 211016 2746
rect 211264 2446 211292 2926
rect 211068 2440 211120 2446
rect 211068 2382 211120 2388
rect 211252 2440 211304 2446
rect 211252 2382 211304 2388
rect 210976 944 211028 950
rect 208950 912 209006 921
rect 208950 847 209006 856
rect 209778 912 209834 921
rect 210976 886 211028 892
rect 209778 847 209834 856
rect 208860 672 208912 678
rect 208860 614 208912 620
rect 211080 542 211108 2382
rect 211160 2100 211212 2106
rect 211160 2042 211212 2048
rect 211172 882 211200 2042
rect 211160 876 211212 882
rect 211160 818 211212 824
rect 187148 536 187200 542
rect 187148 478 187200 484
rect 211068 536 211120 542
rect 211068 478 211120 484
rect 211356 474 211384 6734
rect 211448 2990 211476 6734
rect 212080 6656 212132 6662
rect 212080 6598 212132 6604
rect 212092 6390 212120 6598
rect 212080 6384 212132 6390
rect 212080 6326 212132 6332
rect 211804 4072 211856 4078
rect 211804 4014 211856 4020
rect 211436 2984 211488 2990
rect 211436 2926 211488 2932
rect 211712 1964 211764 1970
rect 211712 1906 211764 1912
rect 211528 1352 211580 1358
rect 211526 1320 211528 1329
rect 211580 1320 211582 1329
rect 211526 1255 211582 1264
rect 211724 1057 211752 1906
rect 211816 1222 211844 4014
rect 212184 3058 212212 9046
rect 212368 8906 212396 9046
rect 212356 8900 212408 8906
rect 212356 8842 212408 8848
rect 212448 8900 212500 8906
rect 212448 8842 212500 8848
rect 212356 8424 212408 8430
rect 212356 8366 212408 8372
rect 212368 7206 212396 8366
rect 212460 7886 212488 8842
rect 212448 7880 212500 7886
rect 212448 7822 212500 7828
rect 212356 7200 212408 7206
rect 212356 7142 212408 7148
rect 212446 6896 212502 6905
rect 212552 6882 212580 9522
rect 212724 9376 212776 9382
rect 212724 9318 212776 9324
rect 213276 9376 213328 9382
rect 213276 9318 213328 9324
rect 213920 9376 213972 9382
rect 213920 9318 213972 9324
rect 212736 6914 212764 9318
rect 212502 6854 212580 6882
rect 212644 6886 212764 6914
rect 212446 6831 212502 6840
rect 212540 5704 212592 5710
rect 212538 5672 212540 5681
rect 212592 5672 212594 5681
rect 212538 5607 212594 5616
rect 212644 4146 212672 6886
rect 213000 6724 213052 6730
rect 213000 6666 213052 6672
rect 213012 5642 213040 6666
rect 213000 5636 213052 5642
rect 213000 5578 213052 5584
rect 213288 4690 213316 9318
rect 213932 8974 213960 9318
rect 213920 8968 213972 8974
rect 213920 8910 213972 8916
rect 214196 7744 214248 7750
rect 214196 7686 214248 7692
rect 214208 7342 214236 7686
rect 214196 7336 214248 7342
rect 214196 7278 214248 7284
rect 213920 7268 213972 7274
rect 213920 7210 213972 7216
rect 213932 6866 213960 7210
rect 213920 6860 213972 6866
rect 213920 6802 213972 6808
rect 214300 6662 214328 10814
rect 233608 10872 233660 10878
rect 229100 10814 229152 10820
rect 231858 10840 231914 10849
rect 227442 10775 227498 10784
rect 225328 10668 225380 10674
rect 225328 10610 225380 10616
rect 226432 10668 226484 10674
rect 226432 10610 226484 10616
rect 218610 10568 218666 10577
rect 218610 10503 218666 10512
rect 224592 10532 224644 10538
rect 215482 10296 215538 10305
rect 215482 10231 215538 10240
rect 218164 10266 218376 10282
rect 218164 10260 218388 10266
rect 218164 10254 218336 10260
rect 215298 10160 215354 10169
rect 215298 10095 215354 10104
rect 214932 9648 214984 9654
rect 214932 9590 214984 9596
rect 214380 9580 214432 9586
rect 214380 9522 214432 9528
rect 214392 9110 214420 9522
rect 214472 9376 214524 9382
rect 214472 9318 214524 9324
rect 214380 9104 214432 9110
rect 214380 9046 214432 9052
rect 214380 8832 214432 8838
rect 214380 8774 214432 8780
rect 214288 6656 214340 6662
rect 214288 6598 214340 6604
rect 214104 6248 214156 6254
rect 214104 6190 214156 6196
rect 214012 5160 214064 5166
rect 214116 5148 214144 6190
rect 214196 5160 214248 5166
rect 214116 5120 214196 5148
rect 214012 5102 214064 5108
rect 214196 5102 214248 5108
rect 214024 4826 214052 5102
rect 213920 4820 213972 4826
rect 213920 4762 213972 4768
rect 214012 4820 214064 4826
rect 214012 4762 214064 4768
rect 213460 4752 213512 4758
rect 213460 4694 213512 4700
rect 213932 4706 213960 4762
rect 214208 4706 214236 5102
rect 213276 4684 213328 4690
rect 213276 4626 213328 4632
rect 212632 4140 212684 4146
rect 212632 4082 212684 4088
rect 213472 4078 213500 4694
rect 213932 4678 214236 4706
rect 213920 4616 213972 4622
rect 213920 4558 213972 4564
rect 213932 4282 213960 4558
rect 214104 4548 214156 4554
rect 214104 4490 214156 4496
rect 213920 4276 213972 4282
rect 213920 4218 213972 4224
rect 213642 4176 213698 4185
rect 213642 4111 213698 4120
rect 214010 4176 214066 4185
rect 214010 4111 214012 4120
rect 213092 4072 213144 4078
rect 212354 4040 212410 4049
rect 213092 4014 213144 4020
rect 213460 4072 213512 4078
rect 213460 4014 213512 4020
rect 212354 3975 212410 3984
rect 212368 3466 212396 3975
rect 213104 3602 213132 4014
rect 213276 3936 213328 3942
rect 213276 3878 213328 3884
rect 213092 3596 213144 3602
rect 213092 3538 213144 3544
rect 212540 3528 212592 3534
rect 212540 3470 212592 3476
rect 212356 3460 212408 3466
rect 212356 3402 212408 3408
rect 212172 3052 212224 3058
rect 212172 2994 212224 3000
rect 212368 2553 212396 3402
rect 212354 2544 212410 2553
rect 212354 2479 212410 2488
rect 212264 1352 212316 1358
rect 212264 1294 212316 1300
rect 211804 1216 211856 1222
rect 211804 1158 211856 1164
rect 211710 1048 211766 1057
rect 211710 983 211766 992
rect 212276 921 212304 1294
rect 212552 1290 212580 3470
rect 212816 2984 212868 2990
rect 212816 2926 212868 2932
rect 212540 1284 212592 1290
rect 212540 1226 212592 1232
rect 212828 1018 212856 2926
rect 213184 2644 213236 2650
rect 213184 2586 213236 2592
rect 213196 2310 213224 2586
rect 213288 2310 213316 3878
rect 213656 3534 213684 4111
rect 214064 4111 214066 4120
rect 214012 4082 214064 4088
rect 213828 4072 213880 4078
rect 213828 4014 213880 4020
rect 213368 3528 213420 3534
rect 213368 3470 213420 3476
rect 213460 3528 213512 3534
rect 213460 3470 213512 3476
rect 213644 3528 213696 3534
rect 213644 3470 213696 3476
rect 213380 3194 213408 3470
rect 213368 3188 213420 3194
rect 213368 3130 213420 3136
rect 213472 2689 213500 3470
rect 213550 3360 213606 3369
rect 213550 3295 213606 3304
rect 213564 3058 213592 3295
rect 213552 3052 213604 3058
rect 213552 2994 213604 3000
rect 213736 3052 213788 3058
rect 213736 2994 213788 3000
rect 213458 2680 213514 2689
rect 213458 2615 213514 2624
rect 213748 2582 213776 2994
rect 213736 2576 213788 2582
rect 213736 2518 213788 2524
rect 213184 2304 213236 2310
rect 213184 2246 213236 2252
rect 213276 2304 213328 2310
rect 213276 2246 213328 2252
rect 213840 1850 213868 4014
rect 214116 3505 214144 4490
rect 214196 4072 214248 4078
rect 214196 4014 214248 4020
rect 214102 3496 214158 3505
rect 214102 3431 214158 3440
rect 213920 3188 213972 3194
rect 213920 3130 213972 3136
rect 213932 2961 213960 3130
rect 213918 2952 213974 2961
rect 213918 2887 213974 2896
rect 214116 2446 214144 3431
rect 214104 2440 214156 2446
rect 214104 2382 214156 2388
rect 213656 1822 213868 1850
rect 213460 1352 213512 1358
rect 213460 1294 213512 1300
rect 212816 1012 212868 1018
rect 212816 954 212868 960
rect 213472 921 213500 1294
rect 212262 912 212318 921
rect 212262 847 212318 856
rect 213458 912 213514 921
rect 213458 847 213514 856
rect 213656 814 213684 1822
rect 213736 1352 213788 1358
rect 213736 1294 213788 1300
rect 213748 921 213776 1294
rect 213828 1216 213880 1222
rect 214208 1204 214236 4014
rect 214392 3602 214420 8774
rect 214484 7410 214512 9318
rect 214564 9104 214616 9110
rect 214564 9046 214616 9052
rect 214576 8294 214604 9046
rect 214564 8288 214616 8294
rect 214564 8230 214616 8236
rect 214656 7880 214708 7886
rect 214656 7822 214708 7828
rect 214472 7404 214524 7410
rect 214472 7346 214524 7352
rect 214562 6352 214618 6361
rect 214562 6287 214618 6296
rect 214576 4865 214604 6287
rect 214668 6254 214696 7822
rect 214838 7712 214894 7721
rect 214838 7647 214894 7656
rect 214852 7274 214880 7647
rect 214840 7268 214892 7274
rect 214840 7210 214892 7216
rect 214656 6248 214708 6254
rect 214656 6190 214708 6196
rect 214656 5704 214708 5710
rect 214654 5672 214656 5681
rect 214708 5672 214710 5681
rect 214654 5607 214710 5616
rect 214668 5574 214696 5607
rect 214656 5568 214708 5574
rect 214656 5510 214708 5516
rect 214562 4856 214618 4865
rect 214562 4791 214618 4800
rect 214564 4616 214616 4622
rect 214564 4558 214616 4564
rect 214470 3768 214526 3777
rect 214470 3703 214526 3712
rect 214380 3596 214432 3602
rect 214380 3538 214432 3544
rect 214484 3194 214512 3703
rect 214472 3188 214524 3194
rect 214472 3130 214524 3136
rect 214380 2984 214432 2990
rect 214380 2926 214432 2932
rect 214392 1222 214420 2926
rect 214472 1352 214524 1358
rect 214472 1294 214524 1300
rect 213880 1176 214236 1204
rect 214380 1216 214432 1222
rect 213828 1158 213880 1164
rect 214380 1158 214432 1164
rect 214484 921 214512 1294
rect 214576 1290 214604 4558
rect 214944 4146 214972 9590
rect 215312 9586 215340 10095
rect 215496 9586 215524 10231
rect 216678 10160 216734 10169
rect 216678 10095 216734 10104
rect 217966 10160 218022 10169
rect 218164 10130 218192 10254
rect 218336 10202 218388 10208
rect 217966 10095 218022 10104
rect 218152 10124 218204 10130
rect 216692 9586 216720 10095
rect 216862 9888 216918 9897
rect 216862 9823 216918 9832
rect 215300 9580 215352 9586
rect 215300 9522 215352 9528
rect 215484 9580 215536 9586
rect 215484 9522 215536 9528
rect 216680 9580 216732 9586
rect 216680 9522 216732 9528
rect 215392 9376 215444 9382
rect 215392 9318 215444 9324
rect 215036 7398 215248 7426
rect 215036 7342 215064 7398
rect 215024 7336 215076 7342
rect 215024 7278 215076 7284
rect 215116 7336 215168 7342
rect 215116 7278 215168 7284
rect 215128 7002 215156 7278
rect 215116 6996 215168 7002
rect 215116 6938 215168 6944
rect 215022 6896 215078 6905
rect 215022 6831 215078 6840
rect 215116 6860 215168 6866
rect 215036 5098 215064 6831
rect 215116 6802 215168 6808
rect 215128 5545 215156 6802
rect 215114 5536 215170 5545
rect 215114 5471 215170 5480
rect 215024 5092 215076 5098
rect 215024 5034 215076 5040
rect 215116 4480 215168 4486
rect 215116 4422 215168 4428
rect 215128 4282 215156 4422
rect 215116 4276 215168 4282
rect 215116 4218 215168 4224
rect 214932 4140 214984 4146
rect 214932 4082 214984 4088
rect 214656 3936 214708 3942
rect 214656 3878 214708 3884
rect 214668 3670 214696 3878
rect 214656 3664 214708 3670
rect 214656 3606 214708 3612
rect 214564 1284 214616 1290
rect 214564 1226 214616 1232
rect 215116 1284 215168 1290
rect 215116 1226 215168 1232
rect 215128 921 215156 1226
rect 215220 1222 215248 7398
rect 215298 7032 215354 7041
rect 215298 6967 215354 6976
rect 215312 6254 215340 6967
rect 215300 6248 215352 6254
rect 215300 6190 215352 6196
rect 215404 5778 215432 9318
rect 216876 8974 216904 9823
rect 217980 9586 218008 10095
rect 218152 10066 218204 10072
rect 218244 10124 218296 10130
rect 218244 10066 218296 10072
rect 217968 9580 218020 9586
rect 217968 9522 218020 9528
rect 218256 9518 218284 10066
rect 218624 9586 218652 10503
rect 224592 10474 224644 10480
rect 221830 10432 221886 10441
rect 221830 10367 221886 10376
rect 220818 10296 220874 10305
rect 220818 10231 220874 10240
rect 219254 10160 219310 10169
rect 219254 10095 219310 10104
rect 220542 10160 220598 10169
rect 220542 10095 220598 10104
rect 219268 9586 219296 10095
rect 220556 9586 220584 10095
rect 220832 9586 220860 10231
rect 221844 9586 221872 10367
rect 222014 10296 222070 10305
rect 222014 10231 222070 10240
rect 223118 10296 223174 10305
rect 223118 10231 223174 10240
rect 218612 9580 218664 9586
rect 218612 9522 218664 9528
rect 219256 9580 219308 9586
rect 219256 9522 219308 9528
rect 220544 9580 220596 9586
rect 220544 9522 220596 9528
rect 220820 9580 220872 9586
rect 220820 9522 220872 9528
rect 221832 9580 221884 9586
rect 221832 9522 221884 9528
rect 218244 9512 218296 9518
rect 218244 9454 218296 9460
rect 219164 9444 219216 9450
rect 219164 9386 219216 9392
rect 217692 9376 217744 9382
rect 217692 9318 217744 9324
rect 217784 9376 217836 9382
rect 217784 9318 217836 9324
rect 215668 8968 215720 8974
rect 215668 8910 215720 8916
rect 216864 8968 216916 8974
rect 216864 8910 216916 8916
rect 215576 7404 215628 7410
rect 215576 7346 215628 7352
rect 215588 7177 215616 7346
rect 215574 7168 215630 7177
rect 215574 7103 215630 7112
rect 215484 6996 215536 7002
rect 215484 6938 215536 6944
rect 215392 5772 215444 5778
rect 215392 5714 215444 5720
rect 215496 5642 215524 6938
rect 215574 6760 215630 6769
rect 215574 6695 215630 6704
rect 215588 6662 215616 6695
rect 215576 6656 215628 6662
rect 215576 6598 215628 6604
rect 215576 5704 215628 5710
rect 215576 5646 215628 5652
rect 215484 5636 215536 5642
rect 215484 5578 215536 5584
rect 215484 4752 215536 4758
rect 215484 4694 215536 4700
rect 215496 4078 215524 4694
rect 215484 4072 215536 4078
rect 215484 4014 215536 4020
rect 215392 3528 215444 3534
rect 215392 3470 215444 3476
rect 215404 2106 215432 3470
rect 215392 2100 215444 2106
rect 215392 2042 215444 2048
rect 215588 1222 215616 5646
rect 215680 2990 215708 8910
rect 216680 8832 216732 8838
rect 216680 8774 216732 8780
rect 216312 7948 216364 7954
rect 216312 7890 216364 7896
rect 215944 6928 215996 6934
rect 215944 6870 215996 6876
rect 215956 5778 215984 6870
rect 216324 6730 216352 7890
rect 216404 7744 216456 7750
rect 216404 7686 216456 7692
rect 216496 7744 216548 7750
rect 216496 7686 216548 7692
rect 216416 7410 216444 7686
rect 216404 7404 216456 7410
rect 216404 7346 216456 7352
rect 216404 7268 216456 7274
rect 216508 7256 216536 7686
rect 216692 7410 216720 8774
rect 216680 7404 216732 7410
rect 216680 7346 216732 7352
rect 216588 7336 216640 7342
rect 216588 7278 216640 7284
rect 216956 7336 217008 7342
rect 216956 7278 217008 7284
rect 216456 7228 216536 7256
rect 216404 7210 216456 7216
rect 216312 6724 216364 6730
rect 216312 6666 216364 6672
rect 216036 5908 216088 5914
rect 216036 5850 216088 5856
rect 215944 5772 215996 5778
rect 215944 5714 215996 5720
rect 215956 5658 215984 5714
rect 215772 5630 215984 5658
rect 215772 3670 215800 5630
rect 216048 5574 216076 5850
rect 216128 5772 216180 5778
rect 216128 5714 216180 5720
rect 215944 5568 215996 5574
rect 215944 5510 215996 5516
rect 216036 5568 216088 5574
rect 216036 5510 216088 5516
rect 215852 5364 215904 5370
rect 215852 5306 215904 5312
rect 215864 4758 215892 5306
rect 215956 5098 215984 5510
rect 215944 5092 215996 5098
rect 215944 5034 215996 5040
rect 215852 4752 215904 4758
rect 216140 4706 216168 5714
rect 216312 5704 216364 5710
rect 216310 5672 216312 5681
rect 216364 5672 216366 5681
rect 216310 5607 216366 5616
rect 215852 4694 215904 4700
rect 216048 4678 216168 4706
rect 216218 4720 216274 4729
rect 216048 4185 216076 4678
rect 216416 4690 216444 7210
rect 216600 6934 216628 7278
rect 216588 6928 216640 6934
rect 216588 6870 216640 6876
rect 216770 6896 216826 6905
rect 216770 6831 216826 6840
rect 216784 6458 216812 6831
rect 216772 6452 216824 6458
rect 216772 6394 216824 6400
rect 216496 5704 216548 5710
rect 216496 5646 216548 5652
rect 216218 4655 216274 4664
rect 216404 4684 216456 4690
rect 216128 4616 216180 4622
rect 216232 4604 216260 4655
rect 216404 4626 216456 4632
rect 216180 4576 216260 4604
rect 216312 4616 216364 4622
rect 216128 4558 216180 4564
rect 216312 4558 216364 4564
rect 216034 4176 216090 4185
rect 215852 4140 215904 4146
rect 216128 4140 216180 4146
rect 216090 4120 216128 4128
rect 216034 4111 216128 4120
rect 216048 4100 216128 4111
rect 215852 4082 215904 4088
rect 216128 4082 216180 4088
rect 215760 3664 215812 3670
rect 215760 3606 215812 3612
rect 215772 2990 215800 3606
rect 215864 3398 215892 4082
rect 216126 3904 216182 3913
rect 216126 3839 216182 3848
rect 216140 3602 216168 3839
rect 216128 3596 216180 3602
rect 216048 3556 216128 3584
rect 215852 3392 215904 3398
rect 215852 3334 215904 3340
rect 215668 2984 215720 2990
rect 215668 2926 215720 2932
rect 215760 2984 215812 2990
rect 215760 2926 215812 2932
rect 215772 2854 215800 2926
rect 215760 2848 215812 2854
rect 215760 2790 215812 2796
rect 215864 2689 215892 3334
rect 216048 3194 216076 3556
rect 216128 3538 216180 3544
rect 216036 3188 216088 3194
rect 216324 3176 216352 4558
rect 216416 3534 216444 4626
rect 216508 4049 216536 5646
rect 216588 5160 216640 5166
rect 216588 5102 216640 5108
rect 216494 4040 216550 4049
rect 216494 3975 216550 3984
rect 216600 3942 216628 5102
rect 216864 4208 216916 4214
rect 216864 4150 216916 4156
rect 216588 3936 216640 3942
rect 216588 3878 216640 3884
rect 216600 3777 216628 3878
rect 216586 3768 216642 3777
rect 216586 3703 216642 3712
rect 216404 3528 216456 3534
rect 216456 3488 216628 3516
rect 216404 3470 216456 3476
rect 216496 3392 216548 3398
rect 216496 3334 216548 3340
rect 216036 3130 216088 3136
rect 216232 3148 216352 3176
rect 215666 2680 215722 2689
rect 215666 2615 215722 2624
rect 215850 2680 215906 2689
rect 215850 2615 215906 2624
rect 215680 2145 215708 2615
rect 216128 2508 216180 2514
rect 216128 2450 216180 2456
rect 215758 2408 215814 2417
rect 215758 2343 215814 2352
rect 215666 2136 215722 2145
rect 215666 2071 215722 2080
rect 215772 1737 215800 2343
rect 216140 1766 216168 2450
rect 216128 1760 216180 1766
rect 215758 1728 215814 1737
rect 216128 1702 216180 1708
rect 215758 1663 215814 1672
rect 215208 1216 215260 1222
rect 215208 1158 215260 1164
rect 215576 1216 215628 1222
rect 215576 1158 215628 1164
rect 213734 912 213790 921
rect 213734 847 213790 856
rect 214470 912 214526 921
rect 214470 847 214526 856
rect 215114 912 215170 921
rect 215114 847 215170 856
rect 213644 808 213696 814
rect 213644 750 213696 756
rect 211344 468 211396 474
rect 211344 410 211396 416
rect 216232 338 216260 3148
rect 216310 3088 216366 3097
rect 216310 3023 216312 3032
rect 216364 3023 216366 3032
rect 216312 2994 216364 3000
rect 216508 2990 216536 3334
rect 216600 3058 216628 3488
rect 216588 3052 216640 3058
rect 216588 2994 216640 3000
rect 216496 2984 216548 2990
rect 216496 2926 216548 2932
rect 216600 2854 216628 2994
rect 216772 2984 216824 2990
rect 216772 2926 216824 2932
rect 216588 2848 216640 2854
rect 216588 2790 216640 2796
rect 216784 2553 216812 2926
rect 216770 2544 216826 2553
rect 216770 2479 216826 2488
rect 216404 2304 216456 2310
rect 216404 2246 216456 2252
rect 216678 2272 216734 2281
rect 216416 1970 216444 2246
rect 216678 2207 216734 2216
rect 216692 2038 216720 2207
rect 216680 2032 216732 2038
rect 216680 1974 216732 1980
rect 216404 1964 216456 1970
rect 216404 1906 216456 1912
rect 216680 1828 216732 1834
rect 216680 1770 216732 1776
rect 216588 1556 216640 1562
rect 216588 1498 216640 1504
rect 216600 474 216628 1498
rect 216692 1465 216720 1770
rect 216678 1456 216734 1465
rect 216678 1391 216734 1400
rect 216680 1352 216732 1358
rect 216680 1294 216732 1300
rect 216692 921 216720 1294
rect 216876 950 216904 4150
rect 216968 2106 216996 7278
rect 217704 6798 217732 9318
rect 217692 6792 217744 6798
rect 217692 6734 217744 6740
rect 217600 6724 217652 6730
rect 217600 6666 217652 6672
rect 217140 6248 217192 6254
rect 217140 6190 217192 6196
rect 217152 5642 217180 6190
rect 217140 5636 217192 5642
rect 217140 5578 217192 5584
rect 217416 4752 217468 4758
rect 217414 4720 217416 4729
rect 217468 4720 217470 4729
rect 217414 4655 217470 4664
rect 217506 3904 217562 3913
rect 217506 3839 217562 3848
rect 217520 3670 217548 3839
rect 217416 3664 217468 3670
rect 217416 3606 217468 3612
rect 217508 3664 217560 3670
rect 217508 3606 217560 3612
rect 217232 3528 217284 3534
rect 217232 3470 217284 3476
rect 217244 3194 217272 3470
rect 217428 3398 217456 3606
rect 217416 3392 217468 3398
rect 217416 3334 217468 3340
rect 217232 3188 217284 3194
rect 217232 3130 217284 3136
rect 217428 2922 217456 3334
rect 217416 2916 217468 2922
rect 217416 2858 217468 2864
rect 217138 2816 217194 2825
rect 217138 2751 217194 2760
rect 217152 2106 217180 2751
rect 216956 2100 217008 2106
rect 216956 2042 217008 2048
rect 217140 2100 217192 2106
rect 217140 2042 217192 2048
rect 217612 1290 217640 6666
rect 217692 6656 217744 6662
rect 217692 6598 217744 6604
rect 217704 4729 217732 6598
rect 217796 6322 217824 9318
rect 217968 8492 218020 8498
rect 217968 8434 218020 8440
rect 217980 8090 218008 8434
rect 217968 8084 218020 8090
rect 217968 8026 218020 8032
rect 218704 7948 218756 7954
rect 218704 7890 218756 7896
rect 217968 7812 218020 7818
rect 217968 7754 218020 7760
rect 217980 7478 218008 7754
rect 218336 7744 218388 7750
rect 218336 7686 218388 7692
rect 218428 7744 218480 7750
rect 218428 7686 218480 7692
rect 217968 7472 218020 7478
rect 217968 7414 218020 7420
rect 218060 7200 218112 7206
rect 218060 7142 218112 7148
rect 218072 6866 218100 7142
rect 218348 6934 218376 7686
rect 218440 7274 218468 7686
rect 218716 7546 218744 7890
rect 218980 7744 219032 7750
rect 218980 7686 219032 7692
rect 218704 7540 218756 7546
rect 218704 7482 218756 7488
rect 218992 7410 219020 7686
rect 218704 7404 218756 7410
rect 218704 7346 218756 7352
rect 218980 7404 219032 7410
rect 218980 7346 219032 7352
rect 218428 7268 218480 7274
rect 218428 7210 218480 7216
rect 218336 6928 218388 6934
rect 218336 6870 218388 6876
rect 218060 6860 218112 6866
rect 218060 6802 218112 6808
rect 217876 6656 217928 6662
rect 217876 6598 217928 6604
rect 217888 6390 217916 6598
rect 218336 6452 218388 6458
rect 218336 6394 218388 6400
rect 217876 6384 217928 6390
rect 217876 6326 217928 6332
rect 217784 6316 217836 6322
rect 217784 6258 217836 6264
rect 218348 6254 218376 6394
rect 217968 6248 218020 6254
rect 217968 6190 218020 6196
rect 218336 6248 218388 6254
rect 218336 6190 218388 6196
rect 217690 4720 217746 4729
rect 217690 4655 217746 4664
rect 217784 2848 217836 2854
rect 217784 2790 217836 2796
rect 217796 1358 217824 2790
rect 217874 2544 217930 2553
rect 217874 2479 217930 2488
rect 217784 1352 217836 1358
rect 217784 1294 217836 1300
rect 217600 1284 217652 1290
rect 217600 1226 217652 1232
rect 217416 1216 217468 1222
rect 217416 1158 217468 1164
rect 216864 944 216916 950
rect 216678 912 216734 921
rect 217428 921 217456 1158
rect 216864 886 216916 892
rect 217414 912 217470 921
rect 216678 847 216734 856
rect 217414 847 217470 856
rect 217324 740 217376 746
rect 217324 682 217376 688
rect 217336 610 217364 682
rect 217324 604 217376 610
rect 217324 546 217376 552
rect 216588 468 216640 474
rect 216588 410 216640 416
rect 217888 406 217916 2479
rect 217980 1018 218008 6190
rect 218060 6180 218112 6186
rect 218060 6122 218112 6128
rect 218072 3126 218100 6122
rect 218440 5386 218468 7210
rect 218716 7177 218744 7346
rect 218518 7168 218574 7177
rect 218518 7103 218574 7112
rect 218702 7168 218758 7177
rect 218702 7103 218758 7112
rect 218164 5370 218468 5386
rect 218152 5364 218468 5370
rect 218204 5358 218468 5364
rect 218152 5306 218204 5312
rect 218152 3936 218204 3942
rect 218152 3878 218204 3884
rect 218060 3120 218112 3126
rect 218060 3062 218112 3068
rect 218164 2990 218192 3878
rect 218152 2984 218204 2990
rect 218152 2926 218204 2932
rect 218060 2440 218112 2446
rect 218060 2382 218112 2388
rect 218072 1902 218100 2382
rect 218152 2304 218204 2310
rect 218152 2246 218204 2252
rect 218060 1896 218112 1902
rect 218060 1838 218112 1844
rect 218164 1358 218192 2246
rect 218152 1352 218204 1358
rect 218152 1294 218204 1300
rect 218060 1284 218112 1290
rect 218060 1226 218112 1232
rect 217968 1012 218020 1018
rect 217968 954 218020 960
rect 218072 950 218100 1226
rect 218532 1193 218560 7103
rect 218888 6792 218940 6798
rect 218886 6760 218888 6769
rect 218940 6760 218942 6769
rect 218886 6695 218942 6704
rect 218992 6338 219020 7346
rect 219072 6792 219124 6798
rect 219072 6734 219124 6740
rect 218900 6310 219020 6338
rect 218796 6248 218848 6254
rect 218796 6190 218848 6196
rect 218704 5024 218756 5030
rect 218704 4966 218756 4972
rect 218716 3194 218744 4966
rect 218808 3777 218836 6190
rect 218900 5778 218928 6310
rect 218980 6248 219032 6254
rect 218978 6216 218980 6225
rect 219032 6216 219034 6225
rect 218978 6151 219034 6160
rect 218888 5772 218940 5778
rect 218888 5714 218940 5720
rect 218888 4480 218940 4486
rect 218888 4422 218940 4428
rect 218794 3768 218850 3777
rect 218794 3703 218850 3712
rect 218900 3602 218928 4422
rect 219084 4282 219112 6734
rect 219176 6254 219204 9386
rect 219348 9376 219400 9382
rect 219348 9318 219400 9324
rect 220360 9376 220412 9382
rect 220360 9318 220412 9324
rect 219360 6866 219388 9318
rect 219624 7744 219676 7750
rect 219624 7686 219676 7692
rect 219636 6905 219664 7686
rect 220372 7410 220400 9318
rect 221924 9036 221976 9042
rect 221924 8978 221976 8984
rect 221936 8838 221964 8978
rect 222028 8974 222056 10231
rect 223132 9586 223160 10231
rect 223302 10160 223358 10169
rect 223302 10095 223358 10104
rect 223316 9586 223344 10095
rect 224316 9716 224368 9722
rect 224316 9658 224368 9664
rect 224328 9586 224356 9658
rect 224604 9586 224632 10474
rect 225340 10334 225368 10610
rect 225420 10532 225472 10538
rect 225420 10474 225472 10480
rect 225328 10328 225380 10334
rect 225328 10270 225380 10276
rect 223120 9580 223172 9586
rect 223120 9522 223172 9528
rect 223304 9580 223356 9586
rect 223304 9522 223356 9528
rect 224316 9580 224368 9586
rect 224316 9522 224368 9528
rect 224592 9580 224644 9586
rect 224592 9522 224644 9528
rect 224776 9580 224828 9586
rect 224776 9522 224828 9528
rect 224408 9512 224460 9518
rect 224788 9489 224816 9522
rect 224408 9454 224460 9460
rect 224774 9480 224830 9489
rect 222108 9444 222160 9450
rect 222108 9386 222160 9392
rect 222200 9444 222252 9450
rect 222200 9386 222252 9392
rect 222016 8968 222068 8974
rect 222016 8910 222068 8916
rect 221832 8832 221884 8838
rect 221832 8774 221884 8780
rect 221924 8832 221976 8838
rect 221924 8774 221976 8780
rect 221844 8498 221872 8774
rect 220912 8492 220964 8498
rect 220912 8434 220964 8440
rect 221832 8492 221884 8498
rect 221832 8434 221884 8440
rect 220634 7848 220690 7857
rect 220634 7783 220690 7792
rect 220360 7404 220412 7410
rect 220360 7346 220412 7352
rect 219992 7268 220044 7274
rect 219992 7210 220044 7216
rect 220544 7268 220596 7274
rect 220544 7210 220596 7216
rect 219716 7200 219768 7206
rect 219714 7168 219716 7177
rect 219768 7168 219770 7177
rect 219714 7103 219770 7112
rect 219622 6896 219678 6905
rect 219348 6860 219400 6866
rect 219622 6831 219678 6840
rect 219348 6802 219400 6808
rect 219900 6792 219952 6798
rect 219900 6734 219952 6740
rect 219912 6458 219940 6734
rect 220004 6497 220032 7210
rect 220556 6866 220584 7210
rect 220648 6905 220676 7783
rect 220728 7336 220780 7342
rect 220728 7278 220780 7284
rect 220818 7304 220874 7313
rect 220634 6896 220690 6905
rect 220544 6860 220596 6866
rect 220634 6831 220690 6840
rect 220544 6802 220596 6808
rect 219990 6488 220046 6497
rect 219900 6452 219952 6458
rect 219990 6423 220046 6432
rect 219900 6394 219952 6400
rect 219164 6248 219216 6254
rect 219164 6190 219216 6196
rect 219912 6186 219940 6394
rect 220360 6248 220412 6254
rect 220360 6190 220412 6196
rect 220544 6248 220596 6254
rect 220544 6190 220596 6196
rect 219900 6180 219952 6186
rect 219900 6122 219952 6128
rect 219164 6112 219216 6118
rect 219164 6054 219216 6060
rect 219440 6112 219492 6118
rect 219440 6054 219492 6060
rect 219072 4276 219124 4282
rect 219072 4218 219124 4224
rect 218888 3596 218940 3602
rect 218888 3538 218940 3544
rect 218704 3188 218756 3194
rect 218704 3130 218756 3136
rect 218716 2774 218744 3130
rect 218900 3126 218928 3538
rect 219176 3534 219204 6054
rect 219256 5636 219308 5642
rect 219256 5578 219308 5584
rect 219268 5409 219296 5578
rect 219254 5400 219310 5409
rect 219254 5335 219310 5344
rect 219452 5250 219480 6054
rect 219268 5234 219480 5250
rect 220176 5296 220228 5302
rect 220176 5238 220228 5244
rect 219256 5228 219480 5234
rect 219308 5222 219480 5228
rect 219256 5170 219308 5176
rect 219714 4856 219770 4865
rect 219714 4791 219716 4800
rect 219768 4791 219770 4800
rect 219716 4762 219768 4768
rect 220188 4554 220216 5238
rect 220176 4548 220228 4554
rect 220176 4490 220228 4496
rect 219164 3528 219216 3534
rect 219164 3470 219216 3476
rect 220188 3466 220216 4490
rect 220176 3460 220228 3466
rect 220176 3402 220228 3408
rect 218888 3120 218940 3126
rect 218888 3062 218940 3068
rect 219072 2984 219124 2990
rect 219072 2926 219124 2932
rect 218624 2746 218744 2774
rect 218624 2514 218652 2746
rect 218612 2508 218664 2514
rect 218612 2450 218664 2456
rect 219084 2446 219112 2926
rect 219440 2848 219492 2854
rect 219440 2790 219492 2796
rect 219072 2440 219124 2446
rect 219072 2382 219124 2388
rect 219452 1970 219480 2790
rect 219808 2304 219860 2310
rect 219808 2246 219860 2252
rect 219440 1964 219492 1970
rect 219440 1906 219492 1912
rect 218980 1284 219032 1290
rect 218980 1226 219032 1232
rect 219440 1284 219492 1290
rect 219440 1226 219492 1232
rect 218518 1184 218574 1193
rect 218518 1119 218574 1128
rect 218992 1057 219020 1226
rect 218978 1048 219034 1057
rect 218978 983 219034 992
rect 218060 944 218112 950
rect 219452 921 219480 1226
rect 219624 1216 219676 1222
rect 219624 1158 219676 1164
rect 219636 1018 219664 1158
rect 219624 1012 219676 1018
rect 219624 954 219676 960
rect 218060 886 218112 892
rect 219438 912 219494 921
rect 219820 882 219848 2246
rect 220082 2000 220138 2009
rect 220082 1935 220084 1944
rect 220136 1935 220138 1944
rect 220084 1906 220136 1912
rect 220372 1222 220400 6190
rect 220556 5137 220584 6190
rect 220636 6112 220688 6118
rect 220636 6054 220688 6060
rect 220542 5128 220598 5137
rect 220542 5063 220598 5072
rect 220648 4690 220676 6054
rect 220636 4684 220688 4690
rect 220636 4626 220688 4632
rect 220740 2496 220768 7278
rect 220818 7239 220874 7248
rect 220832 7002 220860 7239
rect 220924 7177 220952 8434
rect 221096 8016 221148 8022
rect 221096 7958 221148 7964
rect 220910 7168 220966 7177
rect 220910 7103 220966 7112
rect 220820 6996 220872 7002
rect 220820 6938 220872 6944
rect 220912 6928 220964 6934
rect 220964 6888 221044 6916
rect 220912 6870 220964 6876
rect 220912 6656 220964 6662
rect 220912 6598 220964 6604
rect 220648 2468 220768 2496
rect 220648 1562 220676 2468
rect 220728 2372 220780 2378
rect 220728 2314 220780 2320
rect 220740 1970 220768 2314
rect 220728 1964 220780 1970
rect 220728 1906 220780 1912
rect 220820 1964 220872 1970
rect 220820 1906 220872 1912
rect 220636 1556 220688 1562
rect 220636 1498 220688 1504
rect 220832 1465 220860 1906
rect 220818 1456 220874 1465
rect 220818 1391 220874 1400
rect 220728 1284 220780 1290
rect 220728 1226 220780 1232
rect 220360 1216 220412 1222
rect 220360 1158 220412 1164
rect 220084 944 220136 950
rect 220268 944 220320 950
rect 220136 892 220268 898
rect 220084 886 220320 892
rect 219438 847 219494 856
rect 219808 876 219860 882
rect 220096 870 220308 886
rect 219808 818 219860 824
rect 218888 740 218940 746
rect 218888 682 218940 688
rect 217876 400 217928 406
rect 218900 377 218928 682
rect 220740 406 220768 1226
rect 220924 1222 220952 6598
rect 221016 5914 221044 6888
rect 221108 6866 221136 7958
rect 221464 7540 221516 7546
rect 221464 7482 221516 7488
rect 221476 7410 221504 7482
rect 221464 7404 221516 7410
rect 221464 7346 221516 7352
rect 221556 7404 221608 7410
rect 221556 7346 221608 7352
rect 221740 7404 221792 7410
rect 221740 7346 221792 7352
rect 221370 7304 221426 7313
rect 221370 7239 221426 7248
rect 221096 6860 221148 6866
rect 221096 6802 221148 6808
rect 221280 6792 221332 6798
rect 221384 6780 221412 7239
rect 221332 6752 221412 6780
rect 221280 6734 221332 6740
rect 221188 6452 221240 6458
rect 221188 6394 221240 6400
rect 221200 6322 221228 6394
rect 221370 6352 221426 6361
rect 221188 6316 221240 6322
rect 221370 6287 221372 6296
rect 221188 6258 221240 6264
rect 221424 6287 221426 6296
rect 221464 6316 221516 6322
rect 221372 6258 221424 6264
rect 221464 6258 221516 6264
rect 221476 6225 221504 6258
rect 221462 6216 221518 6225
rect 221462 6151 221518 6160
rect 221004 5908 221056 5914
rect 221004 5850 221056 5856
rect 221004 2984 221056 2990
rect 221004 2926 221056 2932
rect 221016 2514 221044 2926
rect 221004 2508 221056 2514
rect 221004 2450 221056 2456
rect 221372 2440 221424 2446
rect 221372 2382 221424 2388
rect 221384 2310 221412 2382
rect 221372 2304 221424 2310
rect 221372 2246 221424 2252
rect 221004 1896 221056 1902
rect 221002 1864 221004 1873
rect 221056 1864 221058 1873
rect 221002 1799 221058 1808
rect 221188 1352 221240 1358
rect 221188 1294 221240 1300
rect 220912 1216 220964 1222
rect 220912 1158 220964 1164
rect 221200 746 221228 1294
rect 221568 814 221596 7346
rect 221752 6866 221780 7346
rect 221922 7304 221978 7313
rect 221922 7239 221978 7248
rect 221936 6866 221964 7239
rect 222120 6866 222148 9386
rect 222212 9110 222240 9386
rect 222844 9376 222896 9382
rect 222844 9318 222896 9324
rect 222936 9376 222988 9382
rect 222936 9318 222988 9324
rect 222200 9104 222252 9110
rect 222200 9046 222252 9052
rect 222856 7410 222884 9318
rect 222844 7404 222896 7410
rect 222844 7346 222896 7352
rect 222198 7304 222254 7313
rect 222198 7239 222254 7248
rect 221740 6860 221792 6866
rect 221740 6802 221792 6808
rect 221924 6860 221976 6866
rect 221924 6802 221976 6808
rect 222108 6860 222160 6866
rect 222108 6802 222160 6808
rect 221752 6225 221780 6802
rect 221844 6730 222148 6746
rect 221844 6724 222160 6730
rect 221844 6718 222108 6724
rect 221738 6216 221794 6225
rect 221738 6151 221794 6160
rect 221648 4072 221700 4078
rect 221648 4014 221700 4020
rect 221660 2378 221688 4014
rect 221648 2372 221700 2378
rect 221648 2314 221700 2320
rect 221844 2106 221872 6718
rect 222108 6666 222160 6672
rect 222016 6656 222068 6662
rect 222016 6598 222068 6604
rect 222028 5778 222056 6598
rect 222108 6384 222160 6390
rect 222108 6326 222160 6332
rect 222120 6225 222148 6326
rect 222106 6216 222162 6225
rect 222106 6151 222162 6160
rect 222016 5772 222068 5778
rect 222016 5714 222068 5720
rect 222016 5636 222068 5642
rect 222016 5578 222068 5584
rect 222028 4758 222056 5578
rect 222016 4752 222068 4758
rect 222016 4694 222068 4700
rect 222028 4554 222056 4694
rect 222016 4548 222068 4554
rect 222016 4490 222068 4496
rect 222016 4276 222068 4282
rect 222016 4218 222068 4224
rect 221924 2644 221976 2650
rect 221924 2586 221976 2592
rect 221936 2514 221964 2586
rect 221924 2508 221976 2514
rect 221924 2450 221976 2456
rect 221832 2100 221884 2106
rect 221832 2042 221884 2048
rect 222028 882 222056 4218
rect 222212 3097 222240 7239
rect 222384 7200 222436 7206
rect 222384 7142 222436 7148
rect 222292 6792 222344 6798
rect 222292 6734 222344 6740
rect 222304 5642 222332 6734
rect 222292 5636 222344 5642
rect 222292 5578 222344 5584
rect 222290 5264 222346 5273
rect 222396 5234 222424 7142
rect 222844 5636 222896 5642
rect 222844 5578 222896 5584
rect 222290 5199 222292 5208
rect 222344 5199 222346 5208
rect 222384 5228 222436 5234
rect 222292 5170 222344 5176
rect 222384 5170 222436 5176
rect 222476 4820 222528 4826
rect 222476 4762 222528 4768
rect 222488 4622 222516 4762
rect 222476 4616 222528 4622
rect 222476 4558 222528 4564
rect 222752 3528 222804 3534
rect 222752 3470 222804 3476
rect 222198 3088 222254 3097
rect 222198 3023 222254 3032
rect 222476 2304 222528 2310
rect 222476 2246 222528 2252
rect 222568 2304 222620 2310
rect 222568 2246 222620 2252
rect 222106 2136 222162 2145
rect 222106 2071 222162 2080
rect 222120 1902 222148 2071
rect 222488 1970 222516 2246
rect 222580 2038 222608 2246
rect 222568 2032 222620 2038
rect 222568 1974 222620 1980
rect 222476 1964 222528 1970
rect 222476 1906 222528 1912
rect 222108 1896 222160 1902
rect 222108 1838 222160 1844
rect 222200 1352 222252 1358
rect 222764 1329 222792 3470
rect 222200 1294 222252 1300
rect 222750 1320 222806 1329
rect 222212 921 222240 1294
rect 222292 1284 222344 1290
rect 222750 1255 222806 1264
rect 222292 1226 222344 1232
rect 222198 912 222254 921
rect 222016 876 222068 882
rect 222198 847 222254 856
rect 222016 818 222068 824
rect 221556 808 221608 814
rect 221556 750 221608 756
rect 221188 740 221240 746
rect 221188 682 221240 688
rect 219624 400 219676 406
rect 217876 342 217928 348
rect 218886 368 218942 377
rect 216220 332 216272 338
rect 218886 303 218942 312
rect 219622 368 219624 377
rect 220728 400 220780 406
rect 219676 368 219678 377
rect 222304 377 222332 1226
rect 222382 1184 222438 1193
rect 222382 1119 222438 1128
rect 222396 921 222424 1119
rect 222382 912 222438 921
rect 222382 847 222438 856
rect 220728 342 220780 348
rect 222290 368 222346 377
rect 219622 303 219678 312
rect 222290 303 222346 312
rect 216220 274 216272 280
rect 222856 270 222884 5578
rect 222948 4078 222976 9318
rect 223486 9208 223542 9217
rect 223486 9143 223542 9152
rect 223500 9110 223528 9143
rect 223488 9104 223540 9110
rect 223488 9046 223540 9052
rect 224420 9042 224448 9454
rect 224774 9415 224830 9424
rect 224408 9036 224460 9042
rect 224408 8978 224460 8984
rect 224040 8968 224092 8974
rect 224040 8910 224092 8916
rect 224684 8968 224736 8974
rect 224788 8956 224816 9415
rect 225144 9376 225196 9382
rect 225144 9318 225196 9324
rect 224736 8928 224816 8956
rect 224684 8910 224736 8916
rect 223946 8800 224002 8809
rect 223946 8735 224002 8744
rect 223960 8566 223988 8735
rect 223948 8560 224000 8566
rect 223948 8502 224000 8508
rect 224052 8514 224080 8910
rect 224788 8566 224816 8928
rect 224776 8560 224828 8566
rect 223672 8492 223724 8498
rect 224052 8486 224448 8514
rect 224776 8502 224828 8508
rect 224868 8560 224920 8566
rect 224868 8502 224920 8508
rect 223672 8434 223724 8440
rect 223488 8424 223540 8430
rect 223488 8366 223540 8372
rect 223396 7948 223448 7954
rect 223396 7890 223448 7896
rect 223120 7336 223172 7342
rect 223120 7278 223172 7284
rect 222936 4072 222988 4078
rect 222936 4014 222988 4020
rect 223028 2440 223080 2446
rect 223028 2382 223080 2388
rect 223040 2106 223068 2382
rect 223028 2100 223080 2106
rect 223028 2042 223080 2048
rect 223040 610 223068 2042
rect 223132 1222 223160 7278
rect 223304 7268 223356 7274
rect 223304 7210 223356 7216
rect 223316 6866 223344 7210
rect 223304 6860 223356 6866
rect 223304 6802 223356 6808
rect 223316 5642 223344 6802
rect 223408 6322 223436 7890
rect 223396 6316 223448 6322
rect 223396 6258 223448 6264
rect 223408 6225 223436 6258
rect 223394 6216 223450 6225
rect 223394 6151 223450 6160
rect 223396 5840 223448 5846
rect 223396 5782 223448 5788
rect 223304 5636 223356 5642
rect 223304 5578 223356 5584
rect 223212 4820 223264 4826
rect 223212 4762 223264 4768
rect 223224 4185 223252 4762
rect 223408 4593 223436 5782
rect 223394 4584 223450 4593
rect 223394 4519 223450 4528
rect 223500 4468 223528 8366
rect 223580 8288 223632 8294
rect 223580 8230 223632 8236
rect 223592 7886 223620 8230
rect 223580 7880 223632 7886
rect 223580 7822 223632 7828
rect 223684 7426 223712 8434
rect 224314 7848 224370 7857
rect 224314 7783 224370 7792
rect 223854 7576 223910 7585
rect 223854 7511 223910 7520
rect 223592 7398 223712 7426
rect 223868 7410 223896 7511
rect 223856 7404 223908 7410
rect 223592 5710 223620 7398
rect 223856 7346 223908 7352
rect 223948 7336 224000 7342
rect 223948 7278 224000 7284
rect 224132 7336 224184 7342
rect 224132 7278 224184 7284
rect 223764 6792 223816 6798
rect 223764 6734 223816 6740
rect 223856 6792 223908 6798
rect 223856 6734 223908 6740
rect 223672 6656 223724 6662
rect 223672 6598 223724 6604
rect 223684 6322 223712 6598
rect 223672 6316 223724 6322
rect 223672 6258 223724 6264
rect 223776 5914 223804 6734
rect 223868 6390 223896 6734
rect 223856 6384 223908 6390
rect 223856 6326 223908 6332
rect 223856 6248 223908 6254
rect 223856 6190 223908 6196
rect 223764 5908 223816 5914
rect 223764 5850 223816 5856
rect 223580 5704 223632 5710
rect 223580 5646 223632 5652
rect 223868 5166 223896 6190
rect 223856 5160 223908 5166
rect 223856 5102 223908 5108
rect 223672 4548 223724 4554
rect 223672 4490 223724 4496
rect 223408 4440 223528 4468
rect 223210 4176 223266 4185
rect 223210 4111 223266 4120
rect 223210 3088 223266 3097
rect 223210 3023 223212 3032
rect 223264 3023 223266 3032
rect 223304 3052 223356 3058
rect 223212 2994 223264 3000
rect 223304 2994 223356 3000
rect 223316 2825 223344 2994
rect 223302 2816 223358 2825
rect 223302 2751 223358 2760
rect 223408 2417 223436 4440
rect 223580 2984 223632 2990
rect 223580 2926 223632 2932
rect 223488 2848 223540 2854
rect 223488 2790 223540 2796
rect 223500 2689 223528 2790
rect 223486 2680 223542 2689
rect 223486 2615 223542 2624
rect 223592 2514 223620 2926
rect 223580 2508 223632 2514
rect 223580 2450 223632 2456
rect 223684 2446 223712 4490
rect 223854 2680 223910 2689
rect 223854 2615 223910 2624
rect 223672 2440 223724 2446
rect 223394 2408 223450 2417
rect 223672 2382 223724 2388
rect 223394 2343 223450 2352
rect 223210 2136 223266 2145
rect 223210 2071 223266 2080
rect 223224 1970 223252 2071
rect 223212 1964 223264 1970
rect 223212 1906 223264 1912
rect 223408 1601 223436 2343
rect 223764 2304 223816 2310
rect 223764 2246 223816 2252
rect 223394 1592 223450 1601
rect 223394 1527 223450 1536
rect 223578 1592 223634 1601
rect 223578 1527 223634 1536
rect 223120 1216 223172 1222
rect 223120 1158 223172 1164
rect 223592 950 223620 1527
rect 223776 1358 223804 2246
rect 223868 1834 223896 2615
rect 223960 2530 223988 7278
rect 224144 6390 224172 7278
rect 224132 6384 224184 6390
rect 224132 6326 224184 6332
rect 224132 6248 224184 6254
rect 224130 6216 224132 6225
rect 224184 6216 224186 6225
rect 224130 6151 224186 6160
rect 224224 6180 224276 6186
rect 224224 6122 224276 6128
rect 224236 5914 224264 6122
rect 224224 5908 224276 5914
rect 224224 5850 224276 5856
rect 223960 2502 224172 2530
rect 224040 2372 224092 2378
rect 224040 2314 224092 2320
rect 223946 2272 224002 2281
rect 223946 2207 224002 2216
rect 223960 2038 223988 2207
rect 223948 2032 224000 2038
rect 223948 1974 224000 1980
rect 223856 1828 223908 1834
rect 223856 1770 223908 1776
rect 224052 1465 224080 2314
rect 224038 1456 224094 1465
rect 224038 1391 224094 1400
rect 223764 1352 223816 1358
rect 223764 1294 223816 1300
rect 224040 1284 224092 1290
rect 224040 1226 224092 1232
rect 223580 944 223632 950
rect 223580 886 223632 892
rect 223028 604 223080 610
rect 223028 546 223080 552
rect 223120 604 223172 610
rect 223120 546 223172 552
rect 223132 338 223160 546
rect 223120 332 223172 338
rect 223120 274 223172 280
rect 222844 264 222896 270
rect 224052 241 224080 1226
rect 224144 406 224172 2502
rect 224224 2304 224276 2310
rect 224224 2246 224276 2252
rect 224236 2106 224264 2246
rect 224224 2100 224276 2106
rect 224224 2042 224276 2048
rect 224328 1766 224356 7783
rect 224420 1970 224448 8486
rect 224774 8392 224830 8401
rect 224774 8327 224776 8336
rect 224828 8327 224830 8336
rect 224776 8298 224828 8304
rect 224880 7041 224908 8502
rect 224958 7576 225014 7585
rect 224958 7511 225014 7520
rect 224972 7342 225000 7511
rect 224960 7336 225012 7342
rect 224960 7278 225012 7284
rect 224866 7032 224922 7041
rect 224866 6967 224922 6976
rect 224960 6928 225012 6934
rect 224958 6896 224960 6905
rect 225012 6896 225014 6905
rect 224868 6860 224920 6866
rect 224958 6831 225014 6840
rect 224868 6802 224920 6808
rect 224592 6656 224644 6662
rect 224592 6598 224644 6604
rect 224604 5846 224632 6598
rect 224880 6225 224908 6802
rect 224866 6216 224922 6225
rect 224866 6151 224922 6160
rect 224592 5840 224644 5846
rect 224592 5782 224644 5788
rect 225052 5704 225104 5710
rect 225052 5646 225104 5652
rect 224868 5636 224920 5642
rect 224868 5578 224920 5584
rect 224684 5296 224736 5302
rect 224684 5238 224736 5244
rect 224696 4826 224724 5238
rect 224880 5114 224908 5578
rect 224880 5086 225000 5114
rect 224868 5024 224920 5030
rect 224868 4966 224920 4972
rect 224880 4865 224908 4966
rect 224866 4856 224922 4865
rect 224684 4820 224736 4826
rect 224866 4791 224922 4800
rect 224684 4762 224736 4768
rect 224696 4321 224724 4762
rect 224682 4312 224738 4321
rect 224682 4247 224738 4256
rect 224500 4072 224552 4078
rect 224500 4014 224552 4020
rect 224512 3738 224540 4014
rect 224972 4010 225000 5086
rect 224960 4004 225012 4010
rect 224960 3946 225012 3952
rect 224500 3732 224552 3738
rect 224500 3674 224552 3680
rect 224972 3602 225000 3946
rect 224960 3596 225012 3602
rect 224960 3538 225012 3544
rect 224866 2816 224922 2825
rect 224922 2774 225000 2802
rect 224866 2751 224922 2760
rect 224972 2650 225000 2774
rect 224960 2644 225012 2650
rect 224960 2586 225012 2592
rect 224682 2544 224738 2553
rect 224682 2479 224738 2488
rect 224696 2281 224724 2479
rect 224682 2272 224738 2281
rect 224682 2207 224738 2216
rect 224408 1964 224460 1970
rect 224408 1906 224460 1912
rect 224776 1964 224828 1970
rect 224776 1906 224828 1912
rect 224316 1760 224368 1766
rect 224788 1737 224816 1906
rect 224868 1896 224920 1902
rect 224868 1838 224920 1844
rect 224316 1702 224368 1708
rect 224774 1728 224830 1737
rect 224774 1663 224830 1672
rect 224788 1494 224816 1663
rect 224776 1488 224828 1494
rect 224776 1430 224828 1436
rect 224880 1034 224908 1838
rect 225064 1222 225092 5646
rect 225156 3602 225184 9318
rect 225236 6996 225288 7002
rect 225236 6938 225288 6944
rect 225248 5030 225276 6938
rect 225328 6384 225380 6390
rect 225328 6326 225380 6332
rect 225340 6254 225368 6326
rect 225328 6248 225380 6254
rect 225328 6190 225380 6196
rect 225236 5024 225288 5030
rect 225236 4966 225288 4972
rect 225236 4072 225288 4078
rect 225236 4014 225288 4020
rect 225328 4072 225380 4078
rect 225328 4014 225380 4020
rect 225248 3738 225276 4014
rect 225236 3732 225288 3738
rect 225236 3674 225288 3680
rect 225144 3596 225196 3602
rect 225144 3538 225196 3544
rect 225340 2530 225368 4014
rect 225248 2502 225368 2530
rect 225248 2281 225276 2502
rect 225328 2440 225380 2446
rect 225328 2382 225380 2388
rect 225234 2272 225290 2281
rect 225234 2207 225290 2216
rect 225340 2106 225368 2382
rect 225328 2100 225380 2106
rect 225328 2042 225380 2048
rect 225432 1426 225460 10474
rect 225512 10328 225564 10334
rect 225512 10270 225564 10276
rect 225524 10130 225552 10270
rect 225512 10124 225564 10130
rect 225512 10066 225564 10072
rect 225604 10124 225656 10130
rect 225604 10066 225656 10072
rect 225616 9178 225644 10066
rect 225694 9752 225750 9761
rect 225694 9687 225696 9696
rect 225748 9687 225750 9696
rect 225696 9658 225748 9664
rect 225970 9480 226026 9489
rect 225970 9415 226026 9424
rect 225696 9376 225748 9382
rect 225696 9318 225748 9324
rect 225604 9172 225656 9178
rect 225604 9114 225656 9120
rect 225604 8968 225656 8974
rect 225602 8936 225604 8945
rect 225656 8936 225658 8945
rect 225602 8871 225658 8880
rect 225708 8838 225736 9318
rect 225880 9104 225932 9110
rect 225880 9046 225932 9052
rect 225696 8832 225748 8838
rect 225696 8774 225748 8780
rect 225788 8832 225840 8838
rect 225788 8774 225840 8780
rect 225800 8498 225828 8774
rect 225892 8634 225920 9046
rect 225984 9042 226012 9415
rect 225972 9036 226024 9042
rect 225972 8978 226024 8984
rect 226444 8974 226472 10610
rect 227536 10600 227588 10606
rect 227536 10542 227588 10548
rect 227548 9722 227576 10542
rect 227720 10532 227772 10538
rect 227720 10474 227772 10480
rect 227732 10334 227760 10474
rect 227720 10328 227772 10334
rect 227720 10270 227772 10276
rect 228088 10328 228140 10334
rect 228088 10270 228140 10276
rect 227536 9716 227588 9722
rect 227536 9658 227588 9664
rect 226432 8968 226484 8974
rect 227260 8968 227312 8974
rect 226432 8910 226484 8916
rect 227166 8936 227222 8945
rect 225970 8664 226026 8673
rect 225880 8628 225932 8634
rect 225970 8599 225972 8608
rect 225880 8570 225932 8576
rect 226024 8599 226026 8608
rect 225972 8570 226024 8576
rect 225788 8492 225840 8498
rect 225788 8434 225840 8440
rect 226444 8362 226472 8910
rect 227732 8956 227760 10270
rect 228100 9382 228128 10270
rect 229112 9722 229140 10814
rect 233700 10872 233752 10878
rect 233608 10814 233660 10820
rect 233698 10840 233700 10849
rect 246764 10872 246816 10878
rect 233752 10840 233754 10849
rect 231858 10775 231914 10784
rect 230848 10532 230900 10538
rect 230848 10474 230900 10480
rect 230860 10334 230888 10474
rect 230848 10328 230900 10334
rect 230848 10270 230900 10276
rect 230664 10260 230716 10266
rect 230664 10202 230716 10208
rect 229192 9920 229244 9926
rect 229192 9862 229244 9868
rect 229468 9920 229520 9926
rect 229468 9862 229520 9868
rect 229204 9722 229232 9862
rect 229100 9716 229152 9722
rect 229100 9658 229152 9664
rect 229192 9716 229244 9722
rect 229192 9658 229244 9664
rect 228364 9580 228416 9586
rect 228364 9522 228416 9528
rect 228270 9480 228326 9489
rect 228270 9415 228326 9424
rect 228284 9382 228312 9415
rect 228088 9376 228140 9382
rect 228088 9318 228140 9324
rect 228272 9376 228324 9382
rect 228272 9318 228324 9324
rect 228100 8974 228128 9318
rect 228376 9178 228404 9522
rect 228364 9172 228416 9178
rect 228364 9114 228416 9120
rect 228456 9172 228508 9178
rect 228456 9114 228508 9120
rect 228088 8968 228140 8974
rect 227312 8928 227852 8956
rect 227260 8910 227312 8916
rect 227166 8871 227222 8880
rect 226524 8832 226576 8838
rect 226524 8774 226576 8780
rect 226536 8498 226564 8774
rect 226706 8664 226762 8673
rect 226706 8599 226708 8608
rect 226760 8599 226762 8608
rect 226708 8570 226760 8576
rect 226524 8492 226576 8498
rect 226524 8434 226576 8440
rect 226432 8356 226484 8362
rect 226432 8298 226484 8304
rect 227076 8356 227128 8362
rect 227076 8298 227128 8304
rect 226338 8256 226394 8265
rect 226338 8191 226394 8200
rect 225880 8084 225932 8090
rect 225880 8026 225932 8032
rect 225512 7268 225564 7274
rect 225512 7210 225564 7216
rect 225524 6866 225552 7210
rect 225512 6860 225564 6866
rect 225512 6802 225564 6808
rect 225604 6452 225656 6458
rect 225604 6394 225656 6400
rect 225616 6225 225644 6394
rect 225892 6322 225920 8026
rect 226064 7880 226116 7886
rect 226064 7822 226116 7828
rect 225972 6724 226024 6730
rect 225972 6666 226024 6672
rect 225880 6316 225932 6322
rect 225880 6258 225932 6264
rect 225602 6216 225658 6225
rect 225602 6151 225658 6160
rect 225984 5166 226012 6666
rect 226076 6322 226104 7822
rect 226248 6996 226300 7002
rect 226248 6938 226300 6944
rect 226260 6497 226288 6938
rect 226352 6934 226380 8191
rect 226984 7472 227036 7478
rect 226984 7414 227036 7420
rect 226996 7206 227024 7414
rect 226984 7200 227036 7206
rect 226984 7142 227036 7148
rect 226340 6928 226392 6934
rect 226340 6870 226392 6876
rect 226246 6488 226302 6497
rect 226246 6423 226302 6432
rect 226984 6384 227036 6390
rect 226064 6316 226116 6322
rect 226064 6258 226116 6264
rect 226444 6310 226932 6338
rect 226984 6326 227036 6332
rect 226076 5778 226104 6258
rect 226338 6216 226394 6225
rect 226248 6180 226300 6186
rect 226338 6151 226394 6160
rect 226248 6122 226300 6128
rect 226260 5914 226288 6122
rect 226156 5908 226208 5914
rect 226156 5850 226208 5856
rect 226248 5908 226300 5914
rect 226248 5850 226300 5856
rect 226168 5794 226196 5850
rect 226064 5772 226116 5778
rect 226168 5766 226288 5794
rect 226064 5714 226116 5720
rect 226260 5522 226288 5766
rect 226352 5681 226380 6151
rect 226444 6118 226472 6310
rect 226708 6248 226760 6254
rect 226708 6190 226760 6196
rect 226432 6112 226484 6118
rect 226432 6054 226484 6060
rect 226524 6112 226576 6118
rect 226524 6054 226576 6060
rect 226536 5710 226564 6054
rect 226720 5710 226748 6190
rect 226524 5704 226576 5710
rect 226338 5672 226394 5681
rect 226708 5704 226760 5710
rect 226524 5646 226576 5652
rect 226614 5672 226670 5681
rect 226338 5607 226394 5616
rect 226708 5646 226760 5652
rect 226614 5607 226670 5616
rect 226260 5494 226380 5522
rect 225972 5160 226024 5166
rect 225972 5102 226024 5108
rect 226352 5098 226380 5494
rect 226628 5250 226656 5607
rect 226444 5222 226656 5250
rect 226340 5092 226392 5098
rect 226340 5034 226392 5040
rect 226444 4978 226472 5222
rect 225616 4950 226472 4978
rect 225616 3466 225644 4950
rect 226340 4820 226392 4826
rect 226340 4762 226392 4768
rect 226156 4616 226208 4622
rect 226156 4558 226208 4564
rect 226246 4584 226302 4593
rect 225878 4176 225934 4185
rect 226168 4146 226196 4558
rect 226246 4519 226248 4528
rect 226300 4519 226302 4528
rect 226248 4490 226300 4496
rect 225878 4111 225934 4120
rect 226156 4140 226208 4146
rect 225892 4060 225920 4111
rect 226156 4082 226208 4088
rect 226064 4072 226116 4078
rect 225892 4032 226064 4060
rect 226064 4014 226116 4020
rect 226352 3754 226380 4762
rect 226616 4480 226668 4486
rect 226616 4422 226668 4428
rect 226628 4214 226656 4422
rect 226616 4208 226668 4214
rect 226720 4185 226748 5646
rect 226800 5160 226852 5166
rect 226800 5102 226852 5108
rect 226812 4554 226840 5102
rect 226800 4548 226852 4554
rect 226800 4490 226852 4496
rect 226616 4150 226668 4156
rect 226706 4176 226762 4185
rect 226706 4111 226762 4120
rect 226616 4004 226668 4010
rect 226720 3992 226748 4111
rect 226668 3964 226748 3992
rect 226616 3946 226668 3952
rect 226168 3726 226380 3754
rect 226168 3602 226196 3726
rect 226248 3664 226300 3670
rect 226248 3606 226300 3612
rect 226156 3596 226208 3602
rect 226156 3538 226208 3544
rect 225696 3528 225748 3534
rect 225696 3470 225748 3476
rect 225604 3460 225656 3466
rect 225604 3402 225656 3408
rect 225708 3194 225736 3470
rect 226260 3194 226288 3606
rect 226720 3534 226748 3964
rect 226904 3942 226932 6310
rect 226996 6186 227024 6326
rect 226984 6180 227036 6186
rect 226984 6122 227036 6128
rect 226984 4072 227036 4078
rect 226984 4014 227036 4020
rect 226800 3936 226852 3942
rect 226800 3878 226852 3884
rect 226892 3936 226944 3942
rect 226892 3878 226944 3884
rect 226432 3528 226484 3534
rect 226432 3470 226484 3476
rect 226708 3528 226760 3534
rect 226708 3470 226760 3476
rect 225696 3188 225748 3194
rect 225696 3130 225748 3136
rect 226248 3188 226300 3194
rect 226248 3130 226300 3136
rect 226064 3120 226116 3126
rect 226064 3062 226116 3068
rect 226076 2990 226104 3062
rect 226064 2984 226116 2990
rect 226064 2926 226116 2932
rect 226246 2816 226302 2825
rect 226246 2751 226302 2760
rect 226260 2650 226288 2751
rect 226248 2644 226300 2650
rect 226248 2586 226300 2592
rect 226156 2440 226208 2446
rect 225878 2408 225934 2417
rect 226156 2382 226208 2388
rect 226248 2440 226300 2446
rect 226248 2382 226300 2388
rect 225878 2343 225934 2352
rect 225604 2304 225656 2310
rect 225604 2246 225656 2252
rect 225512 2032 225564 2038
rect 225512 1974 225564 1980
rect 225524 1766 225552 1974
rect 225512 1760 225564 1766
rect 225512 1702 225564 1708
rect 225616 1465 225644 2246
rect 225892 1970 225920 2343
rect 226168 2106 226196 2382
rect 226156 2100 226208 2106
rect 226156 2042 226208 2048
rect 225880 1964 225932 1970
rect 225880 1906 225932 1912
rect 226260 1562 226288 2382
rect 226444 1562 226472 3470
rect 226812 3126 226840 3878
rect 226996 3126 227024 4014
rect 226800 3120 226852 3126
rect 226800 3062 226852 3068
rect 226984 3120 227036 3126
rect 226984 3062 227036 3068
rect 226892 3052 226944 3058
rect 226892 2994 226944 3000
rect 226524 2848 226576 2854
rect 226522 2816 226524 2825
rect 226576 2816 226578 2825
rect 226522 2751 226578 2760
rect 226708 2304 226760 2310
rect 226708 2246 226760 2252
rect 226720 1970 226748 2246
rect 226708 1964 226760 1970
rect 226708 1906 226760 1912
rect 226616 1896 226668 1902
rect 226616 1838 226668 1844
rect 226248 1556 226300 1562
rect 226248 1498 226300 1504
rect 226432 1556 226484 1562
rect 226432 1498 226484 1504
rect 225602 1456 225658 1465
rect 225420 1420 225472 1426
rect 225602 1391 225658 1400
rect 225420 1362 225472 1368
rect 226628 1358 226656 1838
rect 226904 1358 226932 2994
rect 226984 2440 227036 2446
rect 226984 2382 227036 2388
rect 226996 2106 227024 2382
rect 226984 2100 227036 2106
rect 226984 2042 227036 2048
rect 227088 1426 227116 8298
rect 227180 2310 227208 8871
rect 227626 8120 227682 8129
rect 227626 8055 227628 8064
rect 227680 8055 227682 8064
rect 227628 8026 227680 8032
rect 227628 7812 227680 7818
rect 227628 7754 227680 7760
rect 227640 6798 227668 7754
rect 227628 6792 227680 6798
rect 227628 6734 227680 6740
rect 227640 5914 227668 6734
rect 227720 6384 227772 6390
rect 227720 6326 227772 6332
rect 227732 6118 227760 6326
rect 227720 6112 227772 6118
rect 227720 6054 227772 6060
rect 227628 5908 227680 5914
rect 227628 5850 227680 5856
rect 227732 5710 227760 6054
rect 227720 5704 227772 5710
rect 227720 5646 227772 5652
rect 227352 5568 227404 5574
rect 227352 5510 227404 5516
rect 227364 5302 227392 5510
rect 227352 5296 227404 5302
rect 227352 5238 227404 5244
rect 227536 5296 227588 5302
rect 227536 5238 227588 5244
rect 227548 5030 227576 5238
rect 227536 5024 227588 5030
rect 227536 4966 227588 4972
rect 227720 5024 227772 5030
rect 227720 4966 227772 4972
rect 227732 4865 227760 4966
rect 227718 4856 227774 4865
rect 227718 4791 227774 4800
rect 227352 4072 227404 4078
rect 227352 4014 227404 4020
rect 227364 3738 227392 4014
rect 227444 3936 227496 3942
rect 227442 3904 227444 3913
rect 227496 3904 227498 3913
rect 227442 3839 227498 3848
rect 227352 3732 227404 3738
rect 227352 3674 227404 3680
rect 227720 3596 227772 3602
rect 227720 3538 227772 3544
rect 227732 3398 227760 3538
rect 227720 3392 227772 3398
rect 227720 3334 227772 3340
rect 227628 2984 227680 2990
rect 227628 2926 227680 2932
rect 227260 2848 227312 2854
rect 227260 2790 227312 2796
rect 227168 2304 227220 2310
rect 227168 2246 227220 2252
rect 227076 1420 227128 1426
rect 227076 1362 227128 1368
rect 226616 1352 226668 1358
rect 226616 1294 226668 1300
rect 226892 1352 226944 1358
rect 227272 1329 227300 2790
rect 227640 2446 227668 2926
rect 227824 2774 227852 8928
rect 228008 8928 228088 8956
rect 228008 4706 228036 8928
rect 228468 8945 228496 9114
rect 229112 8974 229140 9658
rect 229480 9518 229508 9862
rect 229834 9752 229890 9761
rect 230676 9722 230704 10202
rect 231582 9752 231638 9761
rect 229834 9687 229836 9696
rect 229888 9687 229890 9696
rect 230664 9716 230716 9722
rect 229836 9658 229888 9664
rect 231582 9687 231638 9696
rect 230664 9658 230716 9664
rect 230020 9580 230072 9586
rect 230020 9522 230072 9528
rect 230204 9580 230256 9586
rect 230204 9522 230256 9528
rect 229468 9512 229520 9518
rect 229468 9454 229520 9460
rect 228824 8968 228876 8974
rect 228088 8910 228140 8916
rect 228454 8936 228510 8945
rect 228824 8910 228876 8916
rect 229100 8968 229152 8974
rect 229100 8910 229152 8916
rect 228454 8871 228510 8880
rect 228088 8832 228140 8838
rect 228836 8809 228864 8910
rect 228916 8832 228968 8838
rect 228088 8774 228140 8780
rect 228822 8800 228878 8809
rect 228100 8498 228128 8774
rect 228916 8774 228968 8780
rect 228822 8735 228878 8744
rect 228270 8664 228326 8673
rect 228270 8599 228272 8608
rect 228324 8599 228326 8608
rect 228272 8570 228324 8576
rect 228088 8492 228140 8498
rect 228088 8434 228140 8440
rect 228088 7744 228140 7750
rect 228088 7686 228140 7692
rect 228100 6089 228128 7686
rect 228180 6656 228232 6662
rect 228180 6598 228232 6604
rect 228086 6080 228142 6089
rect 228086 6015 228142 6024
rect 228100 5710 228128 6015
rect 228088 5704 228140 5710
rect 228088 5646 228140 5652
rect 228192 4865 228220 6598
rect 228456 6248 228508 6254
rect 228456 6190 228508 6196
rect 228468 5642 228496 6190
rect 228456 5636 228508 5642
rect 228456 5578 228508 5584
rect 228836 5522 228864 8735
rect 228928 8498 228956 8774
rect 229098 8664 229154 8673
rect 229098 8599 229100 8608
rect 229152 8599 229154 8608
rect 229100 8570 229152 8576
rect 229480 8498 229508 9454
rect 229836 9376 229888 9382
rect 229836 9318 229888 9324
rect 229848 8974 229876 9318
rect 230032 9042 230060 9522
rect 230020 9036 230072 9042
rect 230020 8978 230072 8984
rect 230216 8974 230244 9522
rect 229652 8968 229704 8974
rect 229652 8910 229704 8916
rect 229836 8968 229888 8974
rect 229836 8910 229888 8916
rect 230204 8968 230256 8974
rect 230204 8910 230256 8916
rect 228916 8492 228968 8498
rect 228916 8434 228968 8440
rect 229468 8492 229520 8498
rect 229468 8434 229520 8440
rect 229560 8424 229612 8430
rect 229560 8366 229612 8372
rect 228916 8288 228968 8294
rect 228916 8230 228968 8236
rect 228928 5642 228956 8230
rect 229192 6996 229244 7002
rect 229192 6938 229244 6944
rect 229008 6724 229060 6730
rect 229008 6666 229060 6672
rect 228916 5636 228968 5642
rect 228916 5578 228968 5584
rect 228836 5494 228956 5522
rect 228272 5296 228324 5302
rect 228270 5264 228272 5273
rect 228824 5296 228876 5302
rect 228324 5264 228326 5273
rect 228824 5238 228876 5244
rect 228270 5199 228326 5208
rect 228178 4856 228234 4865
rect 228178 4791 228234 4800
rect 228272 4752 228324 4758
rect 228008 4678 228220 4706
rect 228272 4694 228324 4700
rect 227902 3768 227958 3777
rect 227902 3703 227958 3712
rect 227732 2746 227852 2774
rect 227628 2440 227680 2446
rect 227628 2382 227680 2388
rect 227732 1970 227760 2746
rect 227812 2372 227864 2378
rect 227812 2314 227864 2320
rect 227720 1964 227772 1970
rect 227720 1906 227772 1912
rect 227824 1494 227852 2314
rect 227812 1488 227864 1494
rect 227812 1430 227864 1436
rect 226892 1294 226944 1300
rect 227258 1320 227314 1329
rect 226248 1284 226300 1290
rect 227258 1255 227314 1264
rect 226248 1226 226300 1232
rect 225052 1216 225104 1222
rect 225052 1158 225104 1164
rect 224880 1006 225000 1034
rect 224868 944 224920 950
rect 224868 886 224920 892
rect 224776 740 224828 746
rect 224776 682 224828 688
rect 224132 400 224184 406
rect 224132 342 224184 348
rect 222844 206 222896 212
rect 224038 232 224094 241
rect 224038 167 224094 176
rect 224788 105 224816 682
rect 224880 377 224908 886
rect 224866 368 224922 377
rect 224866 303 224922 312
rect 224972 105 225000 1006
rect 226260 950 226288 1226
rect 226248 944 226300 950
rect 226248 886 226300 892
rect 227916 338 227944 3703
rect 228088 3052 228140 3058
rect 228088 2994 228140 3000
rect 227996 2644 228048 2650
rect 227996 2586 228048 2592
rect 228008 474 228036 2586
rect 228100 2106 228128 2994
rect 228088 2100 228140 2106
rect 228088 2042 228140 2048
rect 228192 1426 228220 4678
rect 228284 4486 228312 4694
rect 228836 4622 228864 5238
rect 228824 4616 228876 4622
rect 228730 4584 228786 4593
rect 228824 4558 228876 4564
rect 228730 4519 228732 4528
rect 228784 4519 228786 4528
rect 228732 4490 228784 4496
rect 228272 4480 228324 4486
rect 228272 4422 228324 4428
rect 228284 4078 228312 4422
rect 228272 4072 228324 4078
rect 228272 4014 228324 4020
rect 228362 3496 228418 3505
rect 228362 3431 228418 3440
rect 228272 2848 228324 2854
rect 228272 2790 228324 2796
rect 228180 1420 228232 1426
rect 228180 1362 228232 1368
rect 228284 1329 228312 2790
rect 228376 2446 228404 3431
rect 228364 2440 228416 2446
rect 228364 2382 228416 2388
rect 228824 2440 228876 2446
rect 228824 2382 228876 2388
rect 228456 2304 228508 2310
rect 228456 2246 228508 2252
rect 228364 1896 228416 1902
rect 228364 1838 228416 1844
rect 228376 1358 228404 1838
rect 228364 1352 228416 1358
rect 228270 1320 228326 1329
rect 228364 1294 228416 1300
rect 228270 1255 228326 1264
rect 228468 1193 228496 2246
rect 228836 1562 228864 2382
rect 228928 1970 228956 5494
rect 229020 5030 229048 6666
rect 229008 5024 229060 5030
rect 229008 4966 229060 4972
rect 229100 4072 229152 4078
rect 229100 4014 229152 4020
rect 229112 3913 229140 4014
rect 229098 3904 229154 3913
rect 229098 3839 229154 3848
rect 229204 3466 229232 6938
rect 229572 6866 229600 8366
rect 229560 6860 229612 6866
rect 229560 6802 229612 6808
rect 229572 5914 229600 6802
rect 229560 5908 229612 5914
rect 229560 5850 229612 5856
rect 229192 3460 229244 3466
rect 229192 3402 229244 3408
rect 229192 2100 229244 2106
rect 229192 2042 229244 2048
rect 228916 1964 228968 1970
rect 228916 1906 228968 1912
rect 229204 1766 229232 2042
rect 229468 1964 229520 1970
rect 229664 1952 229692 8910
rect 229848 8566 229876 8910
rect 230110 8800 230166 8809
rect 230110 8735 230166 8744
rect 230124 8566 230152 8735
rect 229836 8560 229888 8566
rect 229836 8502 229888 8508
rect 230112 8560 230164 8566
rect 230112 8502 230164 8508
rect 229928 8492 229980 8498
rect 229928 8434 229980 8440
rect 229836 8424 229888 8430
rect 229836 8366 229888 8372
rect 229742 7848 229798 7857
rect 229742 7783 229798 7792
rect 229756 7585 229784 7783
rect 229742 7576 229798 7585
rect 229742 7511 229798 7520
rect 229848 6118 229876 8366
rect 229836 6112 229888 6118
rect 229836 6054 229888 6060
rect 229940 5642 229968 8434
rect 230112 7404 230164 7410
rect 230112 7346 230164 7352
rect 230124 7002 230152 7346
rect 230216 7206 230244 8910
rect 230676 8498 230704 9658
rect 231032 9580 231084 9586
rect 231032 9522 231084 9528
rect 230848 9036 230900 9042
rect 230848 8978 230900 8984
rect 230860 8498 230888 8978
rect 231044 8634 231072 9522
rect 231596 9382 231624 9687
rect 231584 9376 231636 9382
rect 231584 9318 231636 9324
rect 231872 8974 231900 10775
rect 233620 10606 233648 10814
rect 246764 10814 246816 10820
rect 258540 10872 258592 10878
rect 258540 10814 258592 10820
rect 267832 10872 267884 10878
rect 267832 10814 267884 10820
rect 233698 10775 233754 10784
rect 239404 10804 239456 10810
rect 239404 10746 239456 10752
rect 233792 10668 233844 10674
rect 233792 10610 233844 10616
rect 233424 10600 233476 10606
rect 233424 10542 233476 10548
rect 233608 10600 233660 10606
rect 233608 10542 233660 10548
rect 232872 9648 232924 9654
rect 232872 9590 232924 9596
rect 232884 9382 232912 9590
rect 232872 9376 232924 9382
rect 232872 9318 232924 9324
rect 232884 8974 232912 9318
rect 233436 9110 233464 10542
rect 233700 10124 233752 10130
rect 233700 10066 233752 10072
rect 233514 9752 233570 9761
rect 233514 9687 233516 9696
rect 233568 9687 233570 9696
rect 233516 9658 233568 9664
rect 233332 9104 233384 9110
rect 233332 9046 233384 9052
rect 233424 9104 233476 9110
rect 233424 9046 233476 9052
rect 231860 8968 231912 8974
rect 231860 8910 231912 8916
rect 232136 8968 232188 8974
rect 232136 8910 232188 8916
rect 232504 8968 232556 8974
rect 232504 8910 232556 8916
rect 232872 8968 232924 8974
rect 232872 8910 232924 8916
rect 231768 8832 231820 8838
rect 231768 8774 231820 8780
rect 231032 8628 231084 8634
rect 231032 8570 231084 8576
rect 231780 8498 231808 8774
rect 231950 8664 232006 8673
rect 231950 8599 231952 8608
rect 232004 8599 232006 8608
rect 231952 8570 232004 8576
rect 230664 8492 230716 8498
rect 230664 8434 230716 8440
rect 230848 8492 230900 8498
rect 230848 8434 230900 8440
rect 231768 8492 231820 8498
rect 231768 8434 231820 8440
rect 231032 8424 231084 8430
rect 230846 8392 230902 8401
rect 230572 8356 230624 8362
rect 231032 8366 231084 8372
rect 230846 8327 230902 8336
rect 230572 8298 230624 8304
rect 230388 8084 230440 8090
rect 230388 8026 230440 8032
rect 230294 7440 230350 7449
rect 230294 7375 230296 7384
rect 230348 7375 230350 7384
rect 230296 7346 230348 7352
rect 230204 7200 230256 7206
rect 230204 7142 230256 7148
rect 230296 7200 230348 7206
rect 230296 7142 230348 7148
rect 230112 6996 230164 7002
rect 230112 6938 230164 6944
rect 230308 6322 230336 7142
rect 230400 6497 230428 8026
rect 230584 7886 230612 8298
rect 230860 8090 230888 8327
rect 230848 8084 230900 8090
rect 230848 8026 230900 8032
rect 230572 7880 230624 7886
rect 230572 7822 230624 7828
rect 230480 6996 230532 7002
rect 230480 6938 230532 6944
rect 230492 6798 230520 6938
rect 230848 6928 230900 6934
rect 230848 6870 230900 6876
rect 230480 6792 230532 6798
rect 230480 6734 230532 6740
rect 230480 6656 230532 6662
rect 230480 6598 230532 6604
rect 230386 6488 230442 6497
rect 230386 6423 230442 6432
rect 230296 6316 230348 6322
rect 230296 6258 230348 6264
rect 230492 6118 230520 6598
rect 230112 6112 230164 6118
rect 230112 6054 230164 6060
rect 230480 6112 230532 6118
rect 230480 6054 230532 6060
rect 230756 6112 230808 6118
rect 230756 6054 230808 6060
rect 230020 5704 230072 5710
rect 230020 5646 230072 5652
rect 229836 5636 229888 5642
rect 229836 5578 229888 5584
rect 229928 5636 229980 5642
rect 229928 5578 229980 5584
rect 229742 4992 229798 5001
rect 229742 4927 229798 4936
rect 229756 4826 229784 4927
rect 229744 4820 229796 4826
rect 229744 4762 229796 4768
rect 229848 4146 229876 5578
rect 230032 5234 230060 5646
rect 230020 5228 230072 5234
rect 230020 5170 230072 5176
rect 229836 4140 229888 4146
rect 229836 4082 229888 4088
rect 229836 3392 229888 3398
rect 229836 3334 229888 3340
rect 229848 2922 229876 3334
rect 229836 2916 229888 2922
rect 229836 2858 229888 2864
rect 229834 2272 229890 2281
rect 229834 2207 229890 2216
rect 229744 1964 229796 1970
rect 229664 1924 229744 1952
rect 229468 1906 229520 1912
rect 229744 1906 229796 1912
rect 229480 1850 229508 1906
rect 229848 1902 229876 2207
rect 230124 1970 230152 6054
rect 230664 5636 230716 5642
rect 230664 5578 230716 5584
rect 230294 5400 230350 5409
rect 230570 5400 230626 5409
rect 230350 5358 230520 5386
rect 230294 5335 230350 5344
rect 230492 5234 230520 5358
rect 230570 5335 230626 5344
rect 230480 5228 230532 5234
rect 230480 5170 230532 5176
rect 230584 5114 230612 5335
rect 230216 5086 230612 5114
rect 230676 5098 230704 5578
rect 230664 5092 230716 5098
rect 229928 1964 229980 1970
rect 229928 1906 229980 1912
rect 230112 1964 230164 1970
rect 230112 1906 230164 1912
rect 229836 1896 229888 1902
rect 229480 1822 229784 1850
rect 229836 1838 229888 1844
rect 229192 1760 229244 1766
rect 229192 1702 229244 1708
rect 229284 1760 229336 1766
rect 229284 1702 229336 1708
rect 229652 1760 229704 1766
rect 229756 1748 229784 1822
rect 229940 1748 229968 1906
rect 229756 1720 229968 1748
rect 229652 1702 229704 1708
rect 228824 1556 228876 1562
rect 228824 1498 228876 1504
rect 229296 1358 229324 1702
rect 229664 1358 229692 1702
rect 229284 1352 229336 1358
rect 229284 1294 229336 1300
rect 229652 1352 229704 1358
rect 229652 1294 229704 1300
rect 230216 1290 230244 5086
rect 230664 5034 230716 5040
rect 230768 4758 230796 6054
rect 230860 5642 230888 6870
rect 230848 5636 230900 5642
rect 230848 5578 230900 5584
rect 230860 5302 230888 5578
rect 230848 5296 230900 5302
rect 230848 5238 230900 5244
rect 231044 5250 231072 8366
rect 231216 7812 231268 7818
rect 231216 7754 231268 7760
rect 231228 7410 231256 7754
rect 231216 7404 231268 7410
rect 231216 7346 231268 7352
rect 231308 7404 231360 7410
rect 231308 7346 231360 7352
rect 231124 6792 231176 6798
rect 231124 6734 231176 6740
rect 231136 6118 231164 6734
rect 231124 6112 231176 6118
rect 231124 6054 231176 6060
rect 231320 5914 231348 7346
rect 231768 6724 231820 6730
rect 231768 6666 231820 6672
rect 231780 6633 231808 6666
rect 231490 6624 231546 6633
rect 231490 6559 231546 6568
rect 231766 6624 231822 6633
rect 231766 6559 231822 6568
rect 231308 5908 231360 5914
rect 231308 5850 231360 5856
rect 231400 5908 231452 5914
rect 231400 5850 231452 5856
rect 231412 5794 231440 5850
rect 231216 5772 231268 5778
rect 231216 5714 231268 5720
rect 231320 5766 231440 5794
rect 231044 5222 231164 5250
rect 231032 5092 231084 5098
rect 231032 5034 231084 5040
rect 230756 4752 230808 4758
rect 230756 4694 230808 4700
rect 230756 4548 230808 4554
rect 230756 4490 230808 4496
rect 230296 4480 230348 4486
rect 230296 4422 230348 4428
rect 230308 4078 230336 4422
rect 230768 4185 230796 4490
rect 231044 4214 231072 5034
rect 231032 4208 231084 4214
rect 230754 4176 230810 4185
rect 231032 4150 231084 4156
rect 230754 4111 230810 4120
rect 230768 4078 230796 4111
rect 230296 4072 230348 4078
rect 230296 4014 230348 4020
rect 230756 4072 230808 4078
rect 230756 4014 230808 4020
rect 230480 4004 230532 4010
rect 230664 4004 230716 4010
rect 230532 3964 230664 3992
rect 230480 3946 230532 3952
rect 230664 3946 230716 3952
rect 231032 3936 231084 3942
rect 231032 3878 231084 3884
rect 230756 3392 230808 3398
rect 230756 3334 230808 3340
rect 230388 3120 230440 3126
rect 230388 3062 230440 3068
rect 230400 1290 230428 3062
rect 230768 1970 230796 3334
rect 231044 2825 231072 3878
rect 231030 2816 231086 2825
rect 231030 2751 231086 2760
rect 231136 2774 231164 5222
rect 231228 4622 231256 5714
rect 231320 5030 231348 5766
rect 231504 5710 231532 6559
rect 231596 6310 231808 6338
rect 231596 6254 231624 6310
rect 231780 6254 231808 6310
rect 231584 6248 231636 6254
rect 231584 6190 231636 6196
rect 231676 6248 231728 6254
rect 231676 6190 231728 6196
rect 231768 6248 231820 6254
rect 231768 6190 231820 6196
rect 231688 5817 231716 6190
rect 231674 5808 231730 5817
rect 231674 5743 231730 5752
rect 231860 5772 231912 5778
rect 231860 5714 231912 5720
rect 231492 5704 231544 5710
rect 231492 5646 231544 5652
rect 231308 5024 231360 5030
rect 231308 4966 231360 4972
rect 231216 4616 231268 4622
rect 231216 4558 231268 4564
rect 231320 4146 231348 4966
rect 231504 4622 231532 5646
rect 231872 5234 231900 5714
rect 231860 5228 231912 5234
rect 231860 5170 231912 5176
rect 231492 4616 231544 4622
rect 231492 4558 231544 4564
rect 231492 4480 231544 4486
rect 231492 4422 231544 4428
rect 231308 4140 231360 4146
rect 231308 4082 231360 4088
rect 231504 3534 231532 4422
rect 231492 3528 231544 3534
rect 231492 3470 231544 3476
rect 231676 2848 231728 2854
rect 231676 2790 231728 2796
rect 231136 2746 231532 2774
rect 231308 2304 231360 2310
rect 231308 2246 231360 2252
rect 230756 1964 230808 1970
rect 230756 1906 230808 1912
rect 230664 1760 230716 1766
rect 230664 1702 230716 1708
rect 230676 1358 230704 1702
rect 230664 1352 230716 1358
rect 230664 1294 230716 1300
rect 230204 1284 230256 1290
rect 230204 1226 230256 1232
rect 230388 1284 230440 1290
rect 230388 1226 230440 1232
rect 229100 1216 229152 1222
rect 228454 1184 228510 1193
rect 229100 1158 229152 1164
rect 229836 1216 229888 1222
rect 229836 1158 229888 1164
rect 230848 1216 230900 1222
rect 231320 1193 231348 2246
rect 231504 1970 231532 2746
rect 231688 2650 231716 2790
rect 231676 2644 231728 2650
rect 231676 2586 231728 2592
rect 231768 2440 231820 2446
rect 231768 2382 231820 2388
rect 231860 2440 231912 2446
rect 231860 2382 231912 2388
rect 231780 2038 231808 2382
rect 231872 2038 231900 2382
rect 232044 2304 232096 2310
rect 232044 2246 232096 2252
rect 231768 2032 231820 2038
rect 231768 1974 231820 1980
rect 231860 2032 231912 2038
rect 231860 1974 231912 1980
rect 231492 1964 231544 1970
rect 231492 1906 231544 1912
rect 231584 1964 231636 1970
rect 231584 1906 231636 1912
rect 231596 1766 231624 1906
rect 231584 1760 231636 1766
rect 231584 1702 231636 1708
rect 232056 1193 232084 2246
rect 232148 1970 232176 8910
rect 232318 5808 232374 5817
rect 232318 5743 232374 5752
rect 232332 5710 232360 5743
rect 232320 5704 232372 5710
rect 232320 5646 232372 5652
rect 232136 1964 232188 1970
rect 232136 1906 232188 1912
rect 232320 1964 232372 1970
rect 232320 1906 232372 1912
rect 232332 1766 232360 1906
rect 232320 1760 232372 1766
rect 232320 1702 232372 1708
rect 232332 1358 232360 1702
rect 232516 1426 232544 8910
rect 233344 8838 233372 9046
rect 233712 8974 233740 10066
rect 233804 9178 233832 10610
rect 235724 10396 235776 10402
rect 235724 10338 235776 10344
rect 234342 9752 234398 9761
rect 234342 9687 234344 9696
rect 234396 9687 234398 9696
rect 235078 9752 235134 9761
rect 235078 9687 235080 9696
rect 234344 9658 234396 9664
rect 235132 9687 235134 9696
rect 235080 9658 235132 9664
rect 234068 9580 234120 9586
rect 234068 9522 234120 9528
rect 234160 9580 234212 9586
rect 234160 9522 234212 9528
rect 234896 9580 234948 9586
rect 234896 9522 234948 9528
rect 234080 9178 234108 9522
rect 234172 9178 234200 9522
rect 234620 9444 234672 9450
rect 234620 9386 234672 9392
rect 233792 9172 233844 9178
rect 233792 9114 233844 9120
rect 234068 9172 234120 9178
rect 234068 9114 234120 9120
rect 234160 9172 234212 9178
rect 234160 9114 234212 9120
rect 233700 8968 233752 8974
rect 233700 8910 233752 8916
rect 234528 8968 234580 8974
rect 234528 8910 234580 8916
rect 233240 8832 233292 8838
rect 233240 8774 233292 8780
rect 233332 8832 233384 8838
rect 233332 8774 233384 8780
rect 232870 8664 232926 8673
rect 232870 8599 232872 8608
rect 232924 8599 232926 8608
rect 232872 8570 232924 8576
rect 233252 8498 233280 8774
rect 233240 8492 233292 8498
rect 233240 8434 233292 8440
rect 232596 2440 232648 2446
rect 232596 2382 232648 2388
rect 232608 1562 232636 2382
rect 232780 2304 232832 2310
rect 232780 2246 232832 2252
rect 232596 1556 232648 1562
rect 232596 1498 232648 1504
rect 232504 1420 232556 1426
rect 232504 1362 232556 1368
rect 232320 1352 232372 1358
rect 232320 1294 232372 1300
rect 232792 1193 232820 2246
rect 233712 2038 233740 8910
rect 234540 8838 234568 8910
rect 234068 8832 234120 8838
rect 234068 8774 234120 8780
rect 234528 8832 234580 8838
rect 234528 8774 234580 8780
rect 233700 2032 233752 2038
rect 233700 1974 233752 1980
rect 233884 2032 233936 2038
rect 233884 1974 233936 1980
rect 233240 1964 233292 1970
rect 233424 1964 233476 1970
rect 233292 1924 233424 1952
rect 233240 1906 233292 1912
rect 233424 1906 233476 1912
rect 233896 1766 233924 1974
rect 234080 1902 234108 8774
rect 234528 8492 234580 8498
rect 234632 8480 234660 9386
rect 234908 8634 234936 9522
rect 235448 9512 235500 9518
rect 235448 9454 235500 9460
rect 234896 8628 234948 8634
rect 234896 8570 234948 8576
rect 234580 8452 234660 8480
rect 234528 8434 234580 8440
rect 234540 8362 234568 8434
rect 235262 8392 235318 8401
rect 234528 8356 234580 8362
rect 234528 8298 234580 8304
rect 234896 8356 234948 8362
rect 235262 8327 235318 8336
rect 234896 8298 234948 8304
rect 234908 1970 234936 8298
rect 235276 7410 235304 8327
rect 235264 7404 235316 7410
rect 235264 7346 235316 7352
rect 235356 7404 235408 7410
rect 235356 7346 235408 7352
rect 235368 5681 235396 7346
rect 235354 5672 235410 5681
rect 235354 5607 235410 5616
rect 234896 1964 234948 1970
rect 234896 1906 234948 1912
rect 234068 1896 234120 1902
rect 234068 1838 234120 1844
rect 233240 1760 233292 1766
rect 233240 1702 233292 1708
rect 233884 1760 233936 1766
rect 233884 1702 233936 1708
rect 233976 1760 234028 1766
rect 233976 1702 234028 1708
rect 234712 1760 234764 1766
rect 234712 1702 234764 1708
rect 233252 1358 233280 1702
rect 233988 1358 234016 1702
rect 234724 1358 234752 1702
rect 235460 1426 235488 9454
rect 235540 9444 235592 9450
rect 235540 9386 235592 9392
rect 235552 3942 235580 9386
rect 235632 8968 235684 8974
rect 235736 8956 235764 10338
rect 235816 9716 235868 9722
rect 235816 9658 235868 9664
rect 236552 9716 236604 9722
rect 236552 9658 236604 9664
rect 235828 9586 235856 9658
rect 235816 9580 235868 9586
rect 235816 9522 235868 9528
rect 235908 9580 235960 9586
rect 235908 9522 235960 9528
rect 235920 8974 235948 9522
rect 236564 9382 236592 9658
rect 236184 9376 236236 9382
rect 236184 9318 236236 9324
rect 236552 9376 236604 9382
rect 236552 9318 236604 9324
rect 237196 9376 237248 9382
rect 237196 9318 237248 9324
rect 238116 9376 238168 9382
rect 238116 9318 238168 9324
rect 235998 9208 236054 9217
rect 235998 9143 236000 9152
rect 236052 9143 236054 9152
rect 236000 9114 236052 9120
rect 236092 9036 236144 9042
rect 236092 8978 236144 8984
rect 235816 8968 235868 8974
rect 235736 8928 235816 8956
rect 235632 8910 235684 8916
rect 235816 8910 235868 8916
rect 235908 8968 235960 8974
rect 235908 8910 235960 8916
rect 235644 8838 235672 8910
rect 235632 8832 235684 8838
rect 235632 8774 235684 8780
rect 235724 8492 235776 8498
rect 235724 8434 235776 8440
rect 235736 7886 235764 8434
rect 235828 8294 235856 8910
rect 235920 8498 235948 8910
rect 236104 8634 236132 8978
rect 236092 8628 236144 8634
rect 236092 8570 236144 8576
rect 236196 8498 236224 9318
rect 236368 8832 236420 8838
rect 236368 8774 236420 8780
rect 236552 8832 236604 8838
rect 236552 8774 236604 8780
rect 235908 8492 235960 8498
rect 235908 8434 235960 8440
rect 236184 8492 236236 8498
rect 236184 8434 236236 8440
rect 236380 8430 236408 8774
rect 236368 8424 236420 8430
rect 236368 8366 236420 8372
rect 236564 8294 236592 8774
rect 236642 8664 236698 8673
rect 236642 8599 236644 8608
rect 236696 8599 236698 8608
rect 236644 8570 236696 8576
rect 235816 8288 235868 8294
rect 235816 8230 235868 8236
rect 236552 8288 236604 8294
rect 236552 8230 236604 8236
rect 236920 8288 236972 8294
rect 236920 8230 236972 8236
rect 237102 8256 237158 8265
rect 235724 7880 235776 7886
rect 235724 7822 235776 7828
rect 236092 7744 236144 7750
rect 236092 7686 236144 7692
rect 236184 7744 236236 7750
rect 236184 7686 236236 7692
rect 236000 7404 236052 7410
rect 236000 7346 236052 7352
rect 236012 7206 236040 7346
rect 236104 7342 236132 7686
rect 236196 7410 236224 7686
rect 236184 7404 236236 7410
rect 236184 7346 236236 7352
rect 236092 7336 236144 7342
rect 236092 7278 236144 7284
rect 235632 7200 235684 7206
rect 235632 7142 235684 7148
rect 236000 7200 236052 7206
rect 236000 7142 236052 7148
rect 235644 6322 235672 7142
rect 236564 6934 236592 8230
rect 236736 8016 236788 8022
rect 236736 7958 236788 7964
rect 235724 6928 235776 6934
rect 235724 6870 235776 6876
rect 236552 6928 236604 6934
rect 236552 6870 236604 6876
rect 235632 6316 235684 6322
rect 235632 6258 235684 6264
rect 235632 5024 235684 5030
rect 235632 4966 235684 4972
rect 235644 4214 235672 4966
rect 235632 4208 235684 4214
rect 235632 4150 235684 4156
rect 235540 3936 235592 3942
rect 235540 3878 235592 3884
rect 235736 1902 235764 6870
rect 235816 2984 235868 2990
rect 235816 2926 235868 2932
rect 236092 2984 236144 2990
rect 236092 2926 236144 2932
rect 235828 1902 235856 2926
rect 235906 2816 235962 2825
rect 235962 2774 236040 2802
rect 235906 2751 235962 2760
rect 236012 2650 236040 2774
rect 236104 2689 236132 2926
rect 236090 2680 236146 2689
rect 236000 2644 236052 2650
rect 236748 2650 236776 7958
rect 236932 7546 236960 8230
rect 237102 8191 237158 8200
rect 237012 7880 237064 7886
rect 237010 7848 237012 7857
rect 237064 7848 237066 7857
rect 237010 7783 237066 7792
rect 236920 7540 236972 7546
rect 236920 7482 236972 7488
rect 236920 6996 236972 7002
rect 236920 6938 236972 6944
rect 236932 4146 236960 6938
rect 237010 6896 237066 6905
rect 237010 6831 237066 6840
rect 237024 5953 237052 6831
rect 237116 6610 237144 8191
rect 237208 8022 237236 9318
rect 237539 9276 237847 9285
rect 237539 9274 237545 9276
rect 237601 9274 237625 9276
rect 237681 9274 237705 9276
rect 237761 9274 237785 9276
rect 237841 9274 237847 9276
rect 237601 9222 237603 9274
rect 237783 9222 237785 9274
rect 237539 9220 237545 9222
rect 237601 9220 237625 9222
rect 237681 9220 237705 9222
rect 237761 9220 237785 9222
rect 237841 9220 237847 9222
rect 237286 9208 237342 9217
rect 237539 9211 237847 9220
rect 237286 9143 237288 9152
rect 237340 9143 237342 9152
rect 237932 9172 237984 9178
rect 237288 9114 237340 9120
rect 237932 9114 237984 9120
rect 237944 8362 237972 9114
rect 237932 8356 237984 8362
rect 237932 8298 237984 8304
rect 237539 8188 237847 8197
rect 237539 8186 237545 8188
rect 237601 8186 237625 8188
rect 237681 8186 237705 8188
rect 237761 8186 237785 8188
rect 237841 8186 237847 8188
rect 237601 8134 237603 8186
rect 237783 8134 237785 8186
rect 237539 8132 237545 8134
rect 237601 8132 237625 8134
rect 237681 8132 237705 8134
rect 237761 8132 237785 8134
rect 237841 8132 237847 8134
rect 237539 8123 237847 8132
rect 237930 8120 237986 8129
rect 237930 8055 237986 8064
rect 237196 8016 237248 8022
rect 237196 7958 237248 7964
rect 237654 7984 237710 7993
rect 237654 7919 237710 7928
rect 237838 7984 237894 7993
rect 237838 7919 237894 7928
rect 237380 7880 237432 7886
rect 237380 7822 237432 7828
rect 237196 7540 237248 7546
rect 237196 7482 237248 7488
rect 237208 7177 237236 7482
rect 237286 7440 237342 7449
rect 237392 7410 237420 7822
rect 237668 7750 237696 7919
rect 237852 7886 237880 7919
rect 237840 7880 237892 7886
rect 237944 7857 237972 8055
rect 238024 7880 238076 7886
rect 237840 7822 237892 7828
rect 237930 7848 237986 7857
rect 238024 7822 238076 7828
rect 237930 7783 237986 7792
rect 237656 7744 237708 7750
rect 237656 7686 237708 7692
rect 238036 7410 238064 7822
rect 237286 7375 237288 7384
rect 237340 7375 237342 7384
rect 237380 7404 237432 7410
rect 237288 7346 237340 7352
rect 237380 7346 237432 7352
rect 238024 7404 238076 7410
rect 238024 7346 238076 7352
rect 237392 7290 237420 7346
rect 237300 7262 237420 7290
rect 237300 7206 237328 7262
rect 237288 7200 237340 7206
rect 237194 7168 237250 7177
rect 237288 7142 237340 7148
rect 237380 7200 237432 7206
rect 237380 7142 237432 7148
rect 237194 7103 237250 7112
rect 237300 6882 237328 7142
rect 237208 6854 237328 6882
rect 237392 6866 237420 7142
rect 237539 7100 237847 7109
rect 237539 7098 237545 7100
rect 237601 7098 237625 7100
rect 237681 7098 237705 7100
rect 237761 7098 237785 7100
rect 237841 7098 237847 7100
rect 237601 7046 237603 7098
rect 237783 7046 237785 7098
rect 237539 7044 237545 7046
rect 237601 7044 237625 7046
rect 237681 7044 237705 7046
rect 237761 7044 237785 7046
rect 237841 7044 237847 7046
rect 237539 7035 237847 7044
rect 237380 6860 237432 6866
rect 237208 6798 237236 6854
rect 237380 6802 237432 6808
rect 237196 6792 237248 6798
rect 237196 6734 237248 6740
rect 237300 6730 237512 6746
rect 237300 6724 237524 6730
rect 237300 6718 237472 6724
rect 237300 6610 237328 6718
rect 237472 6666 237524 6672
rect 237116 6582 237328 6610
rect 237380 6656 237432 6662
rect 237380 6598 237432 6604
rect 237392 6322 237420 6598
rect 237380 6316 237432 6322
rect 237380 6258 237432 6264
rect 237539 6012 237847 6021
rect 237539 6010 237545 6012
rect 237601 6010 237625 6012
rect 237681 6010 237705 6012
rect 237761 6010 237785 6012
rect 237841 6010 237847 6012
rect 237601 5958 237603 6010
rect 237783 5958 237785 6010
rect 237539 5956 237545 5958
rect 237601 5956 237625 5958
rect 237681 5956 237705 5958
rect 237761 5956 237785 5958
rect 237841 5956 237847 5958
rect 237010 5944 237066 5953
rect 237539 5947 237847 5956
rect 237010 5879 237066 5888
rect 237380 5636 237432 5642
rect 237380 5578 237432 5584
rect 237392 4978 237420 5578
rect 237208 4950 237420 4978
rect 237208 4826 237236 4950
rect 237539 4924 237847 4933
rect 237539 4922 237545 4924
rect 237601 4922 237625 4924
rect 237681 4922 237705 4924
rect 237761 4922 237785 4924
rect 237841 4922 237847 4924
rect 237601 4870 237603 4922
rect 237783 4870 237785 4922
rect 237539 4868 237545 4870
rect 237601 4868 237625 4870
rect 237681 4868 237705 4870
rect 237761 4868 237785 4870
rect 237841 4868 237847 4870
rect 237286 4856 237342 4865
rect 237539 4859 237847 4868
rect 237196 4820 237248 4826
rect 237286 4791 237288 4800
rect 237196 4762 237248 4768
rect 237340 4791 237342 4800
rect 237288 4762 237340 4768
rect 236920 4140 236972 4146
rect 236920 4082 236972 4088
rect 237380 4072 237432 4078
rect 237380 4014 237432 4020
rect 236090 2615 236146 2624
rect 236736 2644 236788 2650
rect 236000 2586 236052 2592
rect 236736 2586 236788 2592
rect 236092 2440 236144 2446
rect 236092 2382 236144 2388
rect 236552 2440 236604 2446
rect 236552 2382 236604 2388
rect 235998 2272 236054 2281
rect 235998 2207 236054 2216
rect 236012 2106 236040 2207
rect 236104 2106 236132 2382
rect 236000 2100 236052 2106
rect 236000 2042 236052 2048
rect 236092 2100 236144 2106
rect 236092 2042 236144 2048
rect 236000 1964 236052 1970
rect 236000 1906 236052 1912
rect 235724 1896 235776 1902
rect 235724 1838 235776 1844
rect 235816 1896 235868 1902
rect 235816 1838 235868 1844
rect 235722 1592 235778 1601
rect 235722 1527 235778 1536
rect 235448 1420 235500 1426
rect 235448 1362 235500 1368
rect 233240 1352 233292 1358
rect 233240 1294 233292 1300
rect 233976 1352 234028 1358
rect 234712 1352 234764 1358
rect 233976 1294 234028 1300
rect 234618 1320 234674 1329
rect 234712 1294 234764 1300
rect 234618 1255 234674 1264
rect 233424 1216 233476 1222
rect 230848 1158 230900 1164
rect 231306 1184 231362 1193
rect 228454 1119 228510 1128
rect 227996 468 228048 474
rect 227996 410 228048 416
rect 229112 377 229140 1158
rect 229744 944 229796 950
rect 229744 886 229796 892
rect 229098 368 229154 377
rect 227904 332 227956 338
rect 229098 303 229154 312
rect 227904 274 227956 280
rect 229756 270 229784 886
rect 229848 377 229876 1158
rect 230860 377 230888 1158
rect 231306 1119 231362 1128
rect 232042 1184 232098 1193
rect 232042 1119 232098 1128
rect 232778 1184 232834 1193
rect 233424 1158 233476 1164
rect 234160 1216 234212 1222
rect 234160 1158 234212 1164
rect 232778 1119 232834 1128
rect 233436 377 233464 1158
rect 234172 377 234200 1158
rect 234632 513 234660 1255
rect 234896 1216 234948 1222
rect 234896 1158 234948 1164
rect 234908 513 234936 1158
rect 234618 504 234674 513
rect 234618 439 234674 448
rect 234894 504 234950 513
rect 234894 439 234950 448
rect 235736 406 235764 1527
rect 236012 1358 236040 1906
rect 236564 1562 236592 2382
rect 237196 2372 237248 2378
rect 237196 2314 237248 2320
rect 236736 2304 236788 2310
rect 236736 2246 236788 2252
rect 236552 1556 236604 1562
rect 236552 1498 236604 1504
rect 236000 1352 236052 1358
rect 236000 1294 236052 1300
rect 236748 1193 236776 2246
rect 237208 1426 237236 2314
rect 237288 1760 237340 1766
rect 237288 1702 237340 1708
rect 237300 1465 237328 1702
rect 237286 1456 237342 1465
rect 237196 1420 237248 1426
rect 237286 1391 237342 1400
rect 237196 1362 237248 1368
rect 237392 1290 237420 4014
rect 237539 3836 237847 3845
rect 237539 3834 237545 3836
rect 237601 3834 237625 3836
rect 237681 3834 237705 3836
rect 237761 3834 237785 3836
rect 237841 3834 237847 3836
rect 237601 3782 237603 3834
rect 237783 3782 237785 3834
rect 237539 3780 237545 3782
rect 237601 3780 237625 3782
rect 237681 3780 237705 3782
rect 237761 3780 237785 3782
rect 237841 3780 237847 3782
rect 237539 3771 237847 3780
rect 237930 3768 237986 3777
rect 237930 3703 237986 3712
rect 237944 3618 237972 3703
rect 238128 3641 238156 9318
rect 238760 8968 238812 8974
rect 238760 8910 238812 8916
rect 238576 8356 238628 8362
rect 238576 8298 238628 8304
rect 238206 4040 238262 4049
rect 238206 3975 238262 3984
rect 237852 3590 237972 3618
rect 238114 3632 238170 3641
rect 237852 3369 237880 3590
rect 238114 3567 238170 3576
rect 237838 3360 237894 3369
rect 237838 3295 237894 3304
rect 238220 2774 238248 3975
rect 238588 3670 238616 8298
rect 238772 7585 238800 8910
rect 239036 8016 239088 8022
rect 239036 7958 239088 7964
rect 238942 7848 238998 7857
rect 238942 7783 238998 7792
rect 238758 7576 238814 7585
rect 238956 7546 238984 7783
rect 239048 7585 239076 7958
rect 239416 7886 239444 10746
rect 239678 10296 239734 10305
rect 239678 10231 239734 10240
rect 240230 10296 240286 10305
rect 240230 10231 240286 10240
rect 241242 10296 241298 10305
rect 241242 10231 241298 10240
rect 241978 10296 242034 10305
rect 241978 10231 242034 10240
rect 242714 10296 242770 10305
rect 242714 10231 242770 10240
rect 243450 10296 243506 10305
rect 243450 10231 243506 10240
rect 244186 10296 244242 10305
rect 244186 10231 244242 10240
rect 244922 10296 244978 10305
rect 244922 10231 244978 10240
rect 246118 10296 246174 10305
rect 246118 10231 246174 10240
rect 246394 10296 246450 10305
rect 246394 10231 246450 10240
rect 239692 9586 239720 10231
rect 240244 9654 240272 10231
rect 240232 9648 240284 9654
rect 240232 9590 240284 9596
rect 241256 9586 241284 10231
rect 239680 9580 239732 9586
rect 239680 9522 239732 9528
rect 241244 9580 241296 9586
rect 241244 9522 241296 9528
rect 241520 9512 241572 9518
rect 241520 9454 241572 9460
rect 239404 7880 239456 7886
rect 239404 7822 239456 7828
rect 239034 7576 239090 7585
rect 238758 7511 238814 7520
rect 238944 7540 238996 7546
rect 239034 7511 239090 7520
rect 238944 7482 238996 7488
rect 238668 7404 238720 7410
rect 238668 7346 238720 7352
rect 238680 5370 238708 7346
rect 239128 7336 239180 7342
rect 239128 7278 239180 7284
rect 239140 7206 239168 7278
rect 238760 7200 238812 7206
rect 238760 7142 238812 7148
rect 239128 7200 239180 7206
rect 239128 7142 239180 7148
rect 238772 6118 238800 7142
rect 239140 6662 239168 7142
rect 239128 6656 239180 6662
rect 239128 6598 239180 6604
rect 238760 6112 238812 6118
rect 238760 6054 238812 6060
rect 238668 5364 238720 5370
rect 238668 5306 238720 5312
rect 239232 5358 239720 5386
rect 238680 5234 238708 5306
rect 239232 5302 239260 5358
rect 239692 5302 239720 5358
rect 239220 5296 239272 5302
rect 239680 5296 239732 5302
rect 239220 5238 239272 5244
rect 239324 5234 239628 5250
rect 239680 5238 239732 5244
rect 240322 5264 240378 5273
rect 238668 5228 238720 5234
rect 238668 5170 238720 5176
rect 239312 5228 239640 5234
rect 239364 5222 239588 5228
rect 239312 5170 239364 5176
rect 240322 5199 240378 5208
rect 240506 5264 240562 5273
rect 240506 5199 240562 5208
rect 239588 5170 239640 5176
rect 239220 5160 239272 5166
rect 239272 5108 239352 5114
rect 239220 5102 239352 5108
rect 239232 5086 239352 5102
rect 239220 5024 239272 5030
rect 239324 5012 239352 5086
rect 239588 5024 239640 5030
rect 239324 4984 239588 5012
rect 239220 4966 239272 4972
rect 239588 4966 239640 4972
rect 239232 4622 239260 4966
rect 240336 4826 240364 5199
rect 240324 4820 240376 4826
rect 240324 4762 240376 4768
rect 239220 4616 239272 4622
rect 239220 4558 239272 4564
rect 239680 4480 239732 4486
rect 239680 4422 239732 4428
rect 239692 4214 239720 4422
rect 240048 4276 240100 4282
rect 240048 4218 240100 4224
rect 239680 4208 239732 4214
rect 239680 4150 239732 4156
rect 238576 3664 238628 3670
rect 238576 3606 238628 3612
rect 238666 3224 238722 3233
rect 238666 3159 238722 3168
rect 238680 2854 238708 3159
rect 238668 2848 238720 2854
rect 238668 2790 238720 2796
rect 237539 2748 237847 2757
rect 237539 2746 237545 2748
rect 237601 2746 237625 2748
rect 237681 2746 237705 2748
rect 237761 2746 237785 2748
rect 237841 2746 237847 2748
rect 237601 2694 237603 2746
rect 237783 2694 237785 2746
rect 237539 2692 237545 2694
rect 237601 2692 237625 2694
rect 237681 2692 237705 2694
rect 237761 2692 237785 2694
rect 237841 2692 237847 2694
rect 237539 2683 237847 2692
rect 237944 2746 238248 2774
rect 237944 1970 237972 2746
rect 240060 1970 240088 4218
rect 240520 3233 240548 5199
rect 240968 4820 241020 4826
rect 240968 4762 241020 4768
rect 240980 4622 241008 4762
rect 240968 4616 241020 4622
rect 240968 4558 241020 4564
rect 240784 4140 240836 4146
rect 240784 4082 240836 4088
rect 240796 4049 240824 4082
rect 240782 4040 240838 4049
rect 240782 3975 240838 3984
rect 241532 3369 241560 9454
rect 241992 9042 242020 10231
rect 242728 9586 242756 10231
rect 243084 10056 243136 10062
rect 243084 9998 243136 10004
rect 242716 9580 242768 9586
rect 242716 9522 242768 9528
rect 241980 9036 242032 9042
rect 241980 8978 242032 8984
rect 242992 8628 243044 8634
rect 242992 8570 243044 8576
rect 242900 8424 242952 8430
rect 242900 8366 242952 8372
rect 242912 8022 242940 8366
rect 242900 8016 242952 8022
rect 242900 7958 242952 7964
rect 242900 7744 242952 7750
rect 243004 7721 243032 8570
rect 243096 8090 243124 9998
rect 243176 9376 243228 9382
rect 243176 9318 243228 9324
rect 243188 8294 243216 9318
rect 243464 9042 243492 10231
rect 243820 9512 243872 9518
rect 243820 9454 243872 9460
rect 243544 9444 243596 9450
rect 243544 9386 243596 9392
rect 243556 9042 243584 9386
rect 243452 9036 243504 9042
rect 243452 8978 243504 8984
rect 243544 9036 243596 9042
rect 243544 8978 243596 8984
rect 243728 8968 243780 8974
rect 243728 8910 243780 8916
rect 243176 8288 243228 8294
rect 243176 8230 243228 8236
rect 243084 8084 243136 8090
rect 243084 8026 243136 8032
rect 242900 7686 242952 7692
rect 242990 7712 243046 7721
rect 242912 6633 242940 7686
rect 242990 7647 243046 7656
rect 242898 6624 242954 6633
rect 242898 6559 242954 6568
rect 242256 5024 242308 5030
rect 242256 4966 242308 4972
rect 242624 5024 242676 5030
rect 242624 4966 242676 4972
rect 242716 5024 242768 5030
rect 242716 4966 242768 4972
rect 242268 4622 242296 4966
rect 242636 4826 242664 4966
rect 242624 4820 242676 4826
rect 242624 4762 242676 4768
rect 242256 4616 242308 4622
rect 242254 4584 242256 4593
rect 242308 4584 242310 4593
rect 242254 4519 242310 4528
rect 241612 4480 241664 4486
rect 241612 4422 241664 4428
rect 241624 4214 241652 4422
rect 241612 4208 241664 4214
rect 241612 4150 241664 4156
rect 242728 4026 242756 4966
rect 243268 4480 243320 4486
rect 243268 4422 243320 4428
rect 242898 4312 242954 4321
rect 242898 4247 242954 4256
rect 242992 4276 243044 4282
rect 242452 3998 242756 4026
rect 242452 3942 242480 3998
rect 242440 3936 242492 3942
rect 242532 3936 242584 3942
rect 242440 3878 242492 3884
rect 242530 3904 242532 3913
rect 242808 3936 242860 3942
rect 242584 3904 242586 3913
rect 242808 3878 242860 3884
rect 242530 3839 242586 3848
rect 241518 3360 241574 3369
rect 241518 3295 241574 3304
rect 240506 3224 240562 3233
rect 240506 3159 240562 3168
rect 242532 3052 242584 3058
rect 242532 2994 242584 3000
rect 241518 2680 241574 2689
rect 241518 2615 241574 2624
rect 237932 1964 237984 1970
rect 237932 1906 237984 1912
rect 240048 1964 240100 1970
rect 240048 1906 240100 1912
rect 241244 1896 241296 1902
rect 241244 1838 241296 1844
rect 239496 1828 239548 1834
rect 239496 1770 239548 1776
rect 237539 1660 237847 1669
rect 237539 1658 237545 1660
rect 237601 1658 237625 1660
rect 237681 1658 237705 1660
rect 237761 1658 237785 1660
rect 237841 1658 237847 1660
rect 237601 1606 237603 1658
rect 237783 1606 237785 1658
rect 237539 1604 237545 1606
rect 237601 1604 237625 1606
rect 237681 1604 237705 1606
rect 237761 1604 237785 1606
rect 237841 1604 237847 1606
rect 237539 1595 237847 1604
rect 239508 1494 239536 1770
rect 239496 1488 239548 1494
rect 239496 1430 239548 1436
rect 239956 1420 240008 1426
rect 239956 1362 240008 1368
rect 237380 1284 237432 1290
rect 237380 1226 237432 1232
rect 236734 1184 236790 1193
rect 236734 1119 236790 1128
rect 235724 400 235776 406
rect 229834 368 229890 377
rect 229834 303 229890 312
rect 230846 368 230902 377
rect 230846 303 230902 312
rect 233422 368 233478 377
rect 233422 303 233478 312
rect 234158 368 234214 377
rect 239968 377 239996 1362
rect 240968 1352 241020 1358
rect 240968 1294 241020 1300
rect 241060 1352 241112 1358
rect 241060 1294 241112 1300
rect 240980 377 241008 1294
rect 241072 678 241100 1294
rect 241060 672 241112 678
rect 241060 614 241112 620
rect 241256 513 241284 1838
rect 241532 1329 241560 2615
rect 242544 1834 242572 2994
rect 242820 2650 242848 3878
rect 242912 3602 242940 4247
rect 242992 4218 243044 4224
rect 242900 3596 242952 3602
rect 242900 3538 242952 3544
rect 243004 3398 243032 4218
rect 243280 4214 243308 4422
rect 243268 4208 243320 4214
rect 243268 4150 243320 4156
rect 243176 4004 243228 4010
rect 243176 3946 243228 3952
rect 242992 3392 243044 3398
rect 242992 3334 243044 3340
rect 242808 2644 242860 2650
rect 242808 2586 242860 2592
rect 243188 2038 243216 3946
rect 243740 3777 243768 8910
rect 243832 6905 243860 9454
rect 244200 8974 244228 10231
rect 244936 9586 244964 10231
rect 244924 9580 244976 9586
rect 244924 9522 244976 9528
rect 245660 9512 245712 9518
rect 245660 9454 245712 9460
rect 244188 8968 244240 8974
rect 244188 8910 244240 8916
rect 245016 8968 245068 8974
rect 245016 8910 245068 8916
rect 243818 6896 243874 6905
rect 243818 6831 243874 6840
rect 244280 6384 244332 6390
rect 244280 6326 244332 6332
rect 244188 5840 244240 5846
rect 244188 5782 244240 5788
rect 244200 4706 244228 5782
rect 244292 4826 244320 6326
rect 244280 4820 244332 4826
rect 244280 4762 244332 4768
rect 244200 4678 244320 4706
rect 244186 4176 244242 4185
rect 244186 4111 244242 4120
rect 244200 4010 244228 4111
rect 244188 4004 244240 4010
rect 244188 3946 244240 3952
rect 243726 3768 243782 3777
rect 243726 3703 243782 3712
rect 243818 2544 243874 2553
rect 243818 2479 243874 2488
rect 243452 2440 243504 2446
rect 243452 2382 243504 2388
rect 243176 2032 243228 2038
rect 243176 1974 243228 1980
rect 242900 1896 242952 1902
rect 242900 1838 242952 1844
rect 242532 1828 242584 1834
rect 242532 1770 242584 1776
rect 242912 1465 242940 1838
rect 242898 1456 242954 1465
rect 242898 1391 242954 1400
rect 241980 1352 242032 1358
rect 241518 1320 241574 1329
rect 241980 1294 242032 1300
rect 241518 1255 241574 1264
rect 241992 513 242020 1294
rect 243464 513 243492 2382
rect 243832 1902 243860 2479
rect 244292 2310 244320 4678
rect 245028 2961 245056 8910
rect 245672 6914 245700 9454
rect 246132 8974 246160 10231
rect 246120 8968 246172 8974
rect 246120 8910 246172 8916
rect 246212 8968 246264 8974
rect 246212 8910 246264 8916
rect 245580 6886 245700 6914
rect 245580 5030 245608 6886
rect 245568 5024 245620 5030
rect 245568 4966 245620 4972
rect 245384 4480 245436 4486
rect 245384 4422 245436 4428
rect 245396 4282 245424 4422
rect 245384 4276 245436 4282
rect 245384 4218 245436 4224
rect 246224 3194 246252 8910
rect 246408 8498 246436 10231
rect 246776 9450 246804 10814
rect 255688 10804 255740 10810
rect 255688 10746 255740 10752
rect 247406 10296 247462 10305
rect 247406 10231 247462 10240
rect 247866 10296 247922 10305
rect 247866 10231 247922 10240
rect 248694 10296 248750 10305
rect 248694 10231 248750 10240
rect 249338 10296 249394 10305
rect 249338 10231 249394 10240
rect 250074 10296 250130 10305
rect 250074 10231 250130 10240
rect 250810 10296 250866 10305
rect 250810 10231 250866 10240
rect 251546 10296 251602 10305
rect 251546 10231 251602 10240
rect 252282 10296 252338 10305
rect 252282 10231 252338 10240
rect 253110 10296 253166 10305
rect 253110 10231 253166 10240
rect 253846 10296 253902 10305
rect 253846 10231 253902 10240
rect 254490 10296 254546 10305
rect 254490 10231 254546 10240
rect 255226 10296 255282 10305
rect 255226 10231 255282 10240
rect 246672 9444 246724 9450
rect 246672 9386 246724 9392
rect 246764 9444 246816 9450
rect 246764 9386 246816 9392
rect 246488 8900 246540 8906
rect 246488 8842 246540 8848
rect 246396 8492 246448 8498
rect 246396 8434 246448 8440
rect 246500 4758 246528 8842
rect 246684 8498 246712 9386
rect 247420 8974 247448 10231
rect 247880 9586 247908 10231
rect 247868 9580 247920 9586
rect 247868 9522 247920 9528
rect 248708 8974 248736 10231
rect 248972 9512 249024 9518
rect 248972 9454 249024 9460
rect 247408 8968 247460 8974
rect 247408 8910 247460 8916
rect 248696 8968 248748 8974
rect 248696 8910 248748 8916
rect 247776 8900 247828 8906
rect 247776 8842 247828 8848
rect 247788 8634 247816 8842
rect 247776 8628 247828 8634
rect 247776 8570 247828 8576
rect 246672 8492 246724 8498
rect 246672 8434 246724 8440
rect 248984 7313 249012 9454
rect 249352 8498 249380 10231
rect 250088 9586 250116 10231
rect 250076 9580 250128 9586
rect 250076 9522 250128 9528
rect 250824 8974 250852 10231
rect 251456 9512 251508 9518
rect 251456 9454 251508 9460
rect 250812 8968 250864 8974
rect 250812 8910 250864 8916
rect 251364 8968 251416 8974
rect 251364 8910 251416 8916
rect 249340 8492 249392 8498
rect 249340 8434 249392 8440
rect 249616 8424 249668 8430
rect 249616 8366 249668 8372
rect 248970 7304 249026 7313
rect 248970 7239 249026 7248
rect 249628 6225 249656 8366
rect 251376 7478 251404 8910
rect 251364 7472 251416 7478
rect 251364 7414 251416 7420
rect 251468 6769 251496 9454
rect 251560 8498 251588 10231
rect 252296 8974 252324 10231
rect 253124 9586 253152 10231
rect 253112 9580 253164 9586
rect 253112 9522 253164 9528
rect 253860 8974 253888 10231
rect 254032 9512 254084 9518
rect 254032 9454 254084 9460
rect 253940 9104 253992 9110
rect 253940 9046 253992 9052
rect 252284 8968 252336 8974
rect 252284 8910 252336 8916
rect 252836 8968 252888 8974
rect 252836 8910 252888 8916
rect 253848 8968 253900 8974
rect 253848 8910 253900 8916
rect 251548 8492 251600 8498
rect 251548 8434 251600 8440
rect 251824 8424 251876 8430
rect 251824 8366 251876 8372
rect 251454 6760 251510 6769
rect 251454 6695 251510 6704
rect 249614 6216 249670 6225
rect 249614 6151 249670 6160
rect 251836 5817 251864 8366
rect 252558 6352 252614 6361
rect 252558 6287 252614 6296
rect 251822 5808 251878 5817
rect 251822 5743 251878 5752
rect 252284 5568 252336 5574
rect 252284 5510 252336 5516
rect 251456 5228 251508 5234
rect 251456 5170 251508 5176
rect 246488 4752 246540 4758
rect 246488 4694 246540 4700
rect 250626 4720 250682 4729
rect 250626 4655 250628 4664
rect 250680 4655 250682 4664
rect 250628 4626 250680 4632
rect 251468 4622 251496 5170
rect 251364 4616 251416 4622
rect 251364 4558 251416 4564
rect 251456 4616 251508 4622
rect 251456 4558 251508 4564
rect 251376 4214 251404 4558
rect 251916 4480 251968 4486
rect 251916 4422 251968 4428
rect 251364 4208 251416 4214
rect 251364 4150 251416 4156
rect 251456 4072 251508 4078
rect 251456 4014 251508 4020
rect 251468 3738 251496 4014
rect 251456 3732 251508 3738
rect 251456 3674 251508 3680
rect 251928 3534 251956 4422
rect 248972 3528 249024 3534
rect 248972 3470 249024 3476
rect 251916 3528 251968 3534
rect 251916 3470 251968 3476
rect 246212 3188 246264 3194
rect 246212 3130 246264 3136
rect 245014 2952 245070 2961
rect 245014 2887 245070 2896
rect 246488 2916 246540 2922
rect 246488 2858 246540 2864
rect 246396 2440 246448 2446
rect 246396 2382 246448 2388
rect 244280 2304 244332 2310
rect 244280 2246 244332 2252
rect 243820 1896 243872 1902
rect 243820 1838 243872 1844
rect 244280 1896 244332 1902
rect 244280 1838 244332 1844
rect 246120 1896 246172 1902
rect 246120 1838 246172 1844
rect 244292 1465 244320 1838
rect 244278 1456 244334 1465
rect 244278 1391 244334 1400
rect 243820 1352 243872 1358
rect 243820 1294 243872 1300
rect 244924 1352 244976 1358
rect 244924 1294 244976 1300
rect 243832 542 243860 1294
rect 243820 536 243872 542
rect 241242 504 241298 513
rect 241242 439 241298 448
rect 241978 504 242034 513
rect 241978 439 242034 448
rect 243450 504 243506 513
rect 244936 513 244964 1294
rect 246132 513 246160 1838
rect 246212 1352 246264 1358
rect 246212 1294 246264 1300
rect 246224 1018 246252 1294
rect 246212 1012 246264 1018
rect 246212 954 246264 960
rect 246408 513 246436 2382
rect 246500 1358 246528 2858
rect 248984 1902 249012 3470
rect 251456 3460 251508 3466
rect 251456 3402 251508 3408
rect 251468 2106 251496 3402
rect 252296 2689 252324 5510
rect 252468 5024 252520 5030
rect 252468 4966 252520 4972
rect 252480 4826 252508 4966
rect 252468 4820 252520 4826
rect 252468 4762 252520 4768
rect 252376 3392 252428 3398
rect 252376 3334 252428 3340
rect 252388 3194 252416 3334
rect 252376 3188 252428 3194
rect 252376 3130 252428 3136
rect 252282 2680 252338 2689
rect 252282 2615 252338 2624
rect 251456 2100 251508 2106
rect 251456 2042 251508 2048
rect 252572 1970 252600 6287
rect 252848 6186 252876 8910
rect 253952 8906 253980 9046
rect 253940 8900 253992 8906
rect 253940 8842 253992 8848
rect 254044 7954 254072 9454
rect 254124 9376 254176 9382
rect 254124 9318 254176 9324
rect 254136 9042 254164 9318
rect 254124 9036 254176 9042
rect 254124 8978 254176 8984
rect 254504 8498 254532 10231
rect 255240 9518 255268 10231
rect 255700 9722 255728 10746
rect 258356 10600 258408 10606
rect 258354 10568 258356 10577
rect 258408 10568 258410 10577
rect 258354 10503 258410 10512
rect 258448 10532 258500 10538
rect 258448 10474 258500 10480
rect 255872 10396 255924 10402
rect 255872 10338 255924 10344
rect 255688 9716 255740 9722
rect 255688 9658 255740 9664
rect 255884 9586 255912 10338
rect 258172 10328 258224 10334
rect 256422 10296 256478 10305
rect 256422 10231 256478 10240
rect 256698 10296 256754 10305
rect 256698 10231 256754 10240
rect 257710 10296 257766 10305
rect 258172 10270 258224 10276
rect 258262 10296 258318 10305
rect 257710 10231 257766 10240
rect 255872 9580 255924 9586
rect 255872 9522 255924 9528
rect 255228 9512 255280 9518
rect 255228 9454 255280 9460
rect 256436 9042 256464 10231
rect 256424 9036 256476 9042
rect 256424 8978 256476 8984
rect 256712 8498 256740 10231
rect 256792 9512 256844 9518
rect 256792 9454 256844 9460
rect 254492 8492 254544 8498
rect 254492 8434 254544 8440
rect 256700 8492 256752 8498
rect 256700 8434 256752 8440
rect 254768 8424 254820 8430
rect 254768 8366 254820 8372
rect 254032 7948 254084 7954
rect 254032 7890 254084 7896
rect 254780 6458 254808 8366
rect 256804 7342 256832 9454
rect 257724 9042 257752 10231
rect 257988 10056 258040 10062
rect 257988 9998 258040 10004
rect 257896 9580 257948 9586
rect 257896 9522 257948 9528
rect 257712 9036 257764 9042
rect 257712 8978 257764 8984
rect 256884 8968 256936 8974
rect 256884 8910 256936 8916
rect 257068 8968 257120 8974
rect 257068 8910 257120 8916
rect 256792 7336 256844 7342
rect 256792 7278 256844 7284
rect 254768 6452 254820 6458
rect 254768 6394 254820 6400
rect 252836 6180 252888 6186
rect 252836 6122 252888 6128
rect 256896 5710 256924 8910
rect 256884 5704 256936 5710
rect 256884 5646 256936 5652
rect 255780 5296 255832 5302
rect 255780 5238 255832 5244
rect 253572 5160 253624 5166
rect 253572 5102 253624 5108
rect 253584 4826 253612 5102
rect 255792 4826 255820 5238
rect 256884 5024 256936 5030
rect 256884 4966 256936 4972
rect 253572 4820 253624 4826
rect 253572 4762 253624 4768
rect 255780 4820 255832 4826
rect 255780 4762 255832 4768
rect 256700 4820 256752 4826
rect 256700 4762 256752 4768
rect 255320 4752 255372 4758
rect 255320 4694 255372 4700
rect 255044 4616 255096 4622
rect 255044 4558 255096 4564
rect 254032 4548 254084 4554
rect 254032 4490 254084 4496
rect 254044 4214 254072 4490
rect 255056 4321 255084 4558
rect 255332 4554 255360 4694
rect 256712 4622 256740 4762
rect 256700 4616 256752 4622
rect 256700 4558 256752 4564
rect 255320 4548 255372 4554
rect 255320 4490 255372 4496
rect 255042 4312 255098 4321
rect 255042 4247 255098 4256
rect 255332 4214 255360 4490
rect 256700 4480 256752 4486
rect 256700 4422 256752 4428
rect 254032 4208 254084 4214
rect 254032 4150 254084 4156
rect 255320 4208 255372 4214
rect 255320 4150 255372 4156
rect 256712 4078 256740 4422
rect 253940 4072 253992 4078
rect 253940 4014 253992 4020
rect 256516 4072 256568 4078
rect 256516 4014 256568 4020
rect 256700 4072 256752 4078
rect 256700 4014 256752 4020
rect 253952 3602 253980 4014
rect 256528 3738 256556 4014
rect 256516 3732 256568 3738
rect 256516 3674 256568 3680
rect 253940 3596 253992 3602
rect 253940 3538 253992 3544
rect 255320 2984 255372 2990
rect 255320 2926 255372 2932
rect 255332 2582 255360 2926
rect 255320 2576 255372 2582
rect 255320 2518 255372 2524
rect 256700 2440 256752 2446
rect 256700 2382 256752 2388
rect 255412 2304 255464 2310
rect 255412 2246 255464 2252
rect 255424 1970 255452 2246
rect 251180 1964 251232 1970
rect 251180 1906 251232 1912
rect 252560 1964 252612 1970
rect 252560 1906 252612 1912
rect 255412 1964 255464 1970
rect 255412 1906 255464 1912
rect 248420 1896 248472 1902
rect 248420 1838 248472 1844
rect 248972 1896 249024 1902
rect 248972 1838 249024 1844
rect 249800 1896 249852 1902
rect 249800 1838 249852 1844
rect 248432 1465 248460 1838
rect 249812 1465 249840 1838
rect 251192 1465 251220 1906
rect 252284 1896 252336 1902
rect 252284 1838 252336 1844
rect 253848 1896 253900 1902
rect 253848 1838 253900 1844
rect 254032 1896 254084 1902
rect 254032 1838 254084 1844
rect 255136 1896 255188 1902
rect 255136 1838 255188 1844
rect 256424 1896 256476 1902
rect 256424 1838 256476 1844
rect 248418 1456 248474 1465
rect 248418 1391 248474 1400
rect 249798 1456 249854 1465
rect 249798 1391 249854 1400
rect 251178 1456 251234 1465
rect 251178 1391 251234 1400
rect 246488 1352 246540 1358
rect 246488 1294 246540 1300
rect 248512 1352 248564 1358
rect 248512 1294 248564 1300
rect 248972 1352 249024 1358
rect 248972 1294 249024 1300
rect 251548 1352 251600 1358
rect 251548 1294 251600 1300
rect 251824 1352 251876 1358
rect 251824 1294 251876 1300
rect 248328 1284 248380 1290
rect 248328 1226 248380 1232
rect 248052 1216 248104 1222
rect 248052 1158 248104 1164
rect 248064 921 248092 1158
rect 248050 912 248106 921
rect 248050 847 248106 856
rect 248340 513 248368 1226
rect 248524 1193 248552 1294
rect 248510 1184 248566 1193
rect 248510 1119 248566 1128
rect 248984 610 249012 1294
rect 250168 1284 250220 1290
rect 250168 1226 250220 1232
rect 250180 649 250208 1226
rect 250260 1216 250312 1222
rect 250260 1158 250312 1164
rect 250272 882 250300 1158
rect 250260 876 250312 882
rect 250260 818 250312 824
rect 251560 649 251588 1294
rect 250166 640 250222 649
rect 248972 604 249024 610
rect 250166 575 250222 584
rect 251546 640 251602 649
rect 251546 575 251602 584
rect 248972 546 249024 552
rect 243820 478 243872 484
rect 244922 504 244978 513
rect 243450 439 243506 448
rect 244922 439 244978 448
rect 246118 504 246174 513
rect 246118 439 246174 448
rect 246394 504 246450 513
rect 246394 439 246450 448
rect 248326 504 248382 513
rect 248326 439 248382 448
rect 235724 342 235776 348
rect 239586 368 239642 377
rect 234158 303 234214 312
rect 239586 303 239642 312
rect 239954 368 240010 377
rect 239954 303 240010 312
rect 240966 368 241022 377
rect 251836 338 251864 1294
rect 252296 649 252324 1838
rect 253480 1352 253532 1358
rect 253480 1294 253532 1300
rect 253492 649 253520 1294
rect 253860 649 253888 1838
rect 254044 814 254072 1838
rect 254124 1352 254176 1358
rect 254124 1294 254176 1300
rect 254136 950 254164 1294
rect 254124 944 254176 950
rect 254124 886 254176 892
rect 254032 808 254084 814
rect 254032 750 254084 756
rect 252282 640 252338 649
rect 252282 575 252338 584
rect 253478 640 253534 649
rect 253478 575 253534 584
rect 253846 640 253902 649
rect 253846 575 253902 584
rect 255148 377 255176 1838
rect 255228 1352 255280 1358
rect 255228 1294 255280 1300
rect 255240 649 255268 1294
rect 256436 649 256464 1838
rect 256516 1352 256568 1358
rect 256516 1294 256568 1300
rect 255226 640 255282 649
rect 255226 575 255282 584
rect 256422 640 256478 649
rect 256422 575 256478 584
rect 256528 474 256556 1294
rect 256712 649 256740 2382
rect 256896 1970 256924 4966
rect 256976 2440 257028 2446
rect 256976 2382 257028 2388
rect 256884 1964 256936 1970
rect 256884 1906 256936 1912
rect 256988 1494 257016 2382
rect 257080 1562 257108 8910
rect 257804 4548 257856 4554
rect 257804 4490 257856 4496
rect 257712 4480 257764 4486
rect 257712 4422 257764 4428
rect 257724 4214 257752 4422
rect 257712 4208 257764 4214
rect 257712 4150 257764 4156
rect 257816 4078 257844 4490
rect 257620 4072 257672 4078
rect 257620 4014 257672 4020
rect 257804 4072 257856 4078
rect 257804 4014 257856 4020
rect 257632 3466 257660 4014
rect 257620 3460 257672 3466
rect 257620 3402 257672 3408
rect 257618 2408 257674 2417
rect 257618 2343 257674 2352
rect 257632 2106 257660 2343
rect 257908 2310 257936 9522
rect 258000 9450 258028 9998
rect 258184 9518 258212 10270
rect 258262 10231 258318 10240
rect 258356 10260 258408 10266
rect 258172 9512 258224 9518
rect 258172 9454 258224 9460
rect 257988 9444 258040 9450
rect 257988 9386 258040 9392
rect 258080 9376 258132 9382
rect 258080 9318 258132 9324
rect 258092 8498 258120 9318
rect 258172 9036 258224 9042
rect 258172 8978 258224 8984
rect 258080 8492 258132 8498
rect 258080 8434 258132 8440
rect 258184 8401 258212 8978
rect 258276 8634 258304 10231
rect 258356 10202 258408 10208
rect 258368 8974 258396 10202
rect 258460 9722 258488 10474
rect 258448 9716 258500 9722
rect 258448 9658 258500 9664
rect 258356 8968 258408 8974
rect 258356 8910 258408 8916
rect 258264 8628 258316 8634
rect 258264 8570 258316 8576
rect 258356 8492 258408 8498
rect 258356 8434 258408 8440
rect 258170 8392 258226 8401
rect 258170 8327 258226 8336
rect 258184 7818 258212 8327
rect 258368 8022 258396 8434
rect 258356 8016 258408 8022
rect 258356 7958 258408 7964
rect 258552 7954 258580 10814
rect 267740 10804 267792 10810
rect 267740 10746 267792 10752
rect 264796 10736 264848 10742
rect 264796 10678 264848 10684
rect 258724 10668 258776 10674
rect 258724 10610 258776 10616
rect 258632 10328 258684 10334
rect 258632 10270 258684 10276
rect 258644 10130 258672 10270
rect 258632 10124 258684 10130
rect 258632 10066 258684 10072
rect 258736 9994 258764 10610
rect 260196 10600 260248 10606
rect 260288 10600 260340 10606
rect 260196 10542 260248 10548
rect 260286 10568 260288 10577
rect 263140 10600 263192 10606
rect 260340 10568 260342 10577
rect 258816 10532 258868 10538
rect 258816 10474 258868 10480
rect 258724 9988 258776 9994
rect 258724 9930 258776 9936
rect 258724 9512 258776 9518
rect 258724 9454 258776 9460
rect 258736 8906 258764 9454
rect 258828 9178 258856 10474
rect 258998 10296 259054 10305
rect 258908 10260 258960 10266
rect 258998 10231 259054 10240
rect 260010 10296 260066 10305
rect 260010 10231 260066 10240
rect 258908 10202 258960 10208
rect 258816 9172 258868 9178
rect 258816 9114 258868 9120
rect 258724 8900 258776 8906
rect 258724 8842 258776 8848
rect 258540 7948 258592 7954
rect 258540 7890 258592 7896
rect 258172 7812 258224 7818
rect 258172 7754 258224 7760
rect 258632 6656 258684 6662
rect 258632 6598 258684 6604
rect 258644 6458 258672 6598
rect 258632 6452 258684 6458
rect 258632 6394 258684 6400
rect 258356 5908 258408 5914
rect 258356 5850 258408 5856
rect 258170 5128 258226 5137
rect 258170 5063 258226 5072
rect 258184 4622 258212 5063
rect 258172 4616 258224 4622
rect 258172 4558 258224 4564
rect 258184 4078 258212 4558
rect 258172 4072 258224 4078
rect 258172 4014 258224 4020
rect 258080 3936 258132 3942
rect 258080 3878 258132 3884
rect 258264 3936 258316 3942
rect 258264 3878 258316 3884
rect 258092 3534 258120 3878
rect 258276 3534 258304 3878
rect 258080 3528 258132 3534
rect 258080 3470 258132 3476
rect 258264 3528 258316 3534
rect 258264 3470 258316 3476
rect 257988 3052 258040 3058
rect 257988 2994 258040 3000
rect 257712 2304 257764 2310
rect 257712 2246 257764 2252
rect 257896 2304 257948 2310
rect 257896 2246 257948 2252
rect 257620 2100 257672 2106
rect 257620 2042 257672 2048
rect 257068 1556 257120 1562
rect 257068 1498 257120 1504
rect 256976 1488 257028 1494
rect 256976 1430 257028 1436
rect 257724 1426 257752 2246
rect 257804 2032 257856 2038
rect 257804 1974 257856 1980
rect 257712 1420 257764 1426
rect 257712 1362 257764 1368
rect 257816 1358 257844 1974
rect 257896 1964 257948 1970
rect 257896 1906 257948 1912
rect 257908 1766 257936 1906
rect 257896 1760 257948 1766
rect 257896 1702 257948 1708
rect 257804 1352 257856 1358
rect 257804 1294 257856 1300
rect 257436 1284 257488 1290
rect 257436 1226 257488 1232
rect 257448 649 257476 1226
rect 257908 785 257936 1702
rect 258000 1358 258028 2994
rect 258080 2848 258132 2854
rect 258078 2816 258080 2825
rect 258132 2816 258134 2825
rect 258078 2751 258134 2760
rect 258080 2644 258132 2650
rect 258080 2586 258132 2592
rect 258092 2378 258120 2586
rect 258080 2372 258132 2378
rect 258080 2314 258132 2320
rect 257988 1352 258040 1358
rect 257988 1294 258040 1300
rect 258092 921 258120 2314
rect 258078 912 258134 921
rect 258078 847 258134 856
rect 257894 776 257950 785
rect 258368 746 258396 5850
rect 258540 5024 258592 5030
rect 258540 4966 258592 4972
rect 258552 3942 258580 4966
rect 258540 3936 258592 3942
rect 258540 3878 258592 3884
rect 258552 3738 258580 3878
rect 258540 3732 258592 3738
rect 258540 3674 258592 3680
rect 258736 2514 258764 8842
rect 258920 8838 258948 10202
rect 258908 8832 258960 8838
rect 258908 8774 258960 8780
rect 258908 8424 258960 8430
rect 258908 8366 258960 8372
rect 258816 8288 258868 8294
rect 258816 8230 258868 8236
rect 258828 7886 258856 8230
rect 258816 7880 258868 7886
rect 258816 7822 258868 7828
rect 258816 5840 258868 5846
rect 258816 5782 258868 5788
rect 258828 5574 258856 5782
rect 258816 5568 258868 5574
rect 258816 5510 258868 5516
rect 258724 2508 258776 2514
rect 258724 2450 258776 2456
rect 258920 2106 258948 8366
rect 259012 8090 259040 10231
rect 260024 9722 260052 10231
rect 259920 9716 259972 9722
rect 259920 9658 259972 9664
rect 260012 9716 260064 9722
rect 260012 9658 260064 9664
rect 259932 9586 259960 9658
rect 259184 9580 259236 9586
rect 259184 9522 259236 9528
rect 259920 9580 259972 9586
rect 259920 9522 259972 9528
rect 259092 8900 259144 8906
rect 259092 8842 259144 8848
rect 259000 8084 259052 8090
rect 259000 8026 259052 8032
rect 259104 5642 259132 8842
rect 259196 8498 259224 9522
rect 260208 9178 260236 10542
rect 263140 10542 263192 10548
rect 260286 10503 260342 10512
rect 262218 10432 262274 10441
rect 262218 10367 262274 10376
rect 260470 10296 260526 10305
rect 260470 10231 260526 10240
rect 261758 10296 261814 10305
rect 261758 10231 261814 10240
rect 260196 9172 260248 9178
rect 260196 9114 260248 9120
rect 260104 8900 260156 8906
rect 260104 8842 260156 8848
rect 259184 8492 259236 8498
rect 259184 8434 259236 8440
rect 259644 8424 259696 8430
rect 259644 8366 259696 8372
rect 259276 5772 259328 5778
rect 259276 5714 259328 5720
rect 259092 5636 259144 5642
rect 259092 5578 259144 5584
rect 259288 4758 259316 5714
rect 259460 5024 259512 5030
rect 259460 4966 259512 4972
rect 259472 4826 259500 4966
rect 259460 4820 259512 4826
rect 259460 4762 259512 4768
rect 259276 4752 259328 4758
rect 259276 4694 259328 4700
rect 259274 3496 259330 3505
rect 259274 3431 259330 3440
rect 259000 3052 259052 3058
rect 259000 2994 259052 3000
rect 259012 2106 259040 2994
rect 259184 2848 259236 2854
rect 259184 2790 259236 2796
rect 259092 2440 259144 2446
rect 259092 2382 259144 2388
rect 258908 2100 258960 2106
rect 258908 2042 258960 2048
rect 259000 2100 259052 2106
rect 259000 2042 259052 2048
rect 258920 1970 258948 2042
rect 259104 2038 259132 2382
rect 259092 2032 259144 2038
rect 259092 1974 259144 1980
rect 258908 1964 258960 1970
rect 258908 1906 258960 1912
rect 257894 711 257950 720
rect 258356 740 258408 746
rect 258356 682 258408 688
rect 259196 649 259224 2790
rect 259288 1834 259316 3431
rect 259656 2972 259684 8366
rect 259828 8084 259880 8090
rect 259828 8026 259880 8032
rect 259736 4548 259788 4554
rect 259736 4490 259788 4496
rect 259748 3126 259776 4490
rect 259840 3210 259868 8026
rect 259920 7948 259972 7954
rect 259920 7890 259972 7896
rect 259932 7546 259960 7890
rect 259920 7540 259972 7546
rect 259920 7482 259972 7488
rect 260116 5846 260144 8842
rect 260208 8362 260236 9114
rect 260380 8968 260432 8974
rect 260380 8910 260432 8916
rect 260196 8356 260248 8362
rect 260196 8298 260248 8304
rect 260288 8288 260340 8294
rect 260288 8230 260340 8236
rect 260300 7886 260328 8230
rect 260288 7880 260340 7886
rect 260288 7822 260340 7828
rect 260392 7546 260420 8910
rect 260484 8090 260512 10231
rect 261024 9988 261076 9994
rect 261024 9930 261076 9936
rect 260656 9580 260708 9586
rect 260656 9522 260708 9528
rect 260668 9178 260696 9522
rect 260656 9172 260708 9178
rect 260656 9114 260708 9120
rect 260668 9058 260696 9114
rect 260576 9030 260696 9058
rect 260472 8084 260524 8090
rect 260472 8026 260524 8032
rect 260380 7540 260432 7546
rect 260380 7482 260432 7488
rect 260196 6656 260248 6662
rect 260196 6598 260248 6604
rect 260208 6186 260236 6598
rect 260196 6180 260248 6186
rect 260196 6122 260248 6128
rect 260104 5840 260156 5846
rect 260104 5782 260156 5788
rect 260104 4548 260156 4554
rect 260104 4490 260156 4496
rect 260012 4140 260064 4146
rect 260012 4082 260064 4088
rect 259920 3936 259972 3942
rect 259920 3878 259972 3884
rect 259932 3670 259960 3878
rect 259920 3664 259972 3670
rect 259920 3606 259972 3612
rect 260024 3466 260052 4082
rect 260116 4010 260144 4490
rect 260288 4480 260340 4486
rect 260288 4422 260340 4428
rect 260194 4312 260250 4321
rect 260194 4247 260250 4256
rect 260208 4214 260236 4247
rect 260300 4214 260328 4422
rect 260196 4208 260248 4214
rect 260196 4150 260248 4156
rect 260288 4208 260340 4214
rect 260288 4150 260340 4156
rect 260104 4004 260156 4010
rect 260104 3946 260156 3952
rect 260012 3460 260064 3466
rect 260012 3402 260064 3408
rect 259840 3182 259960 3210
rect 259932 3126 259960 3182
rect 259736 3120 259788 3126
rect 259736 3062 259788 3068
rect 259920 3120 259972 3126
rect 259920 3062 259972 3068
rect 259656 2944 259868 2972
rect 259840 1970 259868 2944
rect 260576 2774 260604 9030
rect 260656 8900 260708 8906
rect 260656 8842 260708 8848
rect 260668 5273 260696 8842
rect 260932 8560 260984 8566
rect 260932 8502 260984 8508
rect 260840 8424 260892 8430
rect 260840 8366 260892 8372
rect 260852 7818 260880 8366
rect 260840 7812 260892 7818
rect 260840 7754 260892 7760
rect 260944 7750 260972 8502
rect 260932 7744 260984 7750
rect 260932 7686 260984 7692
rect 261036 6798 261064 9930
rect 261208 9580 261260 9586
rect 261208 9522 261260 9528
rect 261116 8492 261168 8498
rect 261116 8434 261168 8440
rect 261024 6792 261076 6798
rect 261024 6734 261076 6740
rect 261128 5914 261156 8434
rect 261220 8362 261248 9522
rect 261484 9512 261536 9518
rect 261484 9454 261536 9460
rect 261496 9382 261524 9454
rect 261484 9376 261536 9382
rect 261484 9318 261536 9324
rect 261576 9376 261628 9382
rect 261576 9318 261628 9324
rect 261496 8498 261524 9318
rect 261484 8492 261536 8498
rect 261404 8452 261484 8480
rect 261208 8356 261260 8362
rect 261208 8298 261260 8304
rect 261208 6316 261260 6322
rect 261208 6258 261260 6264
rect 261220 5914 261248 6258
rect 261116 5908 261168 5914
rect 261116 5850 261168 5856
rect 261208 5908 261260 5914
rect 261208 5850 261260 5856
rect 261128 5642 261156 5850
rect 261116 5636 261168 5642
rect 261116 5578 261168 5584
rect 260654 5264 260710 5273
rect 260654 5199 260710 5208
rect 260668 5166 260696 5199
rect 260656 5160 260708 5166
rect 260656 5102 260708 5108
rect 260840 3528 260892 3534
rect 260838 3496 260840 3505
rect 260892 3496 260894 3505
rect 260838 3431 260894 3440
rect 260300 2746 260604 2774
rect 261404 2774 261432 8452
rect 261484 8434 261536 8440
rect 261588 7410 261616 9318
rect 261772 7546 261800 10231
rect 262232 9722 262260 10367
rect 262494 10296 262550 10305
rect 262494 10231 262550 10240
rect 262404 10124 262456 10130
rect 262404 10066 262456 10072
rect 262128 9716 262180 9722
rect 262128 9658 262180 9664
rect 262220 9716 262272 9722
rect 262220 9658 262272 9664
rect 262140 9518 262168 9658
rect 262128 9512 262180 9518
rect 262128 9454 262180 9460
rect 262036 9376 262088 9382
rect 262036 9318 262088 9324
rect 262048 9110 262076 9318
rect 262036 9104 262088 9110
rect 262036 9046 262088 9052
rect 261852 8832 261904 8838
rect 261852 8774 261904 8780
rect 261864 7886 261892 8774
rect 261944 8356 261996 8362
rect 261944 8298 261996 8304
rect 261956 7886 261984 8298
rect 262310 8256 262366 8265
rect 262310 8191 262366 8200
rect 261852 7880 261904 7886
rect 261852 7822 261904 7828
rect 261944 7880 261996 7886
rect 262324 7834 262352 8191
rect 261944 7822 261996 7828
rect 261760 7540 261812 7546
rect 261760 7482 261812 7488
rect 261576 7404 261628 7410
rect 261576 7346 261628 7352
rect 261864 7018 261892 7822
rect 262232 7806 262352 7834
rect 261864 6990 262076 7018
rect 262048 6610 262076 6990
rect 262232 6746 262260 7806
rect 262312 7744 262364 7750
rect 262312 7686 262364 7692
rect 262324 7410 262352 7686
rect 262312 7404 262364 7410
rect 262312 7346 262364 7352
rect 262416 7256 262444 10066
rect 262508 7546 262536 10231
rect 262864 10192 262916 10198
rect 262864 10134 262916 10140
rect 262876 9722 262904 10134
rect 263152 9722 263180 10542
rect 263600 10464 263652 10470
rect 263600 10406 263652 10412
rect 264426 10432 264482 10441
rect 263230 10296 263286 10305
rect 263230 10231 263286 10240
rect 262864 9716 262916 9722
rect 262864 9658 262916 9664
rect 263140 9716 263192 9722
rect 263140 9658 263192 9664
rect 262876 9586 262904 9658
rect 262864 9580 262916 9586
rect 262864 9522 262916 9528
rect 262588 8900 262640 8906
rect 262588 8842 262640 8848
rect 262600 8809 262628 8842
rect 262586 8800 262642 8809
rect 262586 8735 262642 8744
rect 262588 8628 262640 8634
rect 262588 8570 262640 8576
rect 262600 7886 262628 8570
rect 262876 8401 262904 9522
rect 262956 9172 263008 9178
rect 262956 9114 263008 9120
rect 262862 8392 262918 8401
rect 262862 8327 262918 8336
rect 262680 8288 262732 8294
rect 262680 8230 262732 8236
rect 262588 7880 262640 7886
rect 262588 7822 262640 7828
rect 262496 7540 262548 7546
rect 262496 7482 262548 7488
rect 262140 6730 262260 6746
rect 262128 6724 262260 6730
rect 262180 6718 262260 6724
rect 262324 7228 262444 7256
rect 262128 6666 262180 6672
rect 262048 6582 262260 6610
rect 261484 6248 261536 6254
rect 261482 6216 261484 6225
rect 261536 6216 261538 6225
rect 261482 6151 261538 6160
rect 261668 6112 261720 6118
rect 261668 6054 261720 6060
rect 261680 5710 261708 6054
rect 262232 5930 262260 6582
rect 262140 5902 262260 5930
rect 261668 5704 261720 5710
rect 261668 5646 261720 5652
rect 261944 5568 261996 5574
rect 261944 5510 261996 5516
rect 261956 5302 261984 5510
rect 261944 5296 261996 5302
rect 261944 5238 261996 5244
rect 262140 5250 262168 5902
rect 262324 5817 262352 7228
rect 262494 7168 262550 7177
rect 262494 7103 262550 7112
rect 262508 6798 262536 7103
rect 262496 6792 262548 6798
rect 262496 6734 262548 6740
rect 262404 6316 262456 6322
rect 262404 6258 262456 6264
rect 262496 6316 262548 6322
rect 262496 6258 262548 6264
rect 262310 5808 262366 5817
rect 262220 5772 262272 5778
rect 262310 5743 262366 5752
rect 262220 5714 262272 5720
rect 262232 5370 262260 5714
rect 262220 5364 262272 5370
rect 262220 5306 262272 5312
rect 262140 5222 262352 5250
rect 262220 3188 262272 3194
rect 262220 3130 262272 3136
rect 262232 3097 262260 3130
rect 262218 3088 262274 3097
rect 262218 3023 262274 3032
rect 261404 2746 261524 2774
rect 259920 2304 259972 2310
rect 259920 2246 259972 2252
rect 259828 1964 259880 1970
rect 259828 1906 259880 1912
rect 259276 1828 259328 1834
rect 259276 1770 259328 1776
rect 259932 649 259960 2246
rect 260104 2032 260156 2038
rect 260104 1974 260156 1980
rect 260116 1766 260144 1974
rect 260300 1970 260328 2746
rect 261496 1970 261524 2746
rect 261576 2440 261628 2446
rect 261576 2382 261628 2388
rect 261588 2106 261616 2382
rect 261852 2304 261904 2310
rect 261852 2246 261904 2252
rect 261576 2100 261628 2106
rect 261576 2042 261628 2048
rect 260288 1964 260340 1970
rect 260288 1906 260340 1912
rect 261484 1964 261536 1970
rect 261484 1906 261536 1912
rect 260104 1760 260156 1766
rect 260104 1702 260156 1708
rect 260288 1760 260340 1766
rect 260288 1702 260340 1708
rect 261576 1760 261628 1766
rect 261576 1702 261628 1708
rect 260300 1358 260328 1702
rect 261588 1358 261616 1702
rect 260288 1352 260340 1358
rect 260288 1294 260340 1300
rect 261576 1352 261628 1358
rect 261576 1294 261628 1300
rect 260472 1216 260524 1222
rect 260472 1158 260524 1164
rect 261760 1216 261812 1222
rect 261760 1158 261812 1164
rect 260484 649 260512 1158
rect 261772 649 261800 1158
rect 256698 640 256754 649
rect 256698 575 256754 584
rect 257434 640 257490 649
rect 257434 575 257490 584
rect 259182 640 259238 649
rect 259182 575 259238 584
rect 259918 640 259974 649
rect 259918 575 259974 584
rect 260470 640 260526 649
rect 260470 575 260526 584
rect 261758 640 261814 649
rect 261758 575 261814 584
rect 261864 513 261892 2246
rect 262324 1970 262352 5222
rect 262416 2990 262444 6258
rect 262508 5234 262536 6258
rect 262496 5228 262548 5234
rect 262496 5170 262548 5176
rect 262404 2984 262456 2990
rect 262404 2926 262456 2932
rect 262600 1970 262628 7822
rect 262692 7206 262720 8230
rect 262680 7200 262732 7206
rect 262680 7142 262732 7148
rect 262680 6928 262732 6934
rect 262680 6870 262732 6876
rect 262692 5846 262720 6870
rect 262968 6458 262996 9114
rect 263152 7886 263180 9658
rect 263140 7880 263192 7886
rect 263140 7822 263192 7828
rect 263048 7744 263100 7750
rect 263048 7686 263100 7692
rect 263060 7410 263088 7686
rect 263048 7404 263100 7410
rect 263048 7346 263100 7352
rect 262956 6452 263008 6458
rect 262956 6394 263008 6400
rect 263046 5944 263102 5953
rect 263152 5930 263180 7822
rect 263244 7546 263272 10231
rect 263324 10124 263376 10130
rect 263324 10066 263376 10072
rect 263232 7540 263284 7546
rect 263232 7482 263284 7488
rect 263152 5902 263272 5930
rect 263046 5879 263102 5888
rect 262680 5840 262732 5846
rect 262680 5782 262732 5788
rect 262954 5808 263010 5817
rect 262954 5743 263010 5752
rect 262968 5234 262996 5743
rect 262956 5228 263008 5234
rect 262956 5170 263008 5176
rect 263060 4826 263088 5879
rect 263140 5772 263192 5778
rect 263140 5714 263192 5720
rect 263152 5681 263180 5714
rect 263138 5672 263194 5681
rect 263138 5607 263140 5616
rect 263192 5607 263194 5616
rect 263140 5578 263192 5584
rect 263244 5386 263272 5902
rect 263152 5358 263272 5386
rect 263048 4820 263100 4826
rect 263048 4762 263100 4768
rect 263152 4434 263180 5358
rect 263230 5264 263286 5273
rect 263230 5199 263286 5208
rect 263244 5166 263272 5199
rect 263232 5160 263284 5166
rect 263232 5102 263284 5108
rect 263336 4622 263364 10066
rect 263612 8634 263640 10406
rect 264426 10367 264482 10376
rect 264334 10296 264390 10305
rect 264334 10231 264390 10240
rect 263968 9920 264020 9926
rect 263968 9862 264020 9868
rect 263980 9586 264008 9862
rect 263968 9580 264020 9586
rect 263968 9522 264020 9528
rect 263692 9444 263744 9450
rect 263692 9386 263744 9392
rect 263600 8628 263652 8634
rect 263600 8570 263652 8576
rect 263600 8492 263652 8498
rect 263600 8434 263652 8440
rect 263508 6792 263560 6798
rect 263508 6734 263560 6740
rect 263416 6656 263468 6662
rect 263414 6624 263416 6633
rect 263468 6624 263470 6633
rect 263414 6559 263470 6568
rect 263414 6488 263470 6497
rect 263520 6458 263548 6734
rect 263414 6423 263416 6432
rect 263468 6423 263470 6432
rect 263508 6452 263560 6458
rect 263416 6394 263468 6400
rect 263508 6394 263560 6400
rect 263612 5642 263640 8434
rect 263704 6934 263732 9386
rect 263784 9376 263836 9382
rect 263784 9318 263836 9324
rect 263796 8974 263824 9318
rect 263876 9104 263928 9110
rect 263876 9046 263928 9052
rect 263784 8968 263836 8974
rect 263784 8910 263836 8916
rect 263784 7880 263836 7886
rect 263784 7822 263836 7828
rect 263796 7585 263824 7822
rect 263782 7576 263838 7585
rect 263782 7511 263838 7520
rect 263888 7274 263916 9046
rect 263980 8362 264008 9522
rect 264060 9376 264112 9382
rect 264060 9318 264112 9324
rect 263968 8356 264020 8362
rect 263968 8298 264020 8304
rect 263876 7268 263928 7274
rect 263876 7210 263928 7216
rect 263692 6928 263744 6934
rect 263692 6870 263744 6876
rect 263600 5636 263652 5642
rect 263600 5578 263652 5584
rect 263324 4616 263376 4622
rect 263324 4558 263376 4564
rect 263152 4406 263456 4434
rect 262312 1964 262364 1970
rect 262312 1906 262364 1912
rect 262588 1964 262640 1970
rect 262588 1906 262640 1912
rect 263428 1902 263456 4406
rect 263980 2446 264008 8298
rect 264072 6798 264100 9318
rect 264244 8628 264296 8634
rect 264244 8570 264296 8576
rect 264256 8498 264284 8570
rect 264244 8492 264296 8498
rect 264244 8434 264296 8440
rect 264244 8288 264296 8294
rect 264244 8230 264296 8236
rect 264256 7954 264284 8230
rect 264244 7948 264296 7954
rect 264244 7890 264296 7896
rect 264152 7744 264204 7750
rect 264152 7686 264204 7692
rect 264244 7744 264296 7750
rect 264244 7686 264296 7692
rect 264164 7410 264192 7686
rect 264256 7410 264284 7686
rect 264348 7546 264376 10231
rect 264336 7540 264388 7546
rect 264336 7482 264388 7488
rect 264152 7404 264204 7410
rect 264152 7346 264204 7352
rect 264244 7404 264296 7410
rect 264244 7346 264296 7352
rect 264256 6798 264284 7346
rect 264060 6792 264112 6798
rect 264244 6792 264296 6798
rect 264060 6734 264112 6740
rect 264150 6760 264206 6769
rect 264244 6734 264296 6740
rect 264150 6695 264206 6704
rect 264164 6662 264192 6695
rect 264440 6662 264468 10367
rect 264704 9648 264756 9654
rect 264704 9590 264756 9596
rect 264716 9110 264744 9590
rect 264808 9110 264836 10678
rect 266820 10668 266872 10674
rect 266820 10610 266872 10616
rect 266636 10328 266688 10334
rect 265714 10296 265770 10305
rect 266636 10270 266688 10276
rect 265714 10231 265770 10240
rect 264980 9920 265032 9926
rect 264980 9862 265032 9868
rect 264704 9104 264756 9110
rect 264704 9046 264756 9052
rect 264796 9104 264848 9110
rect 264796 9046 264848 9052
rect 264808 8838 264836 9046
rect 264796 8832 264848 8838
rect 264796 8774 264848 8780
rect 264808 8650 264836 8774
rect 264624 8622 264836 8650
rect 264888 8628 264940 8634
rect 264520 8492 264572 8498
rect 264520 8434 264572 8440
rect 264152 6656 264204 6662
rect 264152 6598 264204 6604
rect 264428 6656 264480 6662
rect 264428 6598 264480 6604
rect 264244 6316 264296 6322
rect 264244 6258 264296 6264
rect 264060 5704 264112 5710
rect 264060 5646 264112 5652
rect 264072 5409 264100 5646
rect 264058 5400 264114 5409
rect 264058 5335 264114 5344
rect 264256 4758 264284 6258
rect 264532 5710 264560 8434
rect 264624 6322 264652 8622
rect 264888 8570 264940 8576
rect 264900 7290 264928 8570
rect 264808 7262 264928 7290
rect 264704 6656 264756 6662
rect 264704 6598 264756 6604
rect 264716 6390 264744 6598
rect 264704 6384 264756 6390
rect 264704 6326 264756 6332
rect 264612 6316 264664 6322
rect 264612 6258 264664 6264
rect 264520 5704 264572 5710
rect 264520 5646 264572 5652
rect 264716 5234 264744 6326
rect 264704 5228 264756 5234
rect 264704 5170 264756 5176
rect 264428 5092 264480 5098
rect 264428 5034 264480 5040
rect 264060 4752 264112 4758
rect 264060 4694 264112 4700
rect 264244 4752 264296 4758
rect 264244 4694 264296 4700
rect 264072 3194 264100 4694
rect 264152 4548 264204 4554
rect 264152 4490 264204 4496
rect 264060 3188 264112 3194
rect 264060 3130 264112 3136
rect 263968 2440 264020 2446
rect 263968 2382 264020 2388
rect 264164 2038 264192 4490
rect 264244 2440 264296 2446
rect 264244 2382 264296 2388
rect 264152 2032 264204 2038
rect 264152 1974 264204 1980
rect 264256 1970 264284 2382
rect 264440 2378 264468 5034
rect 264808 3942 264836 7262
rect 264888 7200 264940 7206
rect 264888 7142 264940 7148
rect 264900 5642 264928 7142
rect 264888 5636 264940 5642
rect 264888 5578 264940 5584
rect 264886 4584 264942 4593
rect 264886 4519 264942 4528
rect 264900 4282 264928 4519
rect 264888 4276 264940 4282
rect 264888 4218 264940 4224
rect 264992 4214 265020 9862
rect 265072 9580 265124 9586
rect 265072 9522 265124 9528
rect 265084 9042 265112 9522
rect 265348 9512 265400 9518
rect 265348 9454 265400 9460
rect 265072 9036 265124 9042
rect 265072 8978 265124 8984
rect 265164 9036 265216 9042
rect 265164 8978 265216 8984
rect 265176 8906 265204 8978
rect 265164 8900 265216 8906
rect 265164 8842 265216 8848
rect 265360 8838 265388 9454
rect 265532 9376 265584 9382
rect 265532 9318 265584 9324
rect 265624 9376 265676 9382
rect 265624 9318 265676 9324
rect 265348 8832 265400 8838
rect 265348 8774 265400 8780
rect 265164 8492 265216 8498
rect 265164 8434 265216 8440
rect 265072 7744 265124 7750
rect 265072 7686 265124 7692
rect 265084 7002 265112 7686
rect 265072 6996 265124 7002
rect 265072 6938 265124 6944
rect 265176 6254 265204 8434
rect 265256 7880 265308 7886
rect 265256 7822 265308 7828
rect 265268 7410 265296 7822
rect 265256 7404 265308 7410
rect 265256 7346 265308 7352
rect 265360 7290 265388 8774
rect 265440 7744 265492 7750
rect 265440 7686 265492 7692
rect 265268 7262 265388 7290
rect 265164 6248 265216 6254
rect 265164 6190 265216 6196
rect 265268 6100 265296 7262
rect 265346 6896 265402 6905
rect 265346 6831 265402 6840
rect 265084 6072 265296 6100
rect 264980 4208 265032 4214
rect 264980 4150 265032 4156
rect 264796 3936 264848 3942
rect 264796 3878 264848 3884
rect 264428 2372 264480 2378
rect 264428 2314 264480 2320
rect 264980 2304 265032 2310
rect 264980 2246 265032 2252
rect 264244 1964 264296 1970
rect 264244 1906 264296 1912
rect 263416 1896 263468 1902
rect 263416 1838 263468 1844
rect 262312 1760 262364 1766
rect 262312 1702 262364 1708
rect 263048 1760 263100 1766
rect 263048 1702 263100 1708
rect 264152 1760 264204 1766
rect 264152 1702 264204 1708
rect 262324 1358 262352 1702
rect 263060 1358 263088 1702
rect 264164 1358 264192 1702
rect 264992 1465 265020 2246
rect 265084 1902 265112 6072
rect 265256 5704 265308 5710
rect 265256 5646 265308 5652
rect 265164 5160 265216 5166
rect 265164 5102 265216 5108
rect 265176 4826 265204 5102
rect 265164 4820 265216 4826
rect 265164 4762 265216 4768
rect 265268 2825 265296 5646
rect 265360 3738 265388 6831
rect 265348 3732 265400 3738
rect 265348 3674 265400 3680
rect 265452 3641 265480 7686
rect 265544 6798 265572 9318
rect 265532 6792 265584 6798
rect 265532 6734 265584 6740
rect 265636 6458 265664 9318
rect 265728 6662 265756 10231
rect 265900 10056 265952 10062
rect 265900 9998 265952 10004
rect 266268 10056 266320 10062
rect 266268 9998 266320 10004
rect 265912 9518 265940 9998
rect 265992 9580 266044 9586
rect 265992 9522 266044 9528
rect 265900 9512 265952 9518
rect 265900 9454 265952 9460
rect 265808 8968 265860 8974
rect 265808 8910 265860 8916
rect 265820 8430 265848 8910
rect 265912 8498 265940 9454
rect 266004 8974 266032 9522
rect 265992 8968 266044 8974
rect 265992 8910 266044 8916
rect 265900 8492 265952 8498
rect 265900 8434 265952 8440
rect 265808 8424 265860 8430
rect 265808 8366 265860 8372
rect 265820 7886 265848 8366
rect 265808 7880 265860 7886
rect 265808 7822 265860 7828
rect 265806 7712 265862 7721
rect 265806 7647 265862 7656
rect 265820 7342 265848 7647
rect 265808 7336 265860 7342
rect 265808 7278 265860 7284
rect 265716 6656 265768 6662
rect 265716 6598 265768 6604
rect 265808 6656 265860 6662
rect 265808 6598 265860 6604
rect 265624 6452 265676 6458
rect 265624 6394 265676 6400
rect 265820 6322 265848 6598
rect 265808 6316 265860 6322
rect 265808 6258 265860 6264
rect 265912 6202 265940 8434
rect 265992 7880 266044 7886
rect 265992 7822 266044 7828
rect 266004 7585 266032 7822
rect 266176 7812 266228 7818
rect 266176 7754 266228 7760
rect 266084 7744 266136 7750
rect 266084 7686 266136 7692
rect 265990 7576 266046 7585
rect 265990 7511 266046 7520
rect 265728 6174 265940 6202
rect 265728 4162 265756 6174
rect 265900 5636 265952 5642
rect 265900 5578 265952 5584
rect 265912 4622 265940 5578
rect 265992 5228 266044 5234
rect 265992 5170 266044 5176
rect 265808 4616 265860 4622
rect 265808 4558 265860 4564
rect 265900 4616 265952 4622
rect 265900 4558 265952 4564
rect 265820 4282 265848 4558
rect 265808 4276 265860 4282
rect 265808 4218 265860 4224
rect 265728 4134 265848 4162
rect 265624 4072 265676 4078
rect 265624 4014 265676 4020
rect 265438 3632 265494 3641
rect 265438 3567 265494 3576
rect 265636 3398 265664 4014
rect 265624 3392 265676 3398
rect 265624 3334 265676 3340
rect 265532 2848 265584 2854
rect 265254 2816 265310 2825
rect 265532 2790 265584 2796
rect 265254 2751 265310 2760
rect 265072 1896 265124 1902
rect 265072 1838 265124 1844
rect 265164 1760 265216 1766
rect 265164 1702 265216 1708
rect 264978 1456 265034 1465
rect 264978 1391 265034 1400
rect 265176 1358 265204 1702
rect 262312 1352 262364 1358
rect 262312 1294 262364 1300
rect 263048 1352 263100 1358
rect 263048 1294 263100 1300
rect 264152 1352 264204 1358
rect 264152 1294 264204 1300
rect 265164 1352 265216 1358
rect 265164 1294 265216 1300
rect 262496 1216 262548 1222
rect 262496 1158 262548 1164
rect 263232 1216 263284 1222
rect 263232 1158 263284 1164
rect 264336 1216 264388 1222
rect 264336 1158 264388 1164
rect 265348 1216 265400 1222
rect 265348 1158 265400 1164
rect 262508 649 262536 1158
rect 263244 649 263272 1158
rect 264348 649 264376 1158
rect 265360 649 265388 1158
rect 265544 1018 265572 2790
rect 265820 1902 265848 4134
rect 265900 4140 265952 4146
rect 265900 4082 265952 4088
rect 265912 3233 265940 4082
rect 266004 3738 266032 5170
rect 266096 4622 266124 7686
rect 266188 7585 266216 7754
rect 266174 7576 266230 7585
rect 266174 7511 266230 7520
rect 266188 6934 266216 7511
rect 266176 6928 266228 6934
rect 266176 6870 266228 6876
rect 266176 6452 266228 6458
rect 266176 6394 266228 6400
rect 266188 5642 266216 6394
rect 266176 5636 266228 5642
rect 266176 5578 266228 5584
rect 266188 5234 266216 5578
rect 266176 5228 266228 5234
rect 266176 5170 266228 5176
rect 266280 5114 266308 9998
rect 266648 8838 266676 10270
rect 266728 9512 266780 9518
rect 266728 9454 266780 9460
rect 266636 8832 266688 8838
rect 266636 8774 266688 8780
rect 266452 8492 266504 8498
rect 266452 8434 266504 8440
rect 266464 8401 266492 8434
rect 266450 8392 266506 8401
rect 266450 8327 266506 8336
rect 266648 7342 266676 8774
rect 266636 7336 266688 7342
rect 266636 7278 266688 7284
rect 266360 5568 266412 5574
rect 266360 5510 266412 5516
rect 266188 5086 266308 5114
rect 266084 4616 266136 4622
rect 266084 4558 266136 4564
rect 266188 4434 266216 5086
rect 266268 4684 266320 4690
rect 266268 4626 266320 4632
rect 266096 4406 266216 4434
rect 265992 3732 266044 3738
rect 265992 3674 266044 3680
rect 266096 3534 266124 4406
rect 266176 4276 266228 4282
rect 266176 4218 266228 4224
rect 266188 3534 266216 4218
rect 266084 3528 266136 3534
rect 266084 3470 266136 3476
rect 266176 3528 266228 3534
rect 266176 3470 266228 3476
rect 265898 3224 265954 3233
rect 265898 3159 265954 3168
rect 266280 3058 266308 4626
rect 266372 3942 266400 5510
rect 266648 5250 266676 7278
rect 266740 6118 266768 9454
rect 266832 8906 266860 10610
rect 267004 10260 267056 10266
rect 267004 10202 267056 10208
rect 267016 9382 267044 10202
rect 267648 9512 267700 9518
rect 267646 9480 267648 9489
rect 267700 9480 267702 9489
rect 267646 9415 267702 9424
rect 267004 9376 267056 9382
rect 267004 9318 267056 9324
rect 266820 8900 266872 8906
rect 266820 8842 266872 8848
rect 266912 8560 266964 8566
rect 266912 8502 266964 8508
rect 266924 6254 266952 8502
rect 267016 7342 267044 9318
rect 267556 9104 267608 9110
rect 267556 9046 267608 9052
rect 267464 8968 267516 8974
rect 267464 8910 267516 8916
rect 267188 8900 267240 8906
rect 267188 8842 267240 8848
rect 267372 8900 267424 8906
rect 267372 8842 267424 8848
rect 267096 8492 267148 8498
rect 267096 8434 267148 8440
rect 267004 7336 267056 7342
rect 267004 7278 267056 7284
rect 267108 6905 267136 8434
rect 267094 6896 267150 6905
rect 267094 6831 267150 6840
rect 267004 6792 267056 6798
rect 267004 6734 267056 6740
rect 266912 6248 266964 6254
rect 266912 6190 266964 6196
rect 266728 6112 266780 6118
rect 266728 6054 266780 6060
rect 266728 5772 266780 5778
rect 266728 5714 266780 5720
rect 266740 5370 266768 5714
rect 266910 5672 266966 5681
rect 266910 5607 266966 5616
rect 266728 5364 266780 5370
rect 266728 5306 266780 5312
rect 266648 5222 266768 5250
rect 266636 5092 266688 5098
rect 266636 5034 266688 5040
rect 266450 4312 266506 4321
rect 266450 4247 266506 4256
rect 266360 3936 266412 3942
rect 266360 3878 266412 3884
rect 266268 3052 266320 3058
rect 266268 2994 266320 3000
rect 266464 2650 266492 4247
rect 266648 2854 266676 5034
rect 266636 2848 266688 2854
rect 266636 2790 266688 2796
rect 266634 2680 266690 2689
rect 266452 2644 266504 2650
rect 266634 2615 266690 2624
rect 266452 2586 266504 2592
rect 266648 1902 266676 2615
rect 266740 1902 266768 5222
rect 266820 5024 266872 5030
rect 266820 4966 266872 4972
rect 266832 3058 266860 4966
rect 266924 4826 266952 5607
rect 266912 4820 266964 4826
rect 266912 4762 266964 4768
rect 267016 4010 267044 6734
rect 267096 6112 267148 6118
rect 267096 6054 267148 6060
rect 267108 4146 267136 6054
rect 267200 5710 267228 8842
rect 267278 7848 267334 7857
rect 267278 7783 267280 7792
rect 267332 7783 267334 7792
rect 267280 7754 267332 7760
rect 267384 7410 267412 8842
rect 267476 8634 267504 8910
rect 267464 8628 267516 8634
rect 267464 8570 267516 8576
rect 267464 8288 267516 8294
rect 267464 8230 267516 8236
rect 267476 7886 267504 8230
rect 267464 7880 267516 7886
rect 267464 7822 267516 7828
rect 267464 7744 267516 7750
rect 267464 7686 267516 7692
rect 267372 7404 267424 7410
rect 267372 7346 267424 7352
rect 267280 7336 267332 7342
rect 267476 7290 267504 7686
rect 267280 7278 267332 7284
rect 267292 6225 267320 7278
rect 267384 7262 267504 7290
rect 267278 6216 267334 6225
rect 267278 6151 267334 6160
rect 267188 5704 267240 5710
rect 267188 5646 267240 5652
rect 267186 5536 267242 5545
rect 267186 5471 267242 5480
rect 267200 4146 267228 5471
rect 267278 5400 267334 5409
rect 267278 5335 267334 5344
rect 267292 5302 267320 5335
rect 267280 5296 267332 5302
rect 267280 5238 267332 5244
rect 267384 4622 267412 7262
rect 267464 7200 267516 7206
rect 267464 7142 267516 7148
rect 267476 5234 267504 7142
rect 267464 5228 267516 5234
rect 267464 5170 267516 5176
rect 267464 5092 267516 5098
rect 267464 5034 267516 5040
rect 267372 4616 267424 4622
rect 267372 4558 267424 4564
rect 267278 4448 267334 4457
rect 267278 4383 267334 4392
rect 267096 4140 267148 4146
rect 267096 4082 267148 4088
rect 267188 4140 267240 4146
rect 267188 4082 267240 4088
rect 267004 4004 267056 4010
rect 267004 3946 267056 3952
rect 266820 3052 266872 3058
rect 266820 2994 266872 3000
rect 266818 2952 266874 2961
rect 266818 2887 266874 2896
rect 267188 2916 267240 2922
rect 266832 2854 266860 2887
rect 267188 2858 267240 2864
rect 266820 2848 266872 2854
rect 266820 2790 266872 2796
rect 267200 2689 267228 2858
rect 267186 2680 267242 2689
rect 267186 2615 267242 2624
rect 267292 2448 267320 4383
rect 267370 3768 267426 3777
rect 267370 3703 267426 3712
rect 267384 3534 267412 3703
rect 267372 3528 267424 3534
rect 267372 3470 267424 3476
rect 267476 3058 267504 5034
rect 267568 4622 267596 9046
rect 267752 8838 267780 10746
rect 267844 9586 267872 10814
rect 268200 10532 268252 10538
rect 268200 10474 268252 10480
rect 268016 10396 268068 10402
rect 268016 10338 268068 10344
rect 267924 9988 267976 9994
rect 267924 9930 267976 9936
rect 267832 9580 267884 9586
rect 267832 9522 267884 9528
rect 267936 8945 267964 9930
rect 268028 9217 268056 10338
rect 268108 9648 268160 9654
rect 268108 9590 268160 9596
rect 268014 9208 268070 9217
rect 268014 9143 268070 9152
rect 268120 9081 268148 9590
rect 268212 9382 268240 10474
rect 270408 10192 270460 10198
rect 270408 10134 270460 10140
rect 268936 10124 268988 10130
rect 268936 10066 268988 10072
rect 268476 9920 268528 9926
rect 268476 9862 268528 9868
rect 268488 9625 268516 9862
rect 268474 9616 268530 9625
rect 268474 9551 268530 9560
rect 268844 9580 268896 9586
rect 268844 9522 268896 9528
rect 268476 9512 268528 9518
rect 268476 9454 268528 9460
rect 268660 9512 268712 9518
rect 268660 9454 268712 9460
rect 268200 9376 268252 9382
rect 268200 9318 268252 9324
rect 268106 9072 268162 9081
rect 268106 9007 268162 9016
rect 268292 8968 268344 8974
rect 267922 8936 267978 8945
rect 268292 8910 268344 8916
rect 267922 8871 267978 8880
rect 267740 8832 267792 8838
rect 267740 8774 267792 8780
rect 267648 8628 267700 8634
rect 267648 8570 267700 8576
rect 267660 8498 267688 8570
rect 267752 8498 267780 8774
rect 268304 8634 268332 8910
rect 268292 8628 268344 8634
rect 268292 8570 268344 8576
rect 268120 8498 268424 8514
rect 267648 8492 267700 8498
rect 267648 8434 267700 8440
rect 267740 8492 267792 8498
rect 267740 8434 267792 8440
rect 268016 8492 268068 8498
rect 268016 8434 268068 8440
rect 268120 8492 268436 8498
rect 268120 8486 268384 8492
rect 268028 8242 268056 8434
rect 268120 8430 268148 8486
rect 268384 8434 268436 8440
rect 268108 8424 268160 8430
rect 268108 8366 268160 8372
rect 268028 8214 268148 8242
rect 268120 8090 268148 8214
rect 268016 8084 268068 8090
rect 268016 8026 268068 8032
rect 268108 8084 268160 8090
rect 268108 8026 268160 8032
rect 268028 7857 268056 8026
rect 268292 7880 268344 7886
rect 267830 7848 267886 7857
rect 267648 7812 267700 7818
rect 267830 7783 267886 7792
rect 268014 7848 268070 7857
rect 268292 7822 268344 7828
rect 268014 7783 268070 7792
rect 267648 7754 267700 7760
rect 267660 7721 267688 7754
rect 267646 7712 267702 7721
rect 267646 7647 267702 7656
rect 267646 7576 267702 7585
rect 267646 7511 267702 7520
rect 267660 7410 267688 7511
rect 267648 7404 267700 7410
rect 267648 7346 267700 7352
rect 267738 7304 267794 7313
rect 267738 7239 267740 7248
rect 267792 7239 267794 7248
rect 267740 7210 267792 7216
rect 267648 7200 267700 7206
rect 267648 7142 267700 7148
rect 267556 4616 267608 4622
rect 267556 4558 267608 4564
rect 267660 4146 267688 7142
rect 267844 6798 267872 7783
rect 268016 7472 268068 7478
rect 268014 7440 268016 7449
rect 268068 7440 268070 7449
rect 268014 7375 268070 7384
rect 268016 7336 268068 7342
rect 268014 7304 268016 7313
rect 268200 7336 268252 7342
rect 268068 7304 268070 7313
rect 268200 7278 268252 7284
rect 268014 7239 268070 7248
rect 268014 7032 268070 7041
rect 268014 6967 268070 6976
rect 268028 6866 268056 6967
rect 268106 6896 268162 6905
rect 268016 6860 268068 6866
rect 268106 6831 268162 6840
rect 268016 6802 268068 6808
rect 267832 6792 267884 6798
rect 267832 6734 267884 6740
rect 267832 6316 267884 6322
rect 267832 6258 267884 6264
rect 267740 5840 267792 5846
rect 267738 5808 267740 5817
rect 267792 5808 267794 5817
rect 267738 5743 267794 5752
rect 267738 5672 267794 5681
rect 267738 5607 267794 5616
rect 267752 5370 267780 5607
rect 267844 5370 267872 6258
rect 268120 6186 268148 6831
rect 268212 6497 268240 7278
rect 268198 6488 268254 6497
rect 268198 6423 268254 6432
rect 268304 6202 268332 7822
rect 268384 7404 268436 7410
rect 268384 7346 268436 7352
rect 268396 6361 268424 7346
rect 268382 6352 268438 6361
rect 268488 6322 268516 9454
rect 268568 8832 268620 8838
rect 268568 8774 268620 8780
rect 268580 8498 268608 8774
rect 268568 8492 268620 8498
rect 268568 8434 268620 8440
rect 268568 7812 268620 7818
rect 268568 7754 268620 7760
rect 268382 6287 268438 6296
rect 268476 6316 268528 6322
rect 268476 6258 268528 6264
rect 268108 6180 268160 6186
rect 268108 6122 268160 6128
rect 268212 6174 268332 6202
rect 268212 5953 268240 6174
rect 268198 5944 268254 5953
rect 268198 5879 268254 5888
rect 268474 5944 268530 5953
rect 268474 5879 268530 5888
rect 268014 5808 268070 5817
rect 268014 5743 268070 5752
rect 267922 5672 267978 5681
rect 267922 5607 267978 5616
rect 267740 5364 267792 5370
rect 267740 5306 267792 5312
rect 267832 5364 267884 5370
rect 267832 5306 267884 5312
rect 267738 4720 267794 4729
rect 267738 4655 267740 4664
rect 267792 4655 267794 4664
rect 267740 4626 267792 4632
rect 267648 4140 267700 4146
rect 267648 4082 267700 4088
rect 267936 4010 267964 5607
rect 268028 4162 268056 5743
rect 268292 5160 268344 5166
rect 268292 5102 268344 5108
rect 268382 5128 268438 5137
rect 268106 4992 268162 5001
rect 268106 4927 268162 4936
rect 268120 4282 268148 4927
rect 268200 4616 268252 4622
rect 268200 4558 268252 4564
rect 268212 4282 268240 4558
rect 268108 4276 268160 4282
rect 268108 4218 268160 4224
rect 268200 4276 268252 4282
rect 268200 4218 268252 4224
rect 268028 4134 268240 4162
rect 268014 4040 268070 4049
rect 267924 4004 267976 4010
rect 268014 3975 268070 3984
rect 267924 3946 267976 3952
rect 268028 3777 268056 3975
rect 268014 3768 268070 3777
rect 267660 3726 267964 3754
rect 267660 3466 267688 3726
rect 267936 3641 267964 3726
rect 268014 3703 268070 3712
rect 268016 3664 268068 3670
rect 267738 3632 267794 3641
rect 267738 3567 267794 3576
rect 267922 3632 267978 3641
rect 268016 3606 268068 3612
rect 267922 3567 267978 3576
rect 267752 3534 267780 3567
rect 267740 3528 267792 3534
rect 267740 3470 267792 3476
rect 267648 3460 267700 3466
rect 267648 3402 267700 3408
rect 267740 3392 267792 3398
rect 267738 3360 267740 3369
rect 267792 3360 267794 3369
rect 267738 3295 267794 3304
rect 267464 3052 267516 3058
rect 267464 2994 267516 3000
rect 268028 2961 268056 3606
rect 268108 3596 268160 3602
rect 268108 3538 268160 3544
rect 268120 3233 268148 3538
rect 268212 3534 268240 4134
rect 268200 3528 268252 3534
rect 268200 3470 268252 3476
rect 268106 3224 268162 3233
rect 268106 3159 268162 3168
rect 268304 2990 268332 5102
rect 268382 5063 268438 5072
rect 268396 4162 268424 5063
rect 268488 4554 268516 5879
rect 268580 4826 268608 7754
rect 268672 5642 268700 9454
rect 268856 8537 268884 9522
rect 268948 9353 268976 10066
rect 269028 10056 269080 10062
rect 269026 10024 269028 10033
rect 269080 10024 269082 10033
rect 269026 9959 269082 9968
rect 269488 9580 269540 9586
rect 269488 9522 269540 9528
rect 269304 9376 269356 9382
rect 268934 9344 268990 9353
rect 269304 9318 269356 9324
rect 268934 9279 268990 9288
rect 269316 8838 269344 9318
rect 269500 8906 269528 9522
rect 270420 9518 270448 10134
rect 271337 9820 271645 9829
rect 271337 9818 271343 9820
rect 271399 9818 271423 9820
rect 271479 9818 271503 9820
rect 271559 9818 271583 9820
rect 271639 9818 271645 9820
rect 271399 9766 271401 9818
rect 271581 9766 271583 9818
rect 271337 9764 271343 9766
rect 271399 9764 271423 9766
rect 271479 9764 271503 9766
rect 271559 9764 271583 9766
rect 271639 9764 271645 9766
rect 271337 9755 271645 9764
rect 271236 9580 271288 9586
rect 271236 9522 271288 9528
rect 270408 9512 270460 9518
rect 270408 9454 270460 9460
rect 269856 9376 269908 9382
rect 269856 9318 269908 9324
rect 270408 9376 270460 9382
rect 270408 9318 270460 9324
rect 269488 8900 269540 8906
rect 269488 8842 269540 8848
rect 269304 8832 269356 8838
rect 269304 8774 269356 8780
rect 268842 8528 268898 8537
rect 268752 8492 268804 8498
rect 268842 8463 268898 8472
rect 268752 8434 268804 8440
rect 268764 8294 268792 8434
rect 268752 8288 268804 8294
rect 268752 8230 268804 8236
rect 268750 7984 268806 7993
rect 268750 7919 268806 7928
rect 268764 7818 268792 7919
rect 268752 7812 268804 7818
rect 268752 7754 268804 7760
rect 268750 6488 268806 6497
rect 268750 6423 268806 6432
rect 268660 5636 268712 5642
rect 268660 5578 268712 5584
rect 268660 5228 268712 5234
rect 268660 5170 268712 5176
rect 268568 4820 268620 4826
rect 268568 4762 268620 4768
rect 268476 4548 268528 4554
rect 268476 4490 268528 4496
rect 268568 4548 268620 4554
rect 268568 4490 268620 4496
rect 268580 4321 268608 4490
rect 268566 4312 268622 4321
rect 268566 4247 268622 4256
rect 268396 4134 268608 4162
rect 268672 4146 268700 5170
rect 268384 4072 268436 4078
rect 268384 4014 268436 4020
rect 268474 4040 268530 4049
rect 268292 2984 268344 2990
rect 268014 2952 268070 2961
rect 268292 2926 268344 2932
rect 268014 2887 268070 2896
rect 268198 2816 268254 2825
rect 268198 2751 268254 2760
rect 267280 2442 267332 2448
rect 267280 2384 267332 2390
rect 268212 2310 268240 2751
rect 268396 2650 268424 4014
rect 268474 3975 268530 3984
rect 268488 3194 268516 3975
rect 268476 3188 268528 3194
rect 268476 3130 268528 3136
rect 268476 2848 268528 2854
rect 268476 2790 268528 2796
rect 268384 2644 268436 2650
rect 268384 2586 268436 2592
rect 268488 2553 268516 2790
rect 268290 2544 268346 2553
rect 268290 2479 268346 2488
rect 268474 2544 268530 2553
rect 268474 2479 268530 2488
rect 267556 2304 267608 2310
rect 267556 2246 267608 2252
rect 268200 2304 268252 2310
rect 268200 2246 268252 2252
rect 267568 2038 267596 2246
rect 267556 2032 267608 2038
rect 267556 1974 267608 1980
rect 268304 1902 268332 2479
rect 268580 2446 268608 4134
rect 268660 4140 268712 4146
rect 268660 4082 268712 4088
rect 268764 3534 268792 6423
rect 268856 5642 268884 8463
rect 269316 8430 269344 8774
rect 269500 8498 269528 8842
rect 269488 8492 269540 8498
rect 269488 8434 269540 8440
rect 269304 8424 269356 8430
rect 269304 8366 269356 8372
rect 269672 8424 269724 8430
rect 269672 8366 269724 8372
rect 268936 8356 268988 8362
rect 268936 8298 268988 8304
rect 268948 8129 268976 8298
rect 268934 8120 268990 8129
rect 268934 8055 268990 8064
rect 269028 7948 269080 7954
rect 269028 7890 269080 7896
rect 269040 6633 269068 7890
rect 269488 7404 269540 7410
rect 269488 7346 269540 7352
rect 269396 7200 269448 7206
rect 269396 7142 269448 7148
rect 269212 6792 269264 6798
rect 269212 6734 269264 6740
rect 269026 6624 269082 6633
rect 269026 6559 269082 6568
rect 269224 6458 269252 6734
rect 269212 6452 269264 6458
rect 269212 6394 269264 6400
rect 269118 6352 269174 6361
rect 269118 6287 269174 6296
rect 269132 6254 269160 6287
rect 269120 6248 269172 6254
rect 268934 6216 268990 6225
rect 269120 6190 269172 6196
rect 268934 6151 268990 6160
rect 268844 5636 268896 5642
rect 268844 5578 268896 5584
rect 268948 5545 268976 6151
rect 269028 6112 269080 6118
rect 269026 6080 269028 6089
rect 269080 6080 269082 6089
rect 269026 6015 269082 6024
rect 269028 5704 269080 5710
rect 269028 5646 269080 5652
rect 268934 5536 268990 5545
rect 268934 5471 268990 5480
rect 268842 5400 268898 5409
rect 269040 5370 269068 5646
rect 269224 5642 269252 6394
rect 269408 6322 269436 7142
rect 269500 6798 269528 7346
rect 269488 6792 269540 6798
rect 269488 6734 269540 6740
rect 269396 6316 269448 6322
rect 269396 6258 269448 6264
rect 269488 5704 269540 5710
rect 269394 5672 269450 5681
rect 269212 5636 269264 5642
rect 269488 5646 269540 5652
rect 269578 5672 269634 5681
rect 269394 5607 269450 5616
rect 269212 5578 269264 5584
rect 268842 5335 268898 5344
rect 269028 5364 269080 5370
rect 268856 5098 268884 5335
rect 269028 5306 269080 5312
rect 268934 5264 268990 5273
rect 268934 5199 268990 5208
rect 268844 5092 268896 5098
rect 268844 5034 268896 5040
rect 268842 4856 268898 4865
rect 268842 4791 268898 4800
rect 268856 4214 268884 4791
rect 268844 4208 268896 4214
rect 268844 4150 268896 4156
rect 268844 4072 268896 4078
rect 268844 4014 268896 4020
rect 268752 3528 268804 3534
rect 268752 3470 268804 3476
rect 268856 3346 268884 4014
rect 268672 3318 268884 3346
rect 268672 3058 268700 3318
rect 268660 3052 268712 3058
rect 268660 2994 268712 3000
rect 268948 2774 268976 5199
rect 269304 5160 269356 5166
rect 269304 5102 269356 5108
rect 269212 5092 269264 5098
rect 269212 5034 269264 5040
rect 269120 4616 269172 4622
rect 269120 4558 269172 4564
rect 269028 3936 269080 3942
rect 269028 3878 269080 3884
rect 269040 3466 269068 3878
rect 269028 3460 269080 3466
rect 269028 3402 269080 3408
rect 269132 2922 269160 4558
rect 269224 3670 269252 5034
rect 269212 3664 269264 3670
rect 269212 3606 269264 3612
rect 269316 3194 269344 5102
rect 269408 3942 269436 5607
rect 269396 3936 269448 3942
rect 269396 3878 269448 3884
rect 269500 3738 269528 5646
rect 269578 5607 269634 5616
rect 269488 3732 269540 3738
rect 269488 3674 269540 3680
rect 269592 3670 269620 5607
rect 269684 4146 269712 8366
rect 269764 5228 269816 5234
rect 269764 5170 269816 5176
rect 269776 4622 269804 5170
rect 269764 4616 269816 4622
rect 269764 4558 269816 4564
rect 269672 4140 269724 4146
rect 269672 4082 269724 4088
rect 269868 3670 269896 9318
rect 270420 8974 270448 9318
rect 270592 9036 270644 9042
rect 270592 8978 270644 8984
rect 270316 8968 270368 8974
rect 270316 8910 270368 8916
rect 270408 8968 270460 8974
rect 270408 8910 270460 8916
rect 270224 8628 270276 8634
rect 270224 8570 270276 8576
rect 270132 8424 270184 8430
rect 270132 8366 270184 8372
rect 270144 7993 270172 8366
rect 270130 7984 270186 7993
rect 270130 7919 270186 7928
rect 270040 7472 270092 7478
rect 270092 7432 270172 7460
rect 270040 7414 270092 7420
rect 270040 6248 270092 6254
rect 270040 6190 270092 6196
rect 269580 3664 269632 3670
rect 269580 3606 269632 3612
rect 269856 3664 269908 3670
rect 269856 3606 269908 3612
rect 269948 3528 270000 3534
rect 269948 3470 270000 3476
rect 269960 3194 269988 3470
rect 270052 3398 270080 6190
rect 270040 3392 270092 3398
rect 270040 3334 270092 3340
rect 269304 3188 269356 3194
rect 269304 3130 269356 3136
rect 269948 3188 270000 3194
rect 269948 3130 270000 3136
rect 269856 3052 269908 3058
rect 269856 2994 269908 3000
rect 269120 2916 269172 2922
rect 269120 2858 269172 2864
rect 268856 2746 268976 2774
rect 268568 2440 268620 2446
rect 268568 2382 268620 2388
rect 268856 2378 268884 2746
rect 269028 2576 269080 2582
rect 269028 2518 269080 2524
rect 268844 2372 268896 2378
rect 268844 2314 268896 2320
rect 268750 2272 268806 2281
rect 268750 2207 268806 2216
rect 265808 1896 265860 1902
rect 265808 1838 265860 1844
rect 266636 1896 266688 1902
rect 266636 1838 266688 1844
rect 266728 1896 266780 1902
rect 266728 1838 266780 1844
rect 268292 1896 268344 1902
rect 268292 1838 268344 1844
rect 265900 1760 265952 1766
rect 265900 1702 265952 1708
rect 266728 1760 266780 1766
rect 267832 1760 267884 1766
rect 266728 1702 266780 1708
rect 267646 1728 267702 1737
rect 265912 1358 265940 1702
rect 266740 1358 266768 1702
rect 267832 1702 267884 1708
rect 268200 1760 268252 1766
rect 268200 1702 268252 1708
rect 267646 1663 267702 1672
rect 267660 1442 267688 1663
rect 267660 1426 267780 1442
rect 267660 1420 267792 1426
rect 267660 1414 267740 1420
rect 267740 1362 267792 1368
rect 267844 1358 267872 1702
rect 268212 1358 268240 1702
rect 265900 1352 265952 1358
rect 265900 1294 265952 1300
rect 266728 1352 266780 1358
rect 266728 1294 266780 1300
rect 267832 1352 267884 1358
rect 267832 1294 267884 1300
rect 268200 1352 268252 1358
rect 268200 1294 268252 1300
rect 266084 1216 266136 1222
rect 266084 1158 266136 1164
rect 266912 1216 266964 1222
rect 266912 1158 266964 1164
rect 267648 1216 267700 1222
rect 267648 1158 267700 1164
rect 268384 1216 268436 1222
rect 268384 1158 268436 1164
rect 265532 1012 265584 1018
rect 265532 954 265584 960
rect 266096 649 266124 1158
rect 266924 649 266952 1158
rect 267660 649 267688 1158
rect 268396 649 268424 1158
rect 268764 1057 268792 2207
rect 269040 2145 269068 2518
rect 269212 2440 269264 2446
rect 269212 2382 269264 2388
rect 269672 2440 269724 2446
rect 269672 2382 269724 2388
rect 268842 2136 268898 2145
rect 268842 2071 268898 2080
rect 269026 2136 269082 2145
rect 269026 2071 269082 2080
rect 268856 1465 268884 2071
rect 269224 1970 269252 2382
rect 269684 2106 269712 2382
rect 269672 2100 269724 2106
rect 269672 2042 269724 2048
rect 269764 2100 269816 2106
rect 269764 2042 269816 2048
rect 269776 1970 269804 2042
rect 269212 1964 269264 1970
rect 269212 1906 269264 1912
rect 269764 1964 269816 1970
rect 269764 1906 269816 1912
rect 269028 1828 269080 1834
rect 269028 1770 269080 1776
rect 269040 1601 269068 1770
rect 269026 1592 269082 1601
rect 269026 1527 269082 1536
rect 268842 1456 268898 1465
rect 268842 1391 268898 1400
rect 269224 1358 269252 1906
rect 269868 1358 269896 2994
rect 270144 2514 270172 7432
rect 270236 4554 270264 8570
rect 270328 8129 270356 8910
rect 270604 8537 270632 8978
rect 270776 8900 270828 8906
rect 270776 8842 270828 8848
rect 270590 8528 270646 8537
rect 270590 8463 270646 8472
rect 270498 8256 270554 8265
rect 270498 8191 270554 8200
rect 270314 8120 270370 8129
rect 270314 8055 270370 8064
rect 270512 7410 270540 8191
rect 270684 7540 270736 7546
rect 270684 7482 270736 7488
rect 270500 7404 270552 7410
rect 270500 7346 270552 7352
rect 270500 6792 270552 6798
rect 270500 6734 270552 6740
rect 270408 6724 270460 6730
rect 270408 6666 270460 6672
rect 270420 6322 270448 6666
rect 270408 6316 270460 6322
rect 270408 6258 270460 6264
rect 270316 6112 270368 6118
rect 270316 6054 270368 6060
rect 270328 5817 270356 6054
rect 270314 5808 270370 5817
rect 270314 5743 270370 5752
rect 270420 5710 270448 6258
rect 270512 5914 270540 6734
rect 270500 5908 270552 5914
rect 270500 5850 270552 5856
rect 270590 5808 270646 5817
rect 270590 5743 270646 5752
rect 270408 5704 270460 5710
rect 270408 5646 270460 5652
rect 270498 5672 270554 5681
rect 270420 5234 270448 5646
rect 270498 5607 270554 5616
rect 270408 5228 270460 5234
rect 270408 5170 270460 5176
rect 270224 4548 270276 4554
rect 270224 4490 270276 4496
rect 270512 3942 270540 5607
rect 270500 3936 270552 3942
rect 270500 3878 270552 3884
rect 270604 3738 270632 5743
rect 270696 4146 270724 7482
rect 270684 4140 270736 4146
rect 270684 4082 270736 4088
rect 270788 3738 270816 8842
rect 271052 8832 271104 8838
rect 271052 8774 271104 8780
rect 270868 8492 270920 8498
rect 270868 8434 270920 8440
rect 270880 4146 270908 8434
rect 270960 6996 271012 7002
rect 270960 6938 271012 6944
rect 270972 4826 271000 6938
rect 270960 4820 271012 4826
rect 270960 4762 271012 4768
rect 270868 4140 270920 4146
rect 270868 4082 270920 4088
rect 270592 3732 270644 3738
rect 270592 3674 270644 3680
rect 270776 3732 270828 3738
rect 270776 3674 270828 3680
rect 270774 3224 270830 3233
rect 270774 3159 270830 3168
rect 270500 2848 270552 2854
rect 270498 2816 270500 2825
rect 270788 2825 270816 3159
rect 270552 2816 270554 2825
rect 270498 2751 270554 2760
rect 270774 2816 270830 2825
rect 271064 2774 271092 8774
rect 271248 8401 271276 9522
rect 271786 9480 271842 9489
rect 271842 9438 272012 9466
rect 271786 9415 271842 9424
rect 271984 8945 272012 9438
rect 271970 8936 272026 8945
rect 271970 8871 272026 8880
rect 271337 8732 271645 8741
rect 271337 8730 271343 8732
rect 271399 8730 271423 8732
rect 271479 8730 271503 8732
rect 271559 8730 271583 8732
rect 271639 8730 271645 8732
rect 271399 8678 271401 8730
rect 271581 8678 271583 8730
rect 271337 8676 271343 8678
rect 271399 8676 271423 8678
rect 271479 8676 271503 8678
rect 271559 8676 271583 8678
rect 271639 8676 271645 8678
rect 271337 8667 271645 8676
rect 271234 8392 271290 8401
rect 271234 8327 271290 8336
rect 271788 7948 271840 7954
rect 271788 7890 271840 7896
rect 271800 7721 271828 7890
rect 271786 7712 271842 7721
rect 271337 7644 271645 7653
rect 271786 7647 271842 7656
rect 271337 7642 271343 7644
rect 271399 7642 271423 7644
rect 271479 7642 271503 7644
rect 271559 7642 271583 7644
rect 271639 7642 271645 7644
rect 271399 7590 271401 7642
rect 271581 7590 271583 7642
rect 271337 7588 271343 7590
rect 271399 7588 271423 7590
rect 271479 7588 271503 7590
rect 271559 7588 271583 7590
rect 271639 7588 271645 7590
rect 271142 7576 271198 7585
rect 271337 7579 271645 7588
rect 271142 7511 271198 7520
rect 271786 7576 271842 7585
rect 271786 7511 271842 7520
rect 271156 7342 271184 7511
rect 271144 7336 271196 7342
rect 271800 7313 271828 7511
rect 271972 7336 272024 7342
rect 271144 7278 271196 7284
rect 271786 7304 271842 7313
rect 271786 7239 271842 7248
rect 271970 7304 271972 7313
rect 272024 7304 272026 7313
rect 271970 7239 272026 7248
rect 271694 6760 271750 6769
rect 271694 6695 271750 6704
rect 272062 6760 272118 6769
rect 272062 6695 272118 6704
rect 271337 6556 271645 6565
rect 271337 6554 271343 6556
rect 271399 6554 271423 6556
rect 271479 6554 271503 6556
rect 271559 6554 271583 6556
rect 271639 6554 271645 6556
rect 271399 6502 271401 6554
rect 271581 6502 271583 6554
rect 271337 6500 271343 6502
rect 271399 6500 271423 6502
rect 271479 6500 271503 6502
rect 271559 6500 271583 6502
rect 271639 6500 271645 6502
rect 271337 6491 271645 6500
rect 271708 5953 271736 6695
rect 271878 6624 271934 6633
rect 271878 6559 271934 6568
rect 271786 6080 271842 6089
rect 271786 6015 271842 6024
rect 271694 5944 271750 5953
rect 271694 5879 271750 5888
rect 271800 5760 271828 6015
rect 271708 5732 271828 5760
rect 271337 5468 271645 5477
rect 271337 5466 271343 5468
rect 271399 5466 271423 5468
rect 271479 5466 271503 5468
rect 271559 5466 271583 5468
rect 271639 5466 271645 5468
rect 271399 5414 271401 5466
rect 271581 5414 271583 5466
rect 271337 5412 271343 5414
rect 271399 5412 271423 5414
rect 271479 5412 271503 5414
rect 271559 5412 271583 5414
rect 271639 5412 271645 5414
rect 271142 5400 271198 5409
rect 271337 5403 271645 5412
rect 271142 5335 271144 5344
rect 271196 5335 271198 5344
rect 271144 5306 271196 5312
rect 271144 4616 271196 4622
rect 271144 4558 271196 4564
rect 271156 4457 271184 4558
rect 271142 4448 271198 4457
rect 271142 4383 271198 4392
rect 271337 4380 271645 4389
rect 271337 4378 271343 4380
rect 271399 4378 271423 4380
rect 271479 4378 271503 4380
rect 271559 4378 271583 4380
rect 271639 4378 271645 4380
rect 271399 4326 271401 4378
rect 271581 4326 271583 4378
rect 271337 4324 271343 4326
rect 271399 4324 271423 4326
rect 271479 4324 271503 4326
rect 271559 4324 271583 4326
rect 271639 4324 271645 4326
rect 271337 4315 271645 4324
rect 271708 4214 271736 5732
rect 271786 5536 271842 5545
rect 271786 5471 271842 5480
rect 271800 5137 271828 5471
rect 271786 5128 271842 5137
rect 271786 5063 271842 5072
rect 271696 4208 271748 4214
rect 271696 4150 271748 4156
rect 271142 4040 271198 4049
rect 271198 3998 271644 4026
rect 271142 3975 271198 3984
rect 271616 3777 271644 3998
rect 271602 3768 271658 3777
rect 271602 3703 271658 3712
rect 271142 3360 271198 3369
rect 271142 3295 271198 3304
rect 271156 3194 271184 3295
rect 271337 3292 271645 3301
rect 271337 3290 271343 3292
rect 271399 3290 271423 3292
rect 271479 3290 271503 3292
rect 271559 3290 271583 3292
rect 271639 3290 271645 3292
rect 271399 3238 271401 3290
rect 271581 3238 271583 3290
rect 271337 3236 271343 3238
rect 271399 3236 271423 3238
rect 271479 3236 271503 3238
rect 271559 3236 271583 3238
rect 271639 3236 271645 3238
rect 271337 3227 271645 3236
rect 271786 3224 271842 3233
rect 271144 3188 271196 3194
rect 271786 3159 271842 3168
rect 271144 3130 271196 3136
rect 271800 2961 271828 3159
rect 271892 3058 271920 6559
rect 271970 6352 272026 6361
rect 271970 6287 272026 6296
rect 271984 6118 272012 6287
rect 271972 6112 272024 6118
rect 271972 6054 272024 6060
rect 271970 5400 272026 5409
rect 271970 5335 271972 5344
rect 272024 5335 272026 5344
rect 271972 5306 272024 5312
rect 271970 5128 272026 5137
rect 271970 5063 272026 5072
rect 271984 5030 272012 5063
rect 271972 5024 272024 5030
rect 271972 4966 272024 4972
rect 271970 3496 272026 3505
rect 271970 3431 271972 3440
rect 272024 3431 272026 3440
rect 271972 3402 272024 3408
rect 271972 3188 272024 3194
rect 271972 3130 272024 3136
rect 271880 3052 271932 3058
rect 271880 2994 271932 3000
rect 271984 2961 272012 3130
rect 272076 3126 272104 6695
rect 272154 4720 272210 4729
rect 272154 4655 272210 4664
rect 272168 4622 272196 4655
rect 272156 4616 272208 4622
rect 272156 4558 272208 4564
rect 272064 3120 272116 3126
rect 272064 3062 272116 3068
rect 271786 2952 271842 2961
rect 271786 2887 271842 2896
rect 271970 2952 272026 2961
rect 271970 2887 272026 2896
rect 270774 2751 270830 2760
rect 270880 2746 271092 2774
rect 270132 2508 270184 2514
rect 270132 2450 270184 2456
rect 270500 2440 270552 2446
rect 270500 2382 270552 2388
rect 269948 2304 270000 2310
rect 269948 2246 270000 2252
rect 270040 2304 270092 2310
rect 270040 2246 270092 2252
rect 269960 1358 269988 2246
rect 269212 1352 269264 1358
rect 269212 1294 269264 1300
rect 269856 1352 269908 1358
rect 269856 1294 269908 1300
rect 269948 1352 270000 1358
rect 269948 1294 270000 1300
rect 268936 1284 268988 1290
rect 268936 1226 268988 1232
rect 268750 1048 268806 1057
rect 268750 983 268806 992
rect 262494 640 262550 649
rect 262494 575 262550 584
rect 263230 640 263286 649
rect 263230 575 263286 584
rect 264334 640 264390 649
rect 264334 575 264390 584
rect 265346 640 265402 649
rect 265346 575 265402 584
rect 266082 640 266138 649
rect 266082 575 266138 584
rect 266910 640 266966 649
rect 266910 575 266966 584
rect 267646 640 267702 649
rect 267646 575 267702 584
rect 268382 640 268438 649
rect 268382 575 268438 584
rect 261850 504 261906 513
rect 256516 468 256568 474
rect 261850 439 261906 448
rect 256516 410 256568 416
rect 268948 406 268976 1226
rect 269028 1012 269080 1018
rect 269028 954 269080 960
rect 269040 921 269068 954
rect 269026 912 269082 921
rect 269026 847 269082 856
rect 270052 513 270080 2246
rect 270512 2106 270540 2382
rect 270776 2304 270828 2310
rect 270776 2246 270828 2252
rect 270500 2100 270552 2106
rect 270500 2042 270552 2048
rect 270316 1216 270368 1222
rect 270316 1158 270368 1164
rect 270328 649 270356 1158
rect 270314 640 270370 649
rect 270314 575 270370 584
rect 270038 504 270094 513
rect 270038 439 270094 448
rect 268936 400 268988 406
rect 255134 368 255190 377
rect 240966 303 241022 312
rect 251824 332 251876 338
rect 229744 264 229796 270
rect 229744 206 229796 212
rect 239600 105 239628 303
rect 270788 377 270816 2246
rect 270880 1902 270908 2746
rect 271970 2408 272026 2417
rect 271970 2343 272026 2352
rect 271142 2272 271198 2281
rect 271142 2207 271198 2216
rect 271156 2038 271184 2207
rect 271337 2204 271645 2213
rect 271337 2202 271343 2204
rect 271399 2202 271423 2204
rect 271479 2202 271503 2204
rect 271559 2202 271583 2204
rect 271639 2202 271645 2204
rect 271399 2150 271401 2202
rect 271581 2150 271583 2202
rect 271337 2148 271343 2150
rect 271399 2148 271423 2150
rect 271479 2148 271503 2150
rect 271559 2148 271583 2150
rect 271639 2148 271645 2150
rect 271337 2139 271645 2148
rect 271786 2136 271842 2145
rect 271786 2071 271842 2080
rect 271144 2032 271196 2038
rect 271144 1974 271196 1980
rect 270868 1896 270920 1902
rect 270868 1838 270920 1844
rect 271800 1290 271828 2071
rect 271984 2009 272012 2343
rect 272156 2032 272208 2038
rect 271970 2000 272026 2009
rect 271970 1935 272026 1944
rect 272154 2000 272156 2009
rect 272208 2000 272210 2009
rect 272154 1935 272210 1944
rect 271788 1284 271840 1290
rect 271788 1226 271840 1232
rect 271786 1184 271842 1193
rect 271337 1116 271645 1125
rect 271786 1119 271842 1128
rect 271337 1114 271343 1116
rect 271399 1114 271423 1116
rect 271479 1114 271503 1116
rect 271559 1114 271583 1116
rect 271639 1114 271645 1116
rect 271399 1062 271401 1114
rect 271581 1062 271583 1114
rect 271337 1060 271343 1062
rect 271399 1060 271423 1062
rect 271479 1060 271503 1062
rect 271559 1060 271583 1062
rect 271639 1060 271645 1062
rect 271337 1051 271645 1060
rect 268936 342 268988 348
rect 270774 368 270830 377
rect 255134 303 255190 312
rect 270774 303 270830 312
rect 251824 274 251876 280
rect 271800 105 271828 1119
rect 180890 96 180946 105
rect 180890 31 180946 40
rect 224774 96 224830 105
rect 224774 31 224830 40
rect 224958 96 225014 105
rect 224958 31 225014 40
rect 239586 96 239642 105
rect 239586 31 239642 40
rect 271786 96 271842 105
rect 271786 31 271842 40
<< via2 >>
rect 227442 10820 227444 10840
rect 227444 10820 227496 10840
rect 227496 10820 227498 10840
rect 9678 10512 9734 10568
rect 20718 10512 20774 10568
rect 1674 10104 1730 10160
rect 2410 10104 2466 10160
rect 3238 10104 3294 10160
rect 4342 10104 4398 10160
rect 5078 10104 5134 10160
rect 5814 10104 5870 10160
rect 6826 10104 6882 10160
rect 7562 10104 7618 10160
rect 3146 9832 3202 9888
rect 1398 9172 1454 9208
rect 1398 9152 1400 9172
rect 1400 9152 1452 9172
rect 1452 9152 1454 9172
rect 8390 10104 8446 10160
rect 8206 9832 8262 9888
rect 11978 10104 12034 10160
rect 12714 10104 12770 10160
rect 13726 10104 13782 10160
rect 14646 10104 14702 10160
rect 15382 10104 15438 10160
rect 16118 10104 16174 10160
rect 17130 10104 17186 10160
rect 17866 10104 17922 10160
rect 18602 10104 18658 10160
rect 22374 10104 22430 10160
rect 10506 9832 10562 9888
rect 11242 9832 11298 9888
rect 13450 9832 13506 9888
rect 21454 9832 21510 9888
rect 19246 6840 19302 6896
rect 19982 6840 20038 6896
rect 20718 5072 20774 5128
rect 846 1420 902 1456
rect 846 1400 848 1420
rect 848 1400 900 1420
rect 900 1400 902 1420
rect 1582 1264 1638 1320
rect 2318 992 2374 1048
rect 2962 720 3018 776
rect 4526 992 4582 1048
rect 5170 720 5226 776
rect 4066 584 4122 640
rect 6826 992 6882 1048
rect 6550 720 6606 776
rect 7562 720 7618 776
rect 8206 584 8262 640
rect 9034 720 9090 776
rect 9586 584 9642 640
rect 10414 1128 10470 1184
rect 19338 4392 19394 4448
rect 23478 8628 23534 8664
rect 23478 8608 23480 8628
rect 23480 8608 23532 8628
rect 23532 8608 23534 8628
rect 23478 6840 23534 6896
rect 19246 2932 19248 2952
rect 19248 2932 19300 2952
rect 19300 2932 19302 2952
rect 19246 2896 19302 2932
rect 22926 2916 22982 2952
rect 22926 2896 22928 2916
rect 22928 2896 22980 2916
rect 22980 2896 22982 2916
rect 19982 2796 19984 2816
rect 19984 2796 20036 2816
rect 20036 2796 20038 2816
rect 19982 2760 20038 2796
rect 23386 2760 23442 2816
rect 24030 8780 24032 8800
rect 24032 8780 24084 8800
rect 24084 8780 24086 8800
rect 24030 8744 24086 8780
rect 24766 6840 24822 6896
rect 15842 1964 15898 2000
rect 15842 1944 15844 1964
rect 15844 1944 15896 1964
rect 15896 1944 15898 1964
rect 14094 992 14150 1048
rect 22190 1672 22246 1728
rect 16578 1400 16634 1456
rect 22098 1400 22154 1456
rect 25686 8744 25742 8800
rect 25870 9560 25926 9616
rect 24490 3304 24546 3360
rect 25226 3032 25282 3088
rect 26698 8336 26754 8392
rect 26238 6840 26294 6896
rect 28814 9444 28870 9480
rect 28814 9424 28816 9444
rect 28816 9424 28868 9444
rect 28868 9424 28870 9444
rect 28354 8336 28410 8392
rect 27894 7792 27950 7848
rect 28078 2760 28134 2816
rect 25962 1264 26018 1320
rect 26698 1264 26754 1320
rect 27434 1264 27490 1320
rect 14830 720 14886 776
rect 15658 720 15714 776
rect 10230 584 10286 640
rect 10966 584 11022 640
rect 11978 584 12034 640
rect 12714 584 12770 640
rect 13450 584 13506 640
rect 17130 584 17186 640
rect 17866 584 17922 640
rect 18602 584 18658 640
rect 23938 584 23994 640
rect 29642 8628 29698 8664
rect 29642 8608 29644 8628
rect 29644 8608 29696 8628
rect 29696 8608 29698 8628
rect 54666 10376 54722 10432
rect 31758 10240 31814 10296
rect 35162 10240 35218 10296
rect 35622 10240 35678 10296
rect 36266 10240 36322 10296
rect 36910 10240 36966 10296
rect 38106 10240 38162 10296
rect 38842 10240 38898 10296
rect 39486 10240 39542 10296
rect 40314 10240 40370 10296
rect 40774 10240 40830 10296
rect 41418 10240 41474 10296
rect 42062 10240 42118 10296
rect 43258 10240 43314 10296
rect 43994 10240 44050 10296
rect 44638 10240 44694 10296
rect 45466 10240 45522 10296
rect 45926 10240 45982 10296
rect 46570 10240 46626 10296
rect 47214 10240 47270 10296
rect 48226 10240 48282 10296
rect 49146 10240 49202 10296
rect 49790 10240 49846 10296
rect 50618 10240 50674 10296
rect 51354 10240 51410 10296
rect 52090 10240 52146 10296
rect 53010 10240 53066 10296
rect 53194 10240 53250 10296
rect 30194 8628 30250 8664
rect 30194 8608 30196 8628
rect 30196 8608 30248 8628
rect 30248 8608 30250 8628
rect 31298 8628 31354 8664
rect 31298 8608 31300 8628
rect 31300 8608 31352 8628
rect 31352 8608 31354 8628
rect 32586 9560 32642 9616
rect 34754 9274 34810 9276
rect 34834 9274 34890 9276
rect 34914 9274 34970 9276
rect 34994 9274 35050 9276
rect 34754 9222 34800 9274
rect 34800 9222 34810 9274
rect 34834 9222 34864 9274
rect 34864 9222 34876 9274
rect 34876 9222 34890 9274
rect 34914 9222 34928 9274
rect 34928 9222 34940 9274
rect 34940 9222 34970 9274
rect 34994 9222 35004 9274
rect 35004 9222 35050 9274
rect 34754 9220 34810 9222
rect 34834 9220 34890 9222
rect 34914 9220 34970 9222
rect 34994 9220 35050 9222
rect 34754 8186 34810 8188
rect 34834 8186 34890 8188
rect 34914 8186 34970 8188
rect 34994 8186 35050 8188
rect 34754 8134 34800 8186
rect 34800 8134 34810 8186
rect 34834 8134 34864 8186
rect 34864 8134 34876 8186
rect 34876 8134 34890 8186
rect 34914 8134 34928 8186
rect 34928 8134 34940 8186
rect 34940 8134 34970 8186
rect 34994 8134 35004 8186
rect 35004 8134 35050 8186
rect 34754 8132 34810 8134
rect 34834 8132 34890 8134
rect 34914 8132 34970 8134
rect 34994 8132 35050 8134
rect 34754 7098 34810 7100
rect 34834 7098 34890 7100
rect 34914 7098 34970 7100
rect 34994 7098 35050 7100
rect 34754 7046 34800 7098
rect 34800 7046 34810 7098
rect 34834 7046 34864 7098
rect 34864 7046 34876 7098
rect 34876 7046 34890 7098
rect 34914 7046 34928 7098
rect 34928 7046 34940 7098
rect 34940 7046 34970 7098
rect 34994 7046 35004 7098
rect 35004 7046 35050 7098
rect 34754 7044 34810 7046
rect 34834 7044 34890 7046
rect 34914 7044 34970 7046
rect 34994 7044 35050 7046
rect 34754 6010 34810 6012
rect 34834 6010 34890 6012
rect 34914 6010 34970 6012
rect 34994 6010 35050 6012
rect 34754 5958 34800 6010
rect 34800 5958 34810 6010
rect 34834 5958 34864 6010
rect 34864 5958 34876 6010
rect 34876 5958 34890 6010
rect 34914 5958 34928 6010
rect 34928 5958 34940 6010
rect 34940 5958 34970 6010
rect 34994 5958 35004 6010
rect 35004 5958 35050 6010
rect 34754 5956 34810 5958
rect 34834 5956 34890 5958
rect 34914 5956 34970 5958
rect 34994 5956 35050 5958
rect 34754 4922 34810 4924
rect 34834 4922 34890 4924
rect 34914 4922 34970 4924
rect 34994 4922 35050 4924
rect 34754 4870 34800 4922
rect 34800 4870 34810 4922
rect 34834 4870 34864 4922
rect 34864 4870 34876 4922
rect 34876 4870 34890 4922
rect 34914 4870 34928 4922
rect 34928 4870 34940 4922
rect 34940 4870 34970 4922
rect 34994 4870 35004 4922
rect 35004 4870 35050 4922
rect 34754 4868 34810 4870
rect 34834 4868 34890 4870
rect 34914 4868 34970 4870
rect 34994 4868 35050 4870
rect 34754 3834 34810 3836
rect 34834 3834 34890 3836
rect 34914 3834 34970 3836
rect 34994 3834 35050 3836
rect 34754 3782 34800 3834
rect 34800 3782 34810 3834
rect 34834 3782 34864 3834
rect 34864 3782 34876 3834
rect 34876 3782 34890 3834
rect 34914 3782 34928 3834
rect 34928 3782 34940 3834
rect 34940 3782 34970 3834
rect 34994 3782 35004 3834
rect 35004 3782 35050 3834
rect 34754 3780 34810 3782
rect 34834 3780 34890 3782
rect 34914 3780 34970 3782
rect 34994 3780 35050 3782
rect 34754 2746 34810 2748
rect 34834 2746 34890 2748
rect 34914 2746 34970 2748
rect 34994 2746 35050 2748
rect 34754 2694 34800 2746
rect 34800 2694 34810 2746
rect 34834 2694 34864 2746
rect 34864 2694 34876 2746
rect 34876 2694 34890 2746
rect 34914 2694 34928 2746
rect 34928 2694 34940 2746
rect 34940 2694 34970 2746
rect 34994 2694 35004 2746
rect 35004 2694 35050 2746
rect 34754 2692 34810 2694
rect 34834 2692 34890 2694
rect 34914 2692 34970 2694
rect 34994 2692 35050 2694
rect 34754 1658 34810 1660
rect 34834 1658 34890 1660
rect 34914 1658 34970 1660
rect 34994 1658 35050 1660
rect 34754 1606 34800 1658
rect 34800 1606 34810 1658
rect 34834 1606 34864 1658
rect 34864 1606 34876 1658
rect 34876 1606 34890 1658
rect 34914 1606 34928 1658
rect 34928 1606 34940 1658
rect 34940 1606 34970 1658
rect 34994 1606 35004 1658
rect 35004 1606 35050 1658
rect 34754 1604 34810 1606
rect 34834 1604 34890 1606
rect 34914 1604 34970 1606
rect 34994 1604 35050 1606
rect 35898 6432 35954 6488
rect 33138 1400 33194 1456
rect 28998 584 29054 640
rect 30378 584 30434 640
rect 28722 448 28778 504
rect 29918 448 29974 504
rect 32494 448 32550 504
rect 36818 1708 36820 1728
rect 36820 1708 36872 1728
rect 36872 1708 36874 1728
rect 36818 1672 36874 1708
rect 35622 584 35678 640
rect 36266 584 36322 640
rect 36910 584 36966 640
rect 38198 2352 38254 2408
rect 39118 3440 39174 3496
rect 38106 584 38162 640
rect 38566 584 38622 640
rect 31574 312 31630 368
rect 34426 312 34482 368
rect 39946 584 40002 640
rect 40314 1828 40370 1864
rect 40314 1808 40316 1828
rect 40316 1808 40368 1828
rect 40368 1808 40370 1828
rect 40958 4256 41014 4312
rect 41418 4256 41474 4312
rect 40774 584 40830 640
rect 38842 312 38898 368
rect 41142 2916 41198 2952
rect 41142 2896 41144 2916
rect 41144 2896 41196 2916
rect 41196 2896 41198 2916
rect 42062 5344 42118 5400
rect 42430 5108 42432 5128
rect 42432 5108 42484 5128
rect 42484 5108 42486 5128
rect 42430 5072 42486 5108
rect 42706 5652 42708 5672
rect 42708 5652 42760 5672
rect 42760 5652 42762 5672
rect 42706 5616 42762 5652
rect 42522 4936 42578 4992
rect 42246 4528 42302 4584
rect 43166 5752 43222 5808
rect 43626 5752 43682 5808
rect 43718 5652 43720 5672
rect 43720 5652 43772 5672
rect 43772 5652 43774 5672
rect 43718 5616 43774 5652
rect 43810 4936 43866 4992
rect 44086 6180 44142 6216
rect 44086 6160 44088 6180
rect 44088 6160 44140 6180
rect 44140 6160 44142 6180
rect 44546 5616 44602 5672
rect 44270 5072 44326 5128
rect 44270 4256 44326 4312
rect 41418 584 41474 640
rect 42062 584 42118 640
rect 43258 584 43314 640
rect 44638 5092 44694 5128
rect 44638 5072 44640 5092
rect 44640 5072 44692 5092
rect 44692 5072 44694 5092
rect 44362 992 44418 1048
rect 45374 5752 45430 5808
rect 46018 6452 46074 6488
rect 46018 6432 46020 6452
rect 46020 6432 46072 6452
rect 46072 6432 46074 6452
rect 46938 4428 46940 4448
rect 46940 4428 46992 4448
rect 46992 4428 46994 4448
rect 46938 4392 46994 4428
rect 47950 5344 48006 5400
rect 48134 4392 48190 4448
rect 49790 4020 49792 4040
rect 49792 4020 49844 4040
rect 49844 4020 49846 4040
rect 49790 3984 49846 4020
rect 49054 1944 49110 2000
rect 51630 4020 51632 4040
rect 51632 4020 51684 4040
rect 51684 4020 51686 4040
rect 51630 3984 51686 4020
rect 43994 584 44050 640
rect 44638 584 44694 640
rect 45466 584 45522 640
rect 45926 584 45982 640
rect 46570 584 46626 640
rect 47214 584 47270 640
rect 48318 584 48374 640
rect 49146 584 49202 640
rect 49790 584 49846 640
rect 50618 584 50674 640
rect 51078 584 51134 640
rect 51722 584 51778 640
rect 54758 10240 54814 10296
rect 55494 10240 55550 10296
rect 56230 10240 56286 10296
rect 57058 10240 57114 10296
rect 54390 3032 54446 3088
rect 53930 1400 53986 1456
rect 54390 1944 54446 2000
rect 54206 1400 54262 1456
rect 57794 10240 57850 10296
rect 58622 10240 58678 10296
rect 59266 10240 59322 10296
rect 60002 10240 60058 10296
rect 60830 10240 60886 10296
rect 59358 1536 59414 1592
rect 61566 10240 61622 10296
rect 62302 10240 62358 10296
rect 63406 10240 63462 10296
rect 63774 10240 63830 10296
rect 64602 10240 64658 10296
rect 65430 10240 65486 10296
rect 60738 4256 60794 4312
rect 60738 2760 60794 2816
rect 71318 10512 71374 10568
rect 74262 10512 74318 10568
rect 66166 10240 66222 10296
rect 66902 10240 66958 10296
rect 68552 9818 68608 9820
rect 68632 9818 68688 9820
rect 68712 9818 68768 9820
rect 68792 9818 68848 9820
rect 68552 9766 68598 9818
rect 68598 9766 68608 9818
rect 68632 9766 68662 9818
rect 68662 9766 68674 9818
rect 68674 9766 68688 9818
rect 68712 9766 68726 9818
rect 68726 9766 68738 9818
rect 68738 9766 68768 9818
rect 68792 9766 68802 9818
rect 68802 9766 68848 9818
rect 68552 9764 68608 9766
rect 68632 9764 68688 9766
rect 68712 9764 68768 9766
rect 68792 9764 68848 9766
rect 69110 9580 69166 9616
rect 69110 9560 69112 9580
rect 69112 9560 69164 9580
rect 69164 9560 69166 9580
rect 70306 9580 70362 9616
rect 70306 9560 70308 9580
rect 70308 9560 70360 9580
rect 70360 9560 70362 9580
rect 69570 9036 69626 9072
rect 69570 9016 69572 9036
rect 69572 9016 69624 9036
rect 69624 9016 69626 9036
rect 68552 8730 68608 8732
rect 68632 8730 68688 8732
rect 68712 8730 68768 8732
rect 68792 8730 68848 8732
rect 68552 8678 68598 8730
rect 68598 8678 68608 8730
rect 68632 8678 68662 8730
rect 68662 8678 68674 8730
rect 68674 8678 68688 8730
rect 68712 8678 68726 8730
rect 68726 8678 68738 8730
rect 68738 8678 68768 8730
rect 68792 8678 68802 8730
rect 68802 8678 68848 8730
rect 68552 8676 68608 8678
rect 68632 8676 68688 8678
rect 68712 8676 68768 8678
rect 68792 8676 68848 8678
rect 72054 10376 72110 10432
rect 72146 9580 72202 9616
rect 72146 9560 72148 9580
rect 72148 9560 72200 9580
rect 72200 9560 72202 9580
rect 73434 9036 73490 9072
rect 73434 9016 73436 9036
rect 73436 9016 73488 9036
rect 73488 9016 73490 9036
rect 68552 7642 68608 7644
rect 68632 7642 68688 7644
rect 68712 7642 68768 7644
rect 68792 7642 68848 7644
rect 68552 7590 68598 7642
rect 68598 7590 68608 7642
rect 68632 7590 68662 7642
rect 68662 7590 68674 7642
rect 68674 7590 68688 7642
rect 68712 7590 68726 7642
rect 68726 7590 68738 7642
rect 68738 7590 68768 7642
rect 68792 7590 68802 7642
rect 68802 7590 68848 7642
rect 68552 7588 68608 7590
rect 68632 7588 68688 7590
rect 68712 7588 68768 7590
rect 68792 7588 68848 7590
rect 68552 6554 68608 6556
rect 68632 6554 68688 6556
rect 68712 6554 68768 6556
rect 68792 6554 68848 6556
rect 68552 6502 68598 6554
rect 68598 6502 68608 6554
rect 68632 6502 68662 6554
rect 68662 6502 68674 6554
rect 68674 6502 68688 6554
rect 68712 6502 68726 6554
rect 68726 6502 68738 6554
rect 68738 6502 68768 6554
rect 68792 6502 68802 6554
rect 68802 6502 68848 6554
rect 68552 6500 68608 6502
rect 68632 6500 68688 6502
rect 68712 6500 68768 6502
rect 68792 6500 68848 6502
rect 74722 9580 74778 9616
rect 74722 9560 74724 9580
rect 74724 9560 74776 9580
rect 74776 9560 74778 9580
rect 74722 9036 74778 9072
rect 84566 10512 84622 10568
rect 86774 10512 86830 10568
rect 77206 10376 77262 10432
rect 82358 10376 82414 10432
rect 83830 10376 83886 10432
rect 76470 9696 76526 9752
rect 74722 9016 74724 9036
rect 74724 9016 74776 9036
rect 74776 9016 74778 9036
rect 68552 5466 68608 5468
rect 68632 5466 68688 5468
rect 68712 5466 68768 5468
rect 68792 5466 68848 5468
rect 68552 5414 68598 5466
rect 68598 5414 68608 5466
rect 68632 5414 68662 5466
rect 68662 5414 68674 5466
rect 68674 5414 68688 5466
rect 68712 5414 68726 5466
rect 68726 5414 68738 5466
rect 68738 5414 68768 5466
rect 68792 5414 68802 5466
rect 68802 5414 68848 5466
rect 68552 5412 68608 5414
rect 68632 5412 68688 5414
rect 68712 5412 68768 5414
rect 68792 5412 68848 5414
rect 67546 5208 67602 5264
rect 68552 4378 68608 4380
rect 68632 4378 68688 4380
rect 68712 4378 68768 4380
rect 68792 4378 68848 4380
rect 68552 4326 68598 4378
rect 68598 4326 68608 4378
rect 68632 4326 68662 4378
rect 68662 4326 68674 4378
rect 68674 4326 68688 4378
rect 68712 4326 68726 4378
rect 68726 4326 68738 4378
rect 68738 4326 68768 4378
rect 68792 4326 68802 4378
rect 68802 4326 68848 4378
rect 68552 4324 68608 4326
rect 68632 4324 68688 4326
rect 68712 4324 68768 4326
rect 68792 4324 68848 4326
rect 68552 3290 68608 3292
rect 68632 3290 68688 3292
rect 68712 3290 68768 3292
rect 68792 3290 68848 3292
rect 68552 3238 68598 3290
rect 68598 3238 68608 3290
rect 68632 3238 68662 3290
rect 68662 3238 68674 3290
rect 68674 3238 68688 3290
rect 68712 3238 68726 3290
rect 68726 3238 68738 3290
rect 68738 3238 68768 3290
rect 68792 3238 68802 3290
rect 68802 3238 68848 3290
rect 68552 3236 68608 3238
rect 68632 3236 68688 3238
rect 68712 3236 68768 3238
rect 68792 3236 68848 3238
rect 68552 2202 68608 2204
rect 68632 2202 68688 2204
rect 68712 2202 68768 2204
rect 68792 2202 68848 2204
rect 68552 2150 68598 2202
rect 68598 2150 68608 2202
rect 68632 2150 68662 2202
rect 68662 2150 68674 2202
rect 68674 2150 68688 2202
rect 68712 2150 68726 2202
rect 68726 2150 68738 2202
rect 68738 2150 68768 2202
rect 68792 2150 68802 2202
rect 68802 2150 68848 2202
rect 68552 2148 68608 2150
rect 68632 2148 68688 2150
rect 68712 2148 68768 2150
rect 68792 2148 68848 2150
rect 52366 584 52422 640
rect 53378 584 53434 640
rect 54850 584 54906 640
rect 55678 584 55734 640
rect 56230 584 56286 640
rect 57058 584 57114 640
rect 57794 584 57850 640
rect 58622 584 58678 640
rect 60830 584 60886 640
rect 61566 584 61622 640
rect 62302 584 62358 640
rect 62946 584 63002 640
rect 63774 584 63830 640
rect 64510 584 64566 640
rect 65614 584 65670 640
rect 68552 1114 68608 1116
rect 68632 1114 68688 1116
rect 68712 1114 68768 1116
rect 68792 1114 68848 1116
rect 68552 1062 68598 1114
rect 68598 1062 68608 1114
rect 68632 1062 68662 1114
rect 68662 1062 68674 1114
rect 68674 1062 68688 1114
rect 68712 1062 68726 1114
rect 68726 1062 68738 1114
rect 68738 1062 68768 1114
rect 68792 1062 68802 1114
rect 68802 1062 68848 1114
rect 68552 1060 68608 1062
rect 68632 1060 68688 1062
rect 68712 1060 68768 1062
rect 68792 1060 68848 1062
rect 77298 9580 77354 9616
rect 77298 9560 77300 9580
rect 77300 9560 77352 9580
rect 77352 9560 77354 9580
rect 79414 9696 79470 9752
rect 81622 9696 81678 9752
rect 78586 9036 78642 9072
rect 78586 9016 78588 9036
rect 78588 9016 78640 9036
rect 78640 9016 78642 9036
rect 79966 9580 80022 9616
rect 79966 9560 79968 9580
rect 79968 9560 80020 9580
rect 80020 9560 80022 9580
rect 79966 9036 80022 9072
rect 79966 9016 79968 9036
rect 79968 9016 80020 9036
rect 80020 9016 80022 9036
rect 79322 6704 79378 6760
rect 71318 1264 71374 1320
rect 70582 992 70638 1048
rect 72054 992 72110 1048
rect 69110 720 69166 776
rect 69570 720 69626 776
rect 72146 584 72202 640
rect 66166 448 66222 504
rect 67546 448 67602 504
rect 73526 1264 73582 1320
rect 74262 992 74318 1048
rect 74722 584 74778 640
rect 76470 1264 76526 1320
rect 75734 992 75790 1048
rect 82634 9580 82690 9616
rect 82634 9560 82636 9580
rect 82636 9560 82688 9580
rect 82688 9560 82690 9580
rect 81990 5772 82046 5808
rect 81990 5752 81992 5772
rect 81992 5752 82044 5772
rect 82044 5752 82046 5772
rect 80334 5244 80336 5264
rect 80336 5244 80388 5264
rect 80388 5244 80390 5264
rect 80334 5208 80390 5244
rect 80886 5228 80942 5264
rect 81898 5616 81954 5672
rect 80886 5208 80888 5228
rect 80888 5208 80940 5228
rect 80940 5208 80942 5228
rect 81438 4664 81494 4720
rect 85394 9832 85450 9888
rect 86498 9832 86554 9888
rect 90362 10240 90418 10296
rect 84106 7928 84162 7984
rect 82726 7792 82782 7848
rect 82634 7384 82690 7440
rect 85578 5636 85634 5672
rect 85578 5616 85580 5636
rect 85580 5616 85632 5636
rect 85632 5616 85634 5636
rect 82174 3168 82230 3224
rect 82358 3052 82414 3088
rect 82358 3032 82360 3052
rect 82360 3032 82412 3052
rect 82412 3032 82414 3052
rect 80058 1536 80114 1592
rect 81346 1536 81402 1592
rect 77206 992 77262 1048
rect 77942 1264 77998 1320
rect 79414 1264 79470 1320
rect 77574 856 77630 912
rect 82082 1264 82138 1320
rect 83830 1672 83886 1728
rect 83002 1536 83058 1592
rect 83738 1536 83794 1592
rect 78586 720 78642 776
rect 79966 720 80022 776
rect 82726 584 82782 640
rect 86590 7656 86646 7712
rect 87050 7520 87106 7576
rect 86590 6568 86646 6624
rect 85670 3576 85726 3632
rect 86590 3440 86646 3496
rect 85670 3340 85672 3360
rect 85672 3340 85724 3360
rect 85724 3340 85726 3360
rect 85670 3304 85726 3340
rect 84290 2352 84346 2408
rect 86406 2080 86462 2136
rect 85302 1128 85358 1184
rect 86130 992 86186 1048
rect 84474 720 84530 776
rect 85026 720 85082 776
rect 86774 720 86830 776
rect 83922 448 83978 504
rect 87510 1264 87566 1320
rect 88338 9172 88394 9208
rect 88338 9152 88340 9172
rect 88340 9152 88392 9172
rect 88392 9152 88394 9172
rect 88338 8628 88394 8664
rect 88338 8608 88340 8628
rect 88340 8608 88392 8628
rect 88392 8608 88394 8628
rect 88338 1808 88394 1864
rect 89718 8064 89774 8120
rect 89074 1944 89130 2000
rect 89074 1400 89130 1456
rect 89902 2488 89958 2544
rect 89810 2216 89866 2272
rect 89626 1944 89682 2000
rect 90454 8628 90510 8664
rect 90454 8608 90456 8628
rect 90456 8608 90508 8628
rect 90508 8608 90510 8628
rect 90086 2932 90088 2952
rect 90088 2932 90140 2952
rect 90140 2932 90142 2952
rect 90086 2896 90142 2932
rect 91834 8744 91890 8800
rect 91926 8628 91982 8664
rect 91926 8608 91928 8628
rect 91928 8608 91980 8628
rect 91980 8608 91982 8628
rect 91466 5344 91522 5400
rect 91742 5108 91744 5128
rect 91744 5108 91796 5128
rect 91796 5108 91798 5128
rect 91742 5072 91798 5108
rect 89350 1264 89406 1320
rect 87602 1128 87658 1184
rect 90638 720 90694 776
rect 93490 9716 93546 9752
rect 93490 9696 93492 9716
rect 93492 9696 93544 9716
rect 93544 9696 93546 9716
rect 93306 8336 93362 8392
rect 92662 6160 92718 6216
rect 92478 4428 92480 4448
rect 92480 4428 92532 4448
rect 92532 4428 92534 4448
rect 92478 4392 92534 4428
rect 92202 720 92258 776
rect 95974 9716 96030 9752
rect 95974 9696 95976 9716
rect 95976 9696 96028 9716
rect 96028 9696 96030 9716
rect 96342 9716 96398 9752
rect 96342 9696 96344 9716
rect 96344 9696 96396 9716
rect 96396 9696 96398 9716
rect 94594 8628 94650 8664
rect 94594 8608 94596 8628
rect 94596 8608 94648 8628
rect 94648 8608 94650 8628
rect 94870 8628 94926 8664
rect 94870 8608 94872 8628
rect 94872 8608 94924 8628
rect 94924 8608 94926 8628
rect 94502 6160 94558 6216
rect 94410 4664 94466 4720
rect 94318 4528 94374 4584
rect 95238 6296 95294 6352
rect 95882 3476 95884 3496
rect 95884 3476 95936 3496
rect 95936 3476 95938 3496
rect 95882 3440 95938 3476
rect 96158 4020 96160 4040
rect 96160 4020 96212 4040
rect 96212 4020 96214 4040
rect 96158 3984 96214 4020
rect 96618 3596 96674 3632
rect 96618 3576 96620 3596
rect 96620 3576 96672 3596
rect 96672 3576 96674 3596
rect 93858 1128 93914 1184
rect 94594 1128 94650 1184
rect 95330 1128 95386 1184
rect 96066 1128 96122 1184
rect 93490 720 93546 776
rect 97446 8628 97502 8664
rect 97446 8608 97448 8628
rect 97448 8608 97500 8628
rect 97500 8608 97502 8628
rect 97998 9716 98054 9752
rect 97998 9696 98000 9716
rect 98000 9696 98052 9716
rect 98052 9696 98054 9716
rect 98090 4256 98146 4312
rect 97630 2624 97686 2680
rect 103242 10240 103298 10296
rect 100666 9716 100722 9752
rect 100666 9696 100668 9716
rect 100668 9696 100720 9716
rect 100720 9696 100722 9716
rect 98642 8628 98698 8664
rect 98642 8608 98644 8628
rect 98644 8608 98696 8628
rect 98696 8608 98698 8628
rect 99286 8200 99342 8256
rect 99470 4256 99526 4312
rect 99378 2896 99434 2952
rect 99010 2352 99066 2408
rect 99470 1808 99526 1864
rect 100298 8628 100354 8664
rect 100298 8608 100300 8628
rect 100300 8608 100352 8628
rect 100352 8608 100354 8628
rect 100114 6704 100170 6760
rect 102351 9274 102407 9276
rect 102431 9274 102487 9276
rect 102511 9274 102567 9276
rect 102591 9274 102647 9276
rect 102351 9222 102397 9274
rect 102397 9222 102407 9274
rect 102431 9222 102461 9274
rect 102461 9222 102473 9274
rect 102473 9222 102487 9274
rect 102511 9222 102525 9274
rect 102525 9222 102537 9274
rect 102537 9222 102567 9274
rect 102591 9222 102601 9274
rect 102601 9222 102647 9274
rect 102351 9220 102407 9222
rect 102431 9220 102487 9222
rect 102511 9220 102567 9222
rect 102591 9220 102647 9222
rect 102351 8186 102407 8188
rect 102431 8186 102487 8188
rect 102511 8186 102567 8188
rect 102591 8186 102647 8188
rect 102351 8134 102397 8186
rect 102397 8134 102407 8186
rect 102431 8134 102461 8186
rect 102461 8134 102473 8186
rect 102473 8134 102487 8186
rect 102511 8134 102525 8186
rect 102525 8134 102537 8186
rect 102537 8134 102567 8186
rect 102591 8134 102601 8186
rect 102601 8134 102647 8186
rect 102351 8132 102407 8134
rect 102431 8132 102487 8134
rect 102511 8132 102567 8134
rect 102591 8132 102647 8134
rect 102351 7098 102407 7100
rect 102431 7098 102487 7100
rect 102511 7098 102567 7100
rect 102591 7098 102647 7100
rect 102351 7046 102397 7098
rect 102397 7046 102407 7098
rect 102431 7046 102461 7098
rect 102461 7046 102473 7098
rect 102473 7046 102487 7098
rect 102511 7046 102525 7098
rect 102525 7046 102537 7098
rect 102537 7046 102567 7098
rect 102591 7046 102601 7098
rect 102601 7046 102647 7098
rect 102351 7044 102407 7046
rect 102431 7044 102487 7046
rect 102511 7044 102567 7046
rect 102591 7044 102647 7046
rect 100574 5752 100630 5808
rect 100574 5072 100630 5128
rect 97446 1264 97502 1320
rect 97078 720 97134 776
rect 98458 720 98514 776
rect 98734 720 98790 776
rect 96526 448 96582 504
rect 101862 6840 101918 6896
rect 102230 6568 102286 6624
rect 102351 6010 102407 6012
rect 102431 6010 102487 6012
rect 102511 6010 102567 6012
rect 102591 6010 102647 6012
rect 102351 5958 102397 6010
rect 102397 5958 102407 6010
rect 102431 5958 102461 6010
rect 102461 5958 102473 6010
rect 102473 5958 102487 6010
rect 102511 5958 102525 6010
rect 102525 5958 102537 6010
rect 102537 5958 102567 6010
rect 102591 5958 102601 6010
rect 102601 5958 102647 6010
rect 102351 5956 102407 5958
rect 102431 5956 102487 5958
rect 102511 5956 102567 5958
rect 102591 5956 102647 5958
rect 102351 4922 102407 4924
rect 102431 4922 102487 4924
rect 102511 4922 102567 4924
rect 102591 4922 102647 4924
rect 102351 4870 102397 4922
rect 102397 4870 102407 4922
rect 102431 4870 102461 4922
rect 102461 4870 102473 4922
rect 102473 4870 102487 4922
rect 102511 4870 102525 4922
rect 102525 4870 102537 4922
rect 102537 4870 102567 4922
rect 102591 4870 102601 4922
rect 102601 4870 102647 4922
rect 102351 4868 102407 4870
rect 102431 4868 102487 4870
rect 102511 4868 102567 4870
rect 102591 4868 102647 4870
rect 100850 4256 100906 4312
rect 101402 4256 101458 4312
rect 100758 2624 100814 2680
rect 101218 2372 101274 2408
rect 101218 2352 101220 2372
rect 101220 2352 101272 2372
rect 101272 2352 101274 2372
rect 100758 1536 100814 1592
rect 100574 1128 100630 1184
rect 101678 3168 101734 3224
rect 102351 3834 102407 3836
rect 102431 3834 102487 3836
rect 102511 3834 102567 3836
rect 102591 3834 102647 3836
rect 102351 3782 102397 3834
rect 102397 3782 102407 3834
rect 102431 3782 102461 3834
rect 102461 3782 102473 3834
rect 102473 3782 102487 3834
rect 102511 3782 102525 3834
rect 102525 3782 102537 3834
rect 102537 3782 102567 3834
rect 102591 3782 102601 3834
rect 102601 3782 102647 3834
rect 102351 3780 102407 3782
rect 102431 3780 102487 3782
rect 102511 3780 102567 3782
rect 102591 3780 102647 3782
rect 103886 10240 103942 10296
rect 100574 856 100630 912
rect 101310 856 101366 912
rect 100022 448 100078 504
rect 102351 2746 102407 2748
rect 102431 2746 102487 2748
rect 102511 2746 102567 2748
rect 102591 2746 102647 2748
rect 102351 2694 102397 2746
rect 102397 2694 102407 2746
rect 102431 2694 102461 2746
rect 102461 2694 102473 2746
rect 102473 2694 102487 2746
rect 102511 2694 102525 2746
rect 102525 2694 102537 2746
rect 102537 2694 102567 2746
rect 102591 2694 102601 2746
rect 102601 2694 102647 2746
rect 102351 2692 102407 2694
rect 102431 2692 102487 2694
rect 102511 2692 102567 2694
rect 102591 2692 102647 2694
rect 103426 2508 103482 2544
rect 103426 2488 103428 2508
rect 103428 2488 103480 2508
rect 103480 2488 103482 2508
rect 104898 10240 104954 10296
rect 105634 10240 105690 10296
rect 106278 10240 106334 10296
rect 107198 10240 107254 10296
rect 107750 10240 107806 10296
rect 108394 10240 108450 10296
rect 109038 10240 109094 10296
rect 110050 10240 110106 10296
rect 110786 10240 110842 10296
rect 111522 10240 111578 10296
rect 112350 10240 112406 10296
rect 112902 10240 112958 10296
rect 113546 10240 113602 10296
rect 114190 10240 114246 10296
rect 115202 10240 115258 10296
rect 115938 10240 115994 10296
rect 116674 10240 116730 10296
rect 117318 10240 117374 10296
rect 118054 10240 118110 10296
rect 118698 10240 118754 10296
rect 119342 10240 119398 10296
rect 120354 10240 120410 10296
rect 121090 10240 121146 10296
rect 121366 10240 121422 10296
rect 122654 10240 122710 10296
rect 123206 10240 123262 10296
rect 123942 10240 123998 10296
rect 104898 5480 104954 5536
rect 103794 2216 103850 2272
rect 102351 1658 102407 1660
rect 102431 1658 102487 1660
rect 102511 1658 102567 1660
rect 102591 1658 102647 1660
rect 102351 1606 102397 1658
rect 102397 1606 102407 1658
rect 102431 1606 102461 1658
rect 102461 1606 102473 1658
rect 102473 1606 102487 1658
rect 102511 1606 102525 1658
rect 102525 1606 102537 1658
rect 102537 1606 102567 1658
rect 102591 1606 102601 1658
rect 102601 1606 102647 1658
rect 102351 1604 102407 1606
rect 102431 1604 102487 1606
rect 102511 1604 102567 1606
rect 102591 1604 102647 1606
rect 104622 1264 104678 1320
rect 105450 1808 105506 1864
rect 103242 448 103298 504
rect 103886 448 103942 504
rect 104714 448 104770 504
rect 105634 448 105690 504
rect 106186 448 106242 504
rect 106830 1128 106886 1184
rect 108670 6160 108726 6216
rect 108854 5772 108910 5808
rect 108854 5752 108856 5772
rect 108856 5752 108908 5772
rect 108908 5752 108910 5772
rect 108394 5208 108450 5264
rect 109038 3440 109094 3496
rect 109406 5344 109462 5400
rect 112350 7384 112406 7440
rect 111522 5788 111524 5808
rect 111524 5788 111576 5808
rect 111576 5788 111578 5808
rect 111522 5752 111578 5788
rect 110510 3984 110566 4040
rect 112718 6316 112774 6352
rect 112718 6296 112720 6316
rect 112720 6296 112772 6316
rect 112772 6296 112774 6316
rect 112534 3032 112590 3088
rect 113178 6704 113234 6760
rect 113362 4428 113364 4448
rect 113364 4428 113416 4448
rect 113416 4428 113418 4448
rect 113362 4392 113418 4428
rect 114834 7928 114890 7984
rect 114742 7792 114798 7848
rect 107106 448 107162 504
rect 107750 448 107806 504
rect 108394 448 108450 504
rect 109038 448 109094 504
rect 110050 448 110106 504
rect 110786 448 110842 504
rect 111522 448 111578 504
rect 112258 448 112314 504
rect 112902 448 112958 504
rect 115938 6432 115994 6488
rect 116214 4528 116270 4584
rect 115754 2916 115810 2952
rect 115754 2896 115756 2916
rect 115756 2896 115808 2916
rect 115808 2896 115810 2916
rect 116122 3576 116178 3632
rect 117410 5480 117466 5536
rect 117318 1400 117374 1456
rect 118974 7656 119030 7712
rect 117594 720 117650 776
rect 119434 5636 119490 5672
rect 119434 5616 119436 5636
rect 119436 5616 119488 5636
rect 119488 5616 119490 5636
rect 120354 7520 120410 7576
rect 118422 992 118478 1048
rect 119986 3884 119988 3904
rect 119988 3884 120040 3904
rect 120040 3884 120042 3904
rect 119986 3848 120042 3884
rect 119342 2080 119398 2136
rect 120354 3596 120410 3632
rect 120354 3576 120356 3596
rect 120356 3576 120408 3596
rect 120408 3576 120410 3596
rect 114190 584 114246 640
rect 115202 584 115258 640
rect 115754 584 115810 640
rect 116674 584 116730 640
rect 118054 584 118110 640
rect 118698 584 118754 640
rect 119342 584 119398 640
rect 120354 584 120410 640
rect 120630 3304 120686 3360
rect 122194 5228 122250 5264
rect 122194 5208 122196 5228
rect 122196 5208 122248 5228
rect 122248 5208 122250 5228
rect 121642 1556 121698 1592
rect 121642 1536 121644 1556
rect 121644 1536 121696 1556
rect 121696 1536 121698 1556
rect 120906 856 120962 912
rect 125322 10376 125378 10432
rect 127806 10376 127862 10432
rect 125230 10240 125286 10296
rect 126334 10240 126390 10296
rect 126794 10240 126850 10296
rect 123298 1944 123354 2000
rect 121090 584 121146 640
rect 121826 584 121882 640
rect 122654 584 122710 640
rect 123114 584 123170 640
rect 123942 584 123998 640
rect 127898 10240 127954 10296
rect 128818 10240 128874 10296
rect 129646 10240 129702 10296
rect 130474 10240 130530 10296
rect 131486 10240 131542 10296
rect 132314 10240 132370 10296
rect 130290 7384 130346 7440
rect 128358 1400 128414 1456
rect 130198 5888 130254 5944
rect 124770 584 124826 640
rect 125322 584 125378 640
rect 126334 584 126390 640
rect 126794 584 126850 640
rect 127806 584 127862 640
rect 129278 584 129334 640
rect 130014 584 130070 640
rect 120446 448 120502 504
rect 124034 448 124090 504
rect 133050 10240 133106 10296
rect 133510 10240 133566 10296
rect 148414 10376 148470 10432
rect 134246 10240 134302 10296
rect 134890 10240 134946 10296
rect 138754 10240 138810 10296
rect 143262 10240 143318 10296
rect 136149 9818 136205 9820
rect 136229 9818 136285 9820
rect 136309 9818 136365 9820
rect 136389 9818 136445 9820
rect 136149 9766 136195 9818
rect 136195 9766 136205 9818
rect 136229 9766 136259 9818
rect 136259 9766 136271 9818
rect 136271 9766 136285 9818
rect 136309 9766 136323 9818
rect 136323 9766 136335 9818
rect 136335 9766 136365 9818
rect 136389 9766 136399 9818
rect 136399 9766 136445 9818
rect 136149 9764 136205 9766
rect 136229 9764 136285 9766
rect 136309 9764 136365 9766
rect 136389 9764 136445 9766
rect 137374 9580 137430 9616
rect 138846 10104 138902 10160
rect 140686 10104 140742 10160
rect 141330 10104 141386 10160
rect 141974 10104 142030 10160
rect 139766 9832 139822 9888
rect 137374 9560 137376 9580
rect 137376 9560 137428 9580
rect 137428 9560 137430 9580
rect 136149 8730 136205 8732
rect 136229 8730 136285 8732
rect 136309 8730 136365 8732
rect 136389 8730 136445 8732
rect 136149 8678 136195 8730
rect 136195 8678 136205 8730
rect 136229 8678 136259 8730
rect 136259 8678 136271 8730
rect 136271 8678 136285 8730
rect 136309 8678 136323 8730
rect 136323 8678 136335 8730
rect 136335 8678 136365 8730
rect 136389 8678 136399 8730
rect 136399 8678 136445 8730
rect 136149 8676 136205 8678
rect 136229 8676 136285 8678
rect 136309 8676 136365 8678
rect 136389 8676 136445 8678
rect 136149 7642 136205 7644
rect 136229 7642 136285 7644
rect 136309 7642 136365 7644
rect 136389 7642 136445 7644
rect 136149 7590 136195 7642
rect 136195 7590 136205 7642
rect 136229 7590 136259 7642
rect 136259 7590 136271 7642
rect 136271 7590 136285 7642
rect 136309 7590 136323 7642
rect 136323 7590 136335 7642
rect 136335 7590 136365 7642
rect 136389 7590 136399 7642
rect 136399 7590 136445 7642
rect 136149 7588 136205 7590
rect 136229 7588 136285 7590
rect 136309 7588 136365 7590
rect 136389 7588 136445 7590
rect 136149 6554 136205 6556
rect 136229 6554 136285 6556
rect 136309 6554 136365 6556
rect 136389 6554 136445 6556
rect 136149 6502 136195 6554
rect 136195 6502 136205 6554
rect 136229 6502 136259 6554
rect 136259 6502 136271 6554
rect 136271 6502 136285 6554
rect 136309 6502 136323 6554
rect 136323 6502 136335 6554
rect 136335 6502 136365 6554
rect 136389 6502 136399 6554
rect 136399 6502 136445 6554
rect 136149 6500 136205 6502
rect 136229 6500 136285 6502
rect 136309 6500 136365 6502
rect 136389 6500 136445 6502
rect 136149 5466 136205 5468
rect 136229 5466 136285 5468
rect 136309 5466 136365 5468
rect 136389 5466 136445 5468
rect 136149 5414 136195 5466
rect 136195 5414 136205 5466
rect 136229 5414 136259 5466
rect 136259 5414 136271 5466
rect 136271 5414 136285 5466
rect 136309 5414 136323 5466
rect 136323 5414 136335 5466
rect 136335 5414 136365 5466
rect 136389 5414 136399 5466
rect 136399 5414 136445 5466
rect 136149 5412 136205 5414
rect 136229 5412 136285 5414
rect 136309 5412 136365 5414
rect 136389 5412 136445 5414
rect 136149 4378 136205 4380
rect 136229 4378 136285 4380
rect 136309 4378 136365 4380
rect 136389 4378 136445 4380
rect 136149 4326 136195 4378
rect 136195 4326 136205 4378
rect 136229 4326 136259 4378
rect 136259 4326 136271 4378
rect 136271 4326 136285 4378
rect 136309 4326 136323 4378
rect 136323 4326 136335 4378
rect 136335 4326 136365 4378
rect 136389 4326 136399 4378
rect 136399 4326 136445 4378
rect 136149 4324 136205 4326
rect 136229 4324 136285 4326
rect 136309 4324 136365 4326
rect 136389 4324 136445 4326
rect 136149 3290 136205 3292
rect 136229 3290 136285 3292
rect 136309 3290 136365 3292
rect 136389 3290 136445 3292
rect 136149 3238 136195 3290
rect 136195 3238 136205 3290
rect 136229 3238 136259 3290
rect 136259 3238 136271 3290
rect 136271 3238 136285 3290
rect 136309 3238 136323 3290
rect 136323 3238 136335 3290
rect 136335 3238 136365 3290
rect 136389 3238 136399 3290
rect 136399 3238 136445 3290
rect 136149 3236 136205 3238
rect 136229 3236 136285 3238
rect 136309 3236 136365 3238
rect 136389 3236 136445 3238
rect 136149 2202 136205 2204
rect 136229 2202 136285 2204
rect 136309 2202 136365 2204
rect 136389 2202 136445 2204
rect 136149 2150 136195 2202
rect 136195 2150 136205 2202
rect 136229 2150 136259 2202
rect 136259 2150 136271 2202
rect 136271 2150 136285 2202
rect 136309 2150 136323 2202
rect 136323 2150 136335 2202
rect 136335 2150 136365 2202
rect 136389 2150 136399 2202
rect 136399 2150 136445 2202
rect 136149 2148 136205 2150
rect 136229 2148 136285 2150
rect 136309 2148 136365 2150
rect 136389 2148 136445 2150
rect 135258 1400 135314 1456
rect 143354 10104 143410 10160
rect 144550 10104 144606 10160
rect 145838 10104 145894 10160
rect 146206 10104 146262 10160
rect 147126 10104 147182 10160
rect 144734 9832 144790 9888
rect 138570 2352 138626 2408
rect 138018 1436 138020 1456
rect 138020 1436 138072 1456
rect 138072 1436 138074 1456
rect 138018 1400 138074 1436
rect 136149 1114 136205 1116
rect 136229 1114 136285 1116
rect 136309 1114 136365 1116
rect 136389 1114 136445 1116
rect 136149 1062 136195 1114
rect 136195 1062 136205 1114
rect 136229 1062 136259 1114
rect 136259 1062 136271 1114
rect 136271 1062 136285 1114
rect 136309 1062 136323 1114
rect 136323 1062 136335 1114
rect 136335 1062 136365 1114
rect 136389 1062 136399 1114
rect 136399 1062 136445 1114
rect 136149 1060 136205 1062
rect 136229 1060 136285 1062
rect 136309 1060 136365 1062
rect 136389 1060 136445 1062
rect 131578 584 131634 640
rect 132130 584 132186 640
rect 132958 584 133014 640
rect 133694 584 133750 640
rect 134430 584 134486 640
rect 139030 2352 139086 2408
rect 138846 2080 138902 2136
rect 139214 1964 139270 2000
rect 140686 2896 140742 2952
rect 139214 1944 139216 1964
rect 139216 1944 139268 1964
rect 139268 1944 139270 1964
rect 140778 1300 140780 1320
rect 140780 1300 140832 1320
rect 140832 1300 140834 1320
rect 138846 720 138902 776
rect 138754 584 138810 640
rect 140778 1264 140834 1300
rect 141698 2080 141754 2136
rect 141422 1808 141478 1864
rect 141974 720 142030 776
rect 143538 5636 143594 5672
rect 143538 5616 143540 5636
rect 143540 5616 143592 5636
rect 143592 5616 143594 5636
rect 144550 7520 144606 7576
rect 144274 3576 144330 3632
rect 143722 3052 143778 3088
rect 143722 3032 143724 3052
rect 143724 3032 143776 3052
rect 143776 3032 143778 3052
rect 143170 1844 143172 1864
rect 143172 1844 143224 1864
rect 143224 1844 143226 1864
rect 143170 1808 143226 1844
rect 142986 992 143042 1048
rect 143538 720 143594 776
rect 143998 2080 144054 2136
rect 144734 3612 144736 3632
rect 144736 3612 144788 3632
rect 144788 3612 144790 3632
rect 144734 3576 144790 3612
rect 144642 2080 144698 2136
rect 144918 1400 144974 1456
rect 148506 10104 148562 10160
rect 146574 7656 146630 7712
rect 146298 5344 146354 5400
rect 144550 720 144606 776
rect 145838 720 145894 776
rect 146206 720 146262 776
rect 148138 6196 148140 6216
rect 148140 6196 148192 6216
rect 148192 6196 148194 6216
rect 148138 6160 148194 6196
rect 147034 856 147090 912
rect 149702 10104 149758 10160
rect 150990 10104 151046 10160
rect 151634 10104 151690 10160
rect 150070 9832 150126 9888
rect 150254 6024 150310 6080
rect 150530 5244 150532 5264
rect 150532 5244 150584 5264
rect 150584 5244 150586 5264
rect 150530 5208 150586 5244
rect 149794 4020 149796 4040
rect 149796 4020 149848 4040
rect 149848 4020 149850 4040
rect 149794 3984 149850 4020
rect 150070 3460 150126 3496
rect 150070 3440 150072 3460
rect 150072 3440 150124 3460
rect 150124 3440 150126 3460
rect 149150 2508 149206 2544
rect 149150 2488 149152 2508
rect 149152 2488 149204 2508
rect 149204 2488 149206 2508
rect 147126 720 147182 776
rect 142066 584 142122 640
rect 148506 720 148562 776
rect 148414 584 148470 640
rect 140686 448 140742 504
rect 150438 1808 150494 1864
rect 152278 10104 152334 10160
rect 154210 10240 154266 10296
rect 157246 10240 157302 10296
rect 153198 10104 153254 10160
rect 154578 10104 154634 10160
rect 155130 9832 155186 9888
rect 151358 7928 151414 7984
rect 151358 5208 151414 5264
rect 150070 992 150126 1048
rect 149702 720 149758 776
rect 150990 720 151046 776
rect 151634 4392 151690 4448
rect 152646 6568 152702 6624
rect 152646 6332 152648 6352
rect 152648 6332 152700 6352
rect 152700 6332 152702 6352
rect 152646 6296 152702 6332
rect 154118 7792 154174 7848
rect 152002 4528 152058 4584
rect 153106 1672 153162 1728
rect 151726 992 151782 1048
rect 151634 720 151690 776
rect 152278 720 152334 776
rect 153198 720 153254 776
rect 154210 584 154266 640
rect 155958 9716 156014 9752
rect 155958 9696 155960 9716
rect 155960 9696 156012 9716
rect 156012 9696 156014 9716
rect 155038 3304 155094 3360
rect 155130 2624 155186 2680
rect 155682 2216 155738 2272
rect 155774 1536 155830 1592
rect 155222 1264 155278 1320
rect 156878 9716 156934 9752
rect 156878 9696 156880 9716
rect 156880 9696 156932 9716
rect 156932 9696 156934 9716
rect 157982 9716 158038 9752
rect 157982 9696 157984 9716
rect 157984 9696 158036 9716
rect 158036 9696 158038 9716
rect 156050 6704 156106 6760
rect 156050 3168 156106 3224
rect 155958 1400 156014 1456
rect 156418 2488 156474 2544
rect 156694 3596 156750 3632
rect 156694 3576 156696 3596
rect 156696 3576 156748 3596
rect 156748 3576 156750 3596
rect 156602 3168 156658 3224
rect 157062 3168 157118 3224
rect 157246 2760 157302 2816
rect 156786 2488 156842 2544
rect 159454 9716 159510 9752
rect 159454 9696 159456 9716
rect 159456 9696 159508 9716
rect 159508 9696 159510 9716
rect 159454 9444 159510 9480
rect 159454 9424 159456 9444
rect 159456 9424 159508 9444
rect 159508 9424 159510 9444
rect 158626 5208 158682 5264
rect 156602 1264 156658 1320
rect 156878 1536 156934 1592
rect 157430 1400 157486 1456
rect 157890 1400 157946 1456
rect 154578 720 154634 776
rect 156786 720 156842 776
rect 158534 2624 158590 2680
rect 160282 8336 160338 8392
rect 160558 5208 160614 5264
rect 159914 3848 159970 3904
rect 160834 4548 160890 4584
rect 160834 4528 160836 4548
rect 160836 4528 160888 4548
rect 160888 4528 160890 4548
rect 160006 3032 160062 3088
rect 160006 2760 160062 2816
rect 158810 584 158866 640
rect 158626 448 158682 504
rect 90822 312 90878 368
rect 91742 312 91798 368
rect 93030 312 93086 368
rect 98734 312 98790 368
rect 113546 312 113602 368
rect 130842 312 130898 368
rect 161294 8336 161350 8392
rect 162306 8472 162362 8528
rect 162122 5092 162178 5128
rect 162122 5072 162124 5092
rect 162124 5072 162176 5092
rect 162176 5072 162178 5092
rect 161662 3576 161718 3632
rect 161938 2352 161994 2408
rect 160926 1128 160982 1184
rect 162582 8336 162638 8392
rect 162766 6296 162822 6352
rect 163134 5072 163190 5128
rect 161754 1128 161810 1184
rect 161294 584 161350 640
rect 162490 584 162546 640
rect 163870 9716 163926 9752
rect 163870 9696 163872 9716
rect 163872 9696 163924 9716
rect 163924 9696 163926 9716
rect 164054 8336 164110 8392
rect 163686 7248 163742 7304
rect 163594 2488 163650 2544
rect 163410 2352 163466 2408
rect 163410 1944 163466 2000
rect 164790 8336 164846 8392
rect 165526 8336 165582 8392
rect 164238 1400 164294 1456
rect 163870 1128 163926 1184
rect 166354 8336 166410 8392
rect 166814 8200 166870 8256
rect 181810 10376 181866 10432
rect 171690 10240 171746 10296
rect 172334 10240 172390 10296
rect 167826 8336 167882 8392
rect 168378 8084 168434 8120
rect 168378 8064 168380 8084
rect 168380 8064 168432 8084
rect 168432 8064 168434 8084
rect 169022 9172 169078 9208
rect 169022 9152 169024 9172
rect 169024 9152 169076 9172
rect 169076 9152 169078 9172
rect 169948 9274 170004 9276
rect 170028 9274 170084 9276
rect 170108 9274 170164 9276
rect 170188 9274 170244 9276
rect 169948 9222 169994 9274
rect 169994 9222 170004 9274
rect 170028 9222 170058 9274
rect 170058 9222 170070 9274
rect 170070 9222 170084 9274
rect 170108 9222 170122 9274
rect 170122 9222 170134 9274
rect 170134 9222 170164 9274
rect 170188 9222 170198 9274
rect 170198 9222 170244 9274
rect 169948 9220 170004 9222
rect 170028 9220 170084 9222
rect 170108 9220 170164 9222
rect 170188 9220 170244 9222
rect 173070 10240 173126 10296
rect 173714 10240 173770 10296
rect 174450 10240 174506 10296
rect 175186 10240 175242 10296
rect 175922 10240 175978 10296
rect 176750 10240 176806 10296
rect 177486 10240 177542 10296
rect 177946 10240 178002 10296
rect 179142 10240 179198 10296
rect 179602 10240 179658 10296
rect 180338 10240 180394 10296
rect 181718 10240 181774 10296
rect 169948 8186 170004 8188
rect 170028 8186 170084 8188
rect 170108 8186 170164 8188
rect 170188 8186 170244 8188
rect 169948 8134 169994 8186
rect 169994 8134 170004 8186
rect 170028 8134 170058 8186
rect 170058 8134 170070 8186
rect 170070 8134 170084 8186
rect 170108 8134 170122 8186
rect 170122 8134 170134 8186
rect 170134 8134 170164 8186
rect 170188 8134 170198 8186
rect 170198 8134 170244 8186
rect 169948 8132 170004 8134
rect 170028 8132 170084 8134
rect 170108 8132 170164 8134
rect 170188 8132 170244 8134
rect 169948 7098 170004 7100
rect 170028 7098 170084 7100
rect 170108 7098 170164 7100
rect 170188 7098 170244 7100
rect 169948 7046 169994 7098
rect 169994 7046 170004 7098
rect 170028 7046 170058 7098
rect 170058 7046 170070 7098
rect 170070 7046 170084 7098
rect 170108 7046 170122 7098
rect 170122 7046 170134 7098
rect 170134 7046 170164 7098
rect 170188 7046 170198 7098
rect 170198 7046 170244 7098
rect 169948 7044 170004 7046
rect 170028 7044 170084 7046
rect 170108 7044 170164 7046
rect 170188 7044 170244 7046
rect 170586 6296 170642 6352
rect 169948 6010 170004 6012
rect 170028 6010 170084 6012
rect 170108 6010 170164 6012
rect 170188 6010 170244 6012
rect 169948 5958 169994 6010
rect 169994 5958 170004 6010
rect 170028 5958 170058 6010
rect 170058 5958 170070 6010
rect 170070 5958 170084 6010
rect 170108 5958 170122 6010
rect 170122 5958 170134 6010
rect 170134 5958 170164 6010
rect 170188 5958 170198 6010
rect 170198 5958 170244 6010
rect 169948 5956 170004 5958
rect 170028 5956 170084 5958
rect 170108 5956 170164 5958
rect 170188 5956 170244 5958
rect 170586 5752 170642 5808
rect 169948 4922 170004 4924
rect 170028 4922 170084 4924
rect 170108 4922 170164 4924
rect 170188 4922 170244 4924
rect 169948 4870 169994 4922
rect 169994 4870 170004 4922
rect 170028 4870 170058 4922
rect 170058 4870 170070 4922
rect 170070 4870 170084 4922
rect 170108 4870 170122 4922
rect 170122 4870 170134 4922
rect 170134 4870 170164 4922
rect 170188 4870 170198 4922
rect 170198 4870 170244 4922
rect 169948 4868 170004 4870
rect 170028 4868 170084 4870
rect 170108 4868 170164 4870
rect 170188 4868 170244 4870
rect 169948 3834 170004 3836
rect 170028 3834 170084 3836
rect 170108 3834 170164 3836
rect 170188 3834 170244 3836
rect 169948 3782 169994 3834
rect 169994 3782 170004 3834
rect 170028 3782 170058 3834
rect 170058 3782 170070 3834
rect 170070 3782 170084 3834
rect 170108 3782 170122 3834
rect 170122 3782 170134 3834
rect 170134 3782 170164 3834
rect 170188 3782 170198 3834
rect 170198 3782 170244 3834
rect 169948 3780 170004 3782
rect 170028 3780 170084 3782
rect 170108 3780 170164 3782
rect 170188 3780 170244 3782
rect 173438 7928 173494 7984
rect 173806 4392 173862 4448
rect 169948 2746 170004 2748
rect 170028 2746 170084 2748
rect 170108 2746 170164 2748
rect 170188 2746 170244 2748
rect 169948 2694 169994 2746
rect 169994 2694 170004 2746
rect 170028 2694 170058 2746
rect 170058 2694 170070 2746
rect 170070 2694 170084 2746
rect 170108 2694 170122 2746
rect 170122 2694 170134 2746
rect 170134 2694 170164 2746
rect 170188 2694 170198 2746
rect 170198 2694 170244 2746
rect 169948 2692 170004 2694
rect 170028 2692 170084 2694
rect 170108 2692 170164 2694
rect 170188 2692 170244 2694
rect 173254 2352 173310 2408
rect 176842 7520 176898 7576
rect 177026 6296 177082 6352
rect 177946 7792 178002 7848
rect 178038 7656 178094 7712
rect 177946 7112 178002 7168
rect 177946 6568 178002 6624
rect 177578 5344 177634 5400
rect 174174 3304 174230 3360
rect 169948 1658 170004 1660
rect 170028 1658 170084 1660
rect 170108 1658 170164 1660
rect 170188 1658 170244 1660
rect 169948 1606 169994 1658
rect 169994 1606 170004 1658
rect 170028 1606 170058 1658
rect 170058 1606 170070 1658
rect 170070 1606 170084 1658
rect 170108 1606 170122 1658
rect 170122 1606 170134 1658
rect 170134 1606 170164 1658
rect 170188 1606 170198 1658
rect 170198 1606 170244 1658
rect 169948 1604 170004 1606
rect 170028 1604 170084 1606
rect 170108 1604 170164 1606
rect 170188 1604 170244 1606
rect 168378 1400 168434 1456
rect 169298 1264 169354 1320
rect 165342 1128 165398 1184
rect 166078 1128 166134 1184
rect 166814 1128 166870 1184
rect 171414 1128 171470 1184
rect 171414 856 171470 912
rect 171690 856 171746 912
rect 172242 856 172298 912
rect 169298 720 169354 776
rect 164698 584 164754 640
rect 168010 584 168066 640
rect 169022 584 169078 640
rect 191286 10376 191342 10432
rect 182546 10240 182602 10296
rect 183282 10240 183338 10296
rect 184294 10240 184350 10296
rect 184754 10240 184810 10296
rect 185490 10240 185546 10296
rect 186226 10240 186282 10296
rect 186962 10240 187018 10296
rect 187698 10240 187754 10296
rect 188434 10240 188490 10296
rect 189446 10240 189502 10296
rect 189906 10240 189962 10296
rect 187698 8064 187754 8120
rect 180062 6432 180118 6488
rect 182086 6024 182142 6080
rect 182914 6160 182970 6216
rect 188434 5888 188490 5944
rect 175922 4120 175978 4176
rect 176842 2080 176898 2136
rect 176658 1264 176714 1320
rect 172978 856 173034 912
rect 173806 856 173862 912
rect 174450 856 174506 912
rect 175186 856 175242 912
rect 176566 856 176622 912
rect 177854 856 177910 912
rect 178406 856 178462 912
rect 179142 856 179198 912
rect 182546 4664 182602 4720
rect 179602 1264 179658 1320
rect 180522 856 180578 912
rect 160098 312 160154 368
rect 163318 312 163374 368
rect 87050 176 87106 232
rect 190366 2760 190422 2816
rect 186318 2488 186374 2544
rect 185030 2216 185086 2272
rect 181994 1808 182050 1864
rect 181902 1264 181958 1320
rect 181902 1164 181904 1184
rect 181904 1164 181956 1184
rect 181956 1164 181958 1184
rect 181902 1128 181958 1164
rect 183282 992 183338 1048
rect 181810 856 181866 912
rect 182546 856 182602 912
rect 184570 1128 184626 1184
rect 186318 1400 186374 1456
rect 190826 2352 190882 2408
rect 184754 992 184810 1048
rect 186962 1264 187018 1320
rect 184294 856 184350 912
rect 185582 856 185638 912
rect 188158 992 188214 1048
rect 191378 10240 191434 10296
rect 194230 10376 194286 10432
rect 192574 10240 192630 10296
rect 192850 10240 192906 10296
rect 193310 9016 193366 9072
rect 191746 2760 191802 2816
rect 191102 1536 191158 1592
rect 189446 992 189502 1048
rect 188526 856 188582 912
rect 194322 10240 194378 10296
rect 195610 10240 195666 10296
rect 195794 10240 195850 10296
rect 196530 10240 196586 10296
rect 194414 7928 194470 7984
rect 208306 10512 208362 10568
rect 199474 10376 199530 10432
rect 200946 10376 201002 10432
rect 202602 10376 202658 10432
rect 197266 10240 197322 10296
rect 198002 10240 198058 10296
rect 197174 7792 197230 7848
rect 194690 1400 194746 1456
rect 195978 1400 196034 1456
rect 198186 9016 198242 9072
rect 200026 10240 200082 10296
rect 200854 10240 200910 10296
rect 191286 1128 191342 1184
rect 202510 10240 202566 10296
rect 199934 1264 199990 1320
rect 198554 1128 198610 1184
rect 204074 10240 204130 10296
rect 203746 9818 203802 9820
rect 203826 9818 203882 9820
rect 203906 9818 203962 9820
rect 203986 9818 204042 9820
rect 203746 9766 203792 9818
rect 203792 9766 203802 9818
rect 203826 9766 203856 9818
rect 203856 9766 203868 9818
rect 203868 9766 203882 9818
rect 203906 9766 203920 9818
rect 203920 9766 203932 9818
rect 203932 9766 203962 9818
rect 203986 9766 203996 9818
rect 203996 9766 204042 9818
rect 203746 9764 203802 9766
rect 203826 9764 203882 9766
rect 203906 9764 203962 9766
rect 203986 9764 204042 9766
rect 206558 10104 206614 10160
rect 207662 10104 207718 10160
rect 205822 9580 205878 9616
rect 210882 10376 210938 10432
rect 211710 10376 211766 10432
rect 205822 9560 205824 9580
rect 205824 9560 205876 9580
rect 205876 9560 205878 9580
rect 203746 8730 203802 8732
rect 203826 8730 203882 8732
rect 203906 8730 203962 8732
rect 203986 8730 204042 8732
rect 203746 8678 203792 8730
rect 203792 8678 203802 8730
rect 203826 8678 203856 8730
rect 203856 8678 203868 8730
rect 203868 8678 203882 8730
rect 203906 8678 203920 8730
rect 203920 8678 203932 8730
rect 203932 8678 203962 8730
rect 203986 8678 203996 8730
rect 203996 8678 204042 8730
rect 203746 8676 203802 8678
rect 203826 8676 203882 8678
rect 203906 8676 203962 8678
rect 203986 8676 204042 8678
rect 203746 7642 203802 7644
rect 203826 7642 203882 7644
rect 203906 7642 203962 7644
rect 203986 7642 204042 7644
rect 203746 7590 203792 7642
rect 203792 7590 203802 7642
rect 203826 7590 203856 7642
rect 203856 7590 203868 7642
rect 203868 7590 203882 7642
rect 203906 7590 203920 7642
rect 203920 7590 203932 7642
rect 203932 7590 203962 7642
rect 203986 7590 203996 7642
rect 203996 7590 204042 7642
rect 203746 7588 203802 7590
rect 203826 7588 203882 7590
rect 203906 7588 203962 7590
rect 203986 7588 204042 7590
rect 203746 6554 203802 6556
rect 203826 6554 203882 6556
rect 203906 6554 203962 6556
rect 203986 6554 204042 6556
rect 203746 6502 203792 6554
rect 203792 6502 203802 6554
rect 203826 6502 203856 6554
rect 203856 6502 203868 6554
rect 203868 6502 203882 6554
rect 203906 6502 203920 6554
rect 203920 6502 203932 6554
rect 203932 6502 203962 6554
rect 203986 6502 203996 6554
rect 203996 6502 204042 6554
rect 203746 6500 203802 6502
rect 203826 6500 203882 6502
rect 203906 6500 203962 6502
rect 203986 6500 204042 6502
rect 203746 5466 203802 5468
rect 203826 5466 203882 5468
rect 203906 5466 203962 5468
rect 203986 5466 204042 5468
rect 203746 5414 203792 5466
rect 203792 5414 203802 5466
rect 203826 5414 203856 5466
rect 203856 5414 203868 5466
rect 203868 5414 203882 5466
rect 203906 5414 203920 5466
rect 203920 5414 203932 5466
rect 203932 5414 203962 5466
rect 203986 5414 203996 5466
rect 203996 5414 204042 5466
rect 203746 5412 203802 5414
rect 203826 5412 203882 5414
rect 203906 5412 203962 5414
rect 203986 5412 204042 5414
rect 204258 4936 204314 4992
rect 203746 4378 203802 4380
rect 203826 4378 203882 4380
rect 203906 4378 203962 4380
rect 203986 4378 204042 4380
rect 203746 4326 203792 4378
rect 203792 4326 203802 4378
rect 203826 4326 203856 4378
rect 203856 4326 203868 4378
rect 203868 4326 203882 4378
rect 203906 4326 203920 4378
rect 203920 4326 203932 4378
rect 203932 4326 203962 4378
rect 203986 4326 203996 4378
rect 203996 4326 204042 4378
rect 203746 4324 203802 4326
rect 203826 4324 203882 4326
rect 203906 4324 203962 4326
rect 203986 4324 204042 4326
rect 207202 3712 207258 3768
rect 203746 3290 203802 3292
rect 203826 3290 203882 3292
rect 203906 3290 203962 3292
rect 203986 3290 204042 3292
rect 203746 3238 203792 3290
rect 203792 3238 203802 3290
rect 203826 3238 203856 3290
rect 203856 3238 203868 3290
rect 203868 3238 203882 3290
rect 203906 3238 203920 3290
rect 203920 3238 203932 3290
rect 203932 3238 203962 3290
rect 203986 3238 203996 3290
rect 203996 3238 204042 3290
rect 203746 3236 203802 3238
rect 203826 3236 203882 3238
rect 203906 3236 203962 3238
rect 203986 3236 204042 3238
rect 203798 2916 203854 2952
rect 203798 2896 203800 2916
rect 203800 2896 203852 2916
rect 203852 2896 203854 2916
rect 204442 2916 204498 2952
rect 204442 2896 204444 2916
rect 204444 2896 204496 2916
rect 204496 2896 204498 2916
rect 202786 2760 202842 2816
rect 203746 2202 203802 2204
rect 203826 2202 203882 2204
rect 203906 2202 203962 2204
rect 203986 2202 204042 2204
rect 203746 2150 203792 2202
rect 203792 2150 203802 2202
rect 203826 2150 203856 2202
rect 203856 2150 203868 2202
rect 203868 2150 203882 2202
rect 203906 2150 203920 2202
rect 203920 2150 203932 2202
rect 203932 2150 203962 2202
rect 203986 2150 203996 2202
rect 203996 2150 204042 2202
rect 203746 2148 203802 2150
rect 203826 2148 203882 2150
rect 203906 2148 203962 2150
rect 203986 2148 204042 2150
rect 202878 1536 202934 1592
rect 201406 1128 201462 1184
rect 203746 1114 203802 1116
rect 203826 1114 203882 1116
rect 203906 1114 203962 1116
rect 203986 1114 204042 1116
rect 203746 1062 203792 1114
rect 203792 1062 203802 1114
rect 203826 1062 203856 1114
rect 203856 1062 203868 1114
rect 203868 1062 203882 1114
rect 203906 1062 203920 1114
rect 203920 1062 203932 1114
rect 203932 1062 203962 1114
rect 203986 1062 203996 1114
rect 203996 1062 204042 1114
rect 203746 1060 203802 1062
rect 203826 1060 203882 1062
rect 203906 1060 203962 1062
rect 203986 1060 204042 1062
rect 192666 856 192722 912
rect 192942 856 192998 912
rect 193678 856 193734 912
rect 195794 856 195850 912
rect 196622 856 196678 912
rect 197266 856 197322 912
rect 199934 856 199990 912
rect 200670 856 200726 912
rect 203338 856 203394 912
rect 205822 856 205878 912
rect 206558 856 206614 912
rect 208950 10104 209006 10160
rect 209318 10104 209374 10160
rect 210790 10104 210846 10160
rect 208398 5616 208454 5672
rect 208674 3576 208730 3632
rect 207662 856 207718 912
rect 208306 856 208362 912
rect 211158 5888 211214 5944
rect 213458 10104 213514 10160
rect 213918 10104 213974 10160
rect 210974 3168 211030 3224
rect 210882 2760 210938 2816
rect 210422 2488 210478 2544
rect 210422 2216 210478 2272
rect 210882 992 210938 1048
rect 208950 856 209006 912
rect 209778 856 209834 912
rect 211526 1300 211528 1320
rect 211528 1300 211580 1320
rect 211580 1300 211582 1320
rect 211526 1264 211582 1300
rect 212446 6840 212502 6896
rect 212538 5652 212540 5672
rect 212540 5652 212592 5672
rect 212592 5652 212594 5672
rect 212538 5616 212594 5652
rect 227442 10784 227498 10820
rect 218610 10512 218666 10568
rect 215482 10240 215538 10296
rect 215298 10104 215354 10160
rect 213642 4120 213698 4176
rect 214010 4140 214066 4176
rect 214010 4120 214012 4140
rect 214012 4120 214064 4140
rect 214064 4120 214066 4140
rect 212354 3984 212410 4040
rect 212354 2488 212410 2544
rect 211710 992 211766 1048
rect 213550 3304 213606 3360
rect 213458 2624 213514 2680
rect 214102 3440 214158 3496
rect 213918 2896 213974 2952
rect 212262 856 212318 912
rect 213458 856 213514 912
rect 214562 6296 214618 6352
rect 214838 7656 214894 7712
rect 214654 5652 214656 5672
rect 214656 5652 214708 5672
rect 214708 5652 214710 5672
rect 214654 5616 214710 5652
rect 214562 4800 214618 4856
rect 214470 3712 214526 3768
rect 216678 10104 216734 10160
rect 217966 10104 218022 10160
rect 216862 9832 216918 9888
rect 215022 6840 215078 6896
rect 215114 5480 215170 5536
rect 215298 6976 215354 7032
rect 221830 10376 221886 10432
rect 220818 10240 220874 10296
rect 219254 10104 219310 10160
rect 220542 10104 220598 10160
rect 222014 10240 222070 10296
rect 223118 10240 223174 10296
rect 215574 7112 215630 7168
rect 215574 6704 215630 6760
rect 216310 5652 216312 5672
rect 216312 5652 216364 5672
rect 216364 5652 216366 5672
rect 216310 5616 216366 5652
rect 216218 4664 216274 4720
rect 216770 6840 216826 6896
rect 216034 4120 216090 4176
rect 216126 3848 216182 3904
rect 216494 3984 216550 4040
rect 216586 3712 216642 3768
rect 215666 2624 215722 2680
rect 215850 2624 215906 2680
rect 215758 2352 215814 2408
rect 215666 2080 215722 2136
rect 215758 1672 215814 1728
rect 213734 856 213790 912
rect 214470 856 214526 912
rect 215114 856 215170 912
rect 216310 3052 216366 3088
rect 216310 3032 216312 3052
rect 216312 3032 216364 3052
rect 216364 3032 216366 3052
rect 216770 2488 216826 2544
rect 216678 2216 216734 2272
rect 216678 1400 216734 1456
rect 217414 4700 217416 4720
rect 217416 4700 217468 4720
rect 217468 4700 217470 4720
rect 217414 4664 217470 4700
rect 217506 3848 217562 3904
rect 217138 2760 217194 2816
rect 217690 4664 217746 4720
rect 217874 2488 217930 2544
rect 216678 856 216734 912
rect 217414 856 217470 912
rect 218518 7112 218574 7168
rect 218702 7112 218758 7168
rect 218886 6740 218888 6760
rect 218888 6740 218940 6760
rect 218940 6740 218942 6760
rect 218886 6704 218942 6740
rect 218978 6196 218980 6216
rect 218980 6196 219032 6216
rect 219032 6196 219034 6216
rect 218978 6160 219034 6196
rect 218794 3712 218850 3768
rect 223302 10104 223358 10160
rect 220634 7792 220690 7848
rect 219714 7148 219716 7168
rect 219716 7148 219768 7168
rect 219768 7148 219770 7168
rect 219714 7112 219770 7148
rect 219622 6840 219678 6896
rect 220634 6840 220690 6896
rect 219990 6432 220046 6488
rect 219254 5344 219310 5400
rect 219714 4820 219770 4856
rect 219714 4800 219716 4820
rect 219716 4800 219768 4820
rect 219768 4800 219770 4820
rect 218518 1128 218574 1184
rect 218978 992 219034 1048
rect 219438 856 219494 912
rect 220082 1964 220138 2000
rect 220082 1944 220084 1964
rect 220084 1944 220136 1964
rect 220136 1944 220138 1964
rect 220542 5072 220598 5128
rect 220818 7248 220874 7304
rect 220910 7112 220966 7168
rect 220818 1400 220874 1456
rect 221370 7248 221426 7304
rect 221370 6316 221426 6352
rect 221370 6296 221372 6316
rect 221372 6296 221424 6316
rect 221424 6296 221426 6316
rect 221462 6160 221518 6216
rect 221002 1844 221004 1864
rect 221004 1844 221056 1864
rect 221056 1844 221058 1864
rect 221002 1808 221058 1844
rect 221922 7248 221978 7304
rect 222198 7248 222254 7304
rect 221738 6160 221794 6216
rect 222106 6160 222162 6216
rect 222290 5228 222346 5264
rect 222290 5208 222292 5228
rect 222292 5208 222344 5228
rect 222344 5208 222346 5228
rect 222198 3032 222254 3088
rect 222106 2080 222162 2136
rect 222750 1264 222806 1320
rect 222198 856 222254 912
rect 218886 312 218942 368
rect 219622 348 219624 368
rect 219624 348 219676 368
rect 219676 348 219678 368
rect 219622 312 219678 348
rect 222382 1128 222438 1184
rect 222382 856 222438 912
rect 222290 312 222346 368
rect 223486 9152 223542 9208
rect 224774 9424 224830 9480
rect 223946 8744 224002 8800
rect 223394 6160 223450 6216
rect 223394 4528 223450 4584
rect 224314 7792 224370 7848
rect 223854 7520 223910 7576
rect 223210 4120 223266 4176
rect 223210 3052 223266 3088
rect 223210 3032 223212 3052
rect 223212 3032 223264 3052
rect 223264 3032 223266 3052
rect 223302 2760 223358 2816
rect 223486 2624 223542 2680
rect 223854 2624 223910 2680
rect 223394 2352 223450 2408
rect 223210 2080 223266 2136
rect 223394 1536 223450 1592
rect 223578 1536 223634 1592
rect 224130 6196 224132 6216
rect 224132 6196 224184 6216
rect 224184 6196 224186 6216
rect 224130 6160 224186 6196
rect 223946 2216 224002 2272
rect 224038 1400 224094 1456
rect 224774 8356 224830 8392
rect 224774 8336 224776 8356
rect 224776 8336 224828 8356
rect 224828 8336 224830 8356
rect 224958 7520 225014 7576
rect 224866 6976 224922 7032
rect 224958 6876 224960 6896
rect 224960 6876 225012 6896
rect 225012 6876 225014 6896
rect 224958 6840 225014 6876
rect 224866 6160 224922 6216
rect 224866 4800 224922 4856
rect 224682 4256 224738 4312
rect 224866 2760 224922 2816
rect 224682 2488 224738 2544
rect 224682 2216 224738 2272
rect 224774 1672 224830 1728
rect 225234 2216 225290 2272
rect 225694 9716 225750 9752
rect 225694 9696 225696 9716
rect 225696 9696 225748 9716
rect 225748 9696 225750 9716
rect 225970 9424 226026 9480
rect 225602 8916 225604 8936
rect 225604 8916 225656 8936
rect 225656 8916 225658 8936
rect 225602 8880 225658 8916
rect 225970 8628 226026 8664
rect 225970 8608 225972 8628
rect 225972 8608 226024 8628
rect 226024 8608 226026 8628
rect 227166 8880 227222 8936
rect 231858 10784 231914 10840
rect 233698 10820 233700 10840
rect 233700 10820 233752 10840
rect 233752 10820 233754 10840
rect 228270 9424 228326 9480
rect 226706 8628 226762 8664
rect 226706 8608 226708 8628
rect 226708 8608 226760 8628
rect 226760 8608 226762 8628
rect 226338 8200 226394 8256
rect 225602 6160 225658 6216
rect 226246 6432 226302 6488
rect 226338 6160 226394 6216
rect 226338 5616 226394 5672
rect 226614 5616 226670 5672
rect 225878 4120 225934 4176
rect 226246 4548 226302 4584
rect 226246 4528 226248 4548
rect 226248 4528 226300 4548
rect 226300 4528 226302 4548
rect 226706 4120 226762 4176
rect 226246 2760 226302 2816
rect 225878 2352 225934 2408
rect 226522 2796 226524 2816
rect 226524 2796 226576 2816
rect 226576 2796 226578 2816
rect 226522 2760 226578 2796
rect 225602 1400 225658 1456
rect 227626 8084 227682 8120
rect 227626 8064 227628 8084
rect 227628 8064 227680 8084
rect 227680 8064 227682 8084
rect 227718 4800 227774 4856
rect 227442 3884 227444 3904
rect 227444 3884 227496 3904
rect 227496 3884 227498 3904
rect 227442 3848 227498 3884
rect 229834 9716 229890 9752
rect 229834 9696 229836 9716
rect 229836 9696 229888 9716
rect 229888 9696 229890 9716
rect 231582 9696 231638 9752
rect 228454 8880 228510 8936
rect 228822 8744 228878 8800
rect 228270 8628 228326 8664
rect 228270 8608 228272 8628
rect 228272 8608 228324 8628
rect 228324 8608 228326 8628
rect 228086 6024 228142 6080
rect 229098 8628 229154 8664
rect 229098 8608 229100 8628
rect 229100 8608 229152 8628
rect 229152 8608 229154 8628
rect 228270 5244 228272 5264
rect 228272 5244 228324 5264
rect 228324 5244 228326 5264
rect 228270 5208 228326 5244
rect 228178 4800 228234 4856
rect 227902 3712 227958 3768
rect 227258 1264 227314 1320
rect 224038 176 224094 232
rect 224866 312 224922 368
rect 228730 4548 228786 4584
rect 228730 4528 228732 4548
rect 228732 4528 228784 4548
rect 228784 4528 228786 4548
rect 228362 3440 228418 3496
rect 228270 1264 228326 1320
rect 229098 3848 229154 3904
rect 230110 8744 230166 8800
rect 229742 7792 229798 7848
rect 229742 7520 229798 7576
rect 233698 10784 233754 10820
rect 233514 9716 233570 9752
rect 233514 9696 233516 9716
rect 233516 9696 233568 9716
rect 233568 9696 233570 9716
rect 231950 8628 232006 8664
rect 231950 8608 231952 8628
rect 231952 8608 232004 8628
rect 232004 8608 232006 8628
rect 230846 8336 230902 8392
rect 230294 7404 230350 7440
rect 230294 7384 230296 7404
rect 230296 7384 230348 7404
rect 230348 7384 230350 7404
rect 230386 6432 230442 6488
rect 229742 4936 229798 4992
rect 229834 2216 229890 2272
rect 230294 5344 230350 5400
rect 230570 5344 230626 5400
rect 231490 6568 231546 6624
rect 231766 6568 231822 6624
rect 230754 4120 230810 4176
rect 231030 2760 231086 2816
rect 231674 5752 231730 5808
rect 228454 1128 228510 1184
rect 232318 5752 232374 5808
rect 234342 9716 234398 9752
rect 234342 9696 234344 9716
rect 234344 9696 234396 9716
rect 234396 9696 234398 9716
rect 235078 9716 235134 9752
rect 235078 9696 235080 9716
rect 235080 9696 235132 9716
rect 235132 9696 235134 9716
rect 232870 8628 232926 8664
rect 232870 8608 232872 8628
rect 232872 8608 232924 8628
rect 232924 8608 232926 8628
rect 235262 8336 235318 8392
rect 235354 5616 235410 5672
rect 235998 9172 236054 9208
rect 235998 9152 236000 9172
rect 236000 9152 236052 9172
rect 236052 9152 236054 9172
rect 236642 8628 236698 8664
rect 236642 8608 236644 8628
rect 236644 8608 236696 8628
rect 236696 8608 236698 8628
rect 235906 2760 235962 2816
rect 236090 2624 236146 2680
rect 237102 8200 237158 8256
rect 237010 7828 237012 7848
rect 237012 7828 237064 7848
rect 237064 7828 237066 7848
rect 237010 7792 237066 7828
rect 237010 6840 237066 6896
rect 237545 9274 237601 9276
rect 237625 9274 237681 9276
rect 237705 9274 237761 9276
rect 237785 9274 237841 9276
rect 237545 9222 237591 9274
rect 237591 9222 237601 9274
rect 237625 9222 237655 9274
rect 237655 9222 237667 9274
rect 237667 9222 237681 9274
rect 237705 9222 237719 9274
rect 237719 9222 237731 9274
rect 237731 9222 237761 9274
rect 237785 9222 237795 9274
rect 237795 9222 237841 9274
rect 237545 9220 237601 9222
rect 237625 9220 237681 9222
rect 237705 9220 237761 9222
rect 237785 9220 237841 9222
rect 237286 9172 237342 9208
rect 237286 9152 237288 9172
rect 237288 9152 237340 9172
rect 237340 9152 237342 9172
rect 237545 8186 237601 8188
rect 237625 8186 237681 8188
rect 237705 8186 237761 8188
rect 237785 8186 237841 8188
rect 237545 8134 237591 8186
rect 237591 8134 237601 8186
rect 237625 8134 237655 8186
rect 237655 8134 237667 8186
rect 237667 8134 237681 8186
rect 237705 8134 237719 8186
rect 237719 8134 237731 8186
rect 237731 8134 237761 8186
rect 237785 8134 237795 8186
rect 237795 8134 237841 8186
rect 237545 8132 237601 8134
rect 237625 8132 237681 8134
rect 237705 8132 237761 8134
rect 237785 8132 237841 8134
rect 237930 8064 237986 8120
rect 237654 7928 237710 7984
rect 237838 7928 237894 7984
rect 237286 7404 237342 7440
rect 237930 7792 237986 7848
rect 237286 7384 237288 7404
rect 237288 7384 237340 7404
rect 237340 7384 237342 7404
rect 237194 7112 237250 7168
rect 237545 7098 237601 7100
rect 237625 7098 237681 7100
rect 237705 7098 237761 7100
rect 237785 7098 237841 7100
rect 237545 7046 237591 7098
rect 237591 7046 237601 7098
rect 237625 7046 237655 7098
rect 237655 7046 237667 7098
rect 237667 7046 237681 7098
rect 237705 7046 237719 7098
rect 237719 7046 237731 7098
rect 237731 7046 237761 7098
rect 237785 7046 237795 7098
rect 237795 7046 237841 7098
rect 237545 7044 237601 7046
rect 237625 7044 237681 7046
rect 237705 7044 237761 7046
rect 237785 7044 237841 7046
rect 237545 6010 237601 6012
rect 237625 6010 237681 6012
rect 237705 6010 237761 6012
rect 237785 6010 237841 6012
rect 237545 5958 237591 6010
rect 237591 5958 237601 6010
rect 237625 5958 237655 6010
rect 237655 5958 237667 6010
rect 237667 5958 237681 6010
rect 237705 5958 237719 6010
rect 237719 5958 237731 6010
rect 237731 5958 237761 6010
rect 237785 5958 237795 6010
rect 237795 5958 237841 6010
rect 237545 5956 237601 5958
rect 237625 5956 237681 5958
rect 237705 5956 237761 5958
rect 237785 5956 237841 5958
rect 237010 5888 237066 5944
rect 237545 4922 237601 4924
rect 237625 4922 237681 4924
rect 237705 4922 237761 4924
rect 237785 4922 237841 4924
rect 237545 4870 237591 4922
rect 237591 4870 237601 4922
rect 237625 4870 237655 4922
rect 237655 4870 237667 4922
rect 237667 4870 237681 4922
rect 237705 4870 237719 4922
rect 237719 4870 237731 4922
rect 237731 4870 237761 4922
rect 237785 4870 237795 4922
rect 237795 4870 237841 4922
rect 237545 4868 237601 4870
rect 237625 4868 237681 4870
rect 237705 4868 237761 4870
rect 237785 4868 237841 4870
rect 237286 4820 237342 4856
rect 237286 4800 237288 4820
rect 237288 4800 237340 4820
rect 237340 4800 237342 4820
rect 235998 2216 236054 2272
rect 235722 1536 235778 1592
rect 234618 1264 234674 1320
rect 229098 312 229154 368
rect 231306 1128 231362 1184
rect 232042 1128 232098 1184
rect 232778 1128 232834 1184
rect 234618 448 234674 504
rect 234894 448 234950 504
rect 237286 1400 237342 1456
rect 237545 3834 237601 3836
rect 237625 3834 237681 3836
rect 237705 3834 237761 3836
rect 237785 3834 237841 3836
rect 237545 3782 237591 3834
rect 237591 3782 237601 3834
rect 237625 3782 237655 3834
rect 237655 3782 237667 3834
rect 237667 3782 237681 3834
rect 237705 3782 237719 3834
rect 237719 3782 237731 3834
rect 237731 3782 237761 3834
rect 237785 3782 237795 3834
rect 237795 3782 237841 3834
rect 237545 3780 237601 3782
rect 237625 3780 237681 3782
rect 237705 3780 237761 3782
rect 237785 3780 237841 3782
rect 237930 3712 237986 3768
rect 238206 3984 238262 4040
rect 238114 3576 238170 3632
rect 237838 3304 237894 3360
rect 238942 7792 238998 7848
rect 238758 7520 238814 7576
rect 239678 10240 239734 10296
rect 240230 10240 240286 10296
rect 241242 10240 241298 10296
rect 241978 10240 242034 10296
rect 242714 10240 242770 10296
rect 243450 10240 243506 10296
rect 244186 10240 244242 10296
rect 244922 10240 244978 10296
rect 246118 10240 246174 10296
rect 246394 10240 246450 10296
rect 239034 7520 239090 7576
rect 240322 5208 240378 5264
rect 240506 5208 240562 5264
rect 238666 3168 238722 3224
rect 237545 2746 237601 2748
rect 237625 2746 237681 2748
rect 237705 2746 237761 2748
rect 237785 2746 237841 2748
rect 237545 2694 237591 2746
rect 237591 2694 237601 2746
rect 237625 2694 237655 2746
rect 237655 2694 237667 2746
rect 237667 2694 237681 2746
rect 237705 2694 237719 2746
rect 237719 2694 237731 2746
rect 237731 2694 237761 2746
rect 237785 2694 237795 2746
rect 237795 2694 237841 2746
rect 237545 2692 237601 2694
rect 237625 2692 237681 2694
rect 237705 2692 237761 2694
rect 237785 2692 237841 2694
rect 240782 3984 240838 4040
rect 242990 7656 243046 7712
rect 242898 6568 242954 6624
rect 242254 4564 242256 4584
rect 242256 4564 242308 4584
rect 242308 4564 242310 4584
rect 242254 4528 242310 4564
rect 242898 4256 242954 4312
rect 242530 3884 242532 3904
rect 242532 3884 242584 3904
rect 242584 3884 242586 3904
rect 242530 3848 242586 3884
rect 241518 3304 241574 3360
rect 240506 3168 240562 3224
rect 241518 2624 241574 2680
rect 237545 1658 237601 1660
rect 237625 1658 237681 1660
rect 237705 1658 237761 1660
rect 237785 1658 237841 1660
rect 237545 1606 237591 1658
rect 237591 1606 237601 1658
rect 237625 1606 237655 1658
rect 237655 1606 237667 1658
rect 237667 1606 237681 1658
rect 237705 1606 237719 1658
rect 237719 1606 237731 1658
rect 237731 1606 237761 1658
rect 237785 1606 237795 1658
rect 237795 1606 237841 1658
rect 237545 1604 237601 1606
rect 237625 1604 237681 1606
rect 237705 1604 237761 1606
rect 237785 1604 237841 1606
rect 236734 1128 236790 1184
rect 229834 312 229890 368
rect 230846 312 230902 368
rect 233422 312 233478 368
rect 234158 312 234214 368
rect 243818 6840 243874 6896
rect 244186 4120 244242 4176
rect 243726 3712 243782 3768
rect 243818 2488 243874 2544
rect 242898 1400 242954 1456
rect 241518 1264 241574 1320
rect 247406 10240 247462 10296
rect 247866 10240 247922 10296
rect 248694 10240 248750 10296
rect 249338 10240 249394 10296
rect 250074 10240 250130 10296
rect 250810 10240 250866 10296
rect 251546 10240 251602 10296
rect 252282 10240 252338 10296
rect 253110 10240 253166 10296
rect 253846 10240 253902 10296
rect 254490 10240 254546 10296
rect 255226 10240 255282 10296
rect 248970 7248 249026 7304
rect 251454 6704 251510 6760
rect 249614 6160 249670 6216
rect 252558 6296 252614 6352
rect 251822 5752 251878 5808
rect 250626 4684 250682 4720
rect 250626 4664 250628 4684
rect 250628 4664 250680 4684
rect 250680 4664 250682 4684
rect 245014 2896 245070 2952
rect 244278 1400 244334 1456
rect 241242 448 241298 504
rect 241978 448 242034 504
rect 243450 448 243506 504
rect 252282 2624 252338 2680
rect 258354 10548 258356 10568
rect 258356 10548 258408 10568
rect 258408 10548 258410 10568
rect 258354 10512 258410 10548
rect 256422 10240 256478 10296
rect 256698 10240 256754 10296
rect 257710 10240 257766 10296
rect 255042 4256 255098 4312
rect 248418 1400 248474 1456
rect 249798 1400 249854 1456
rect 251178 1400 251234 1456
rect 248050 856 248106 912
rect 248510 1128 248566 1184
rect 250166 584 250222 640
rect 251546 584 251602 640
rect 244922 448 244978 504
rect 246118 448 246174 504
rect 246394 448 246450 504
rect 248326 448 248382 504
rect 239586 312 239642 368
rect 239954 312 240010 368
rect 240966 312 241022 368
rect 252282 584 252338 640
rect 253478 584 253534 640
rect 253846 584 253902 640
rect 255226 584 255282 640
rect 256422 584 256478 640
rect 257618 2352 257674 2408
rect 258262 10240 258318 10296
rect 258170 8336 258226 8392
rect 260286 10548 260288 10568
rect 260288 10548 260340 10568
rect 260340 10548 260342 10568
rect 258998 10240 259054 10296
rect 260010 10240 260066 10296
rect 258170 5072 258226 5128
rect 258078 2796 258080 2816
rect 258080 2796 258132 2816
rect 258132 2796 258134 2816
rect 258078 2760 258134 2796
rect 258078 856 258134 912
rect 257894 720 257950 776
rect 260286 10512 260342 10548
rect 262218 10376 262274 10432
rect 260470 10240 260526 10296
rect 261758 10240 261814 10296
rect 259274 3440 259330 3496
rect 260194 4256 260250 4312
rect 260654 5208 260710 5264
rect 260838 3476 260840 3496
rect 260840 3476 260892 3496
rect 260892 3476 260894 3496
rect 260838 3440 260894 3476
rect 262494 10240 262550 10296
rect 262310 8200 262366 8256
rect 263230 10240 263286 10296
rect 262586 8744 262642 8800
rect 262862 8336 262918 8392
rect 261482 6196 261484 6216
rect 261484 6196 261536 6216
rect 261536 6196 261538 6216
rect 261482 6160 261538 6196
rect 262494 7112 262550 7168
rect 262310 5752 262366 5808
rect 262218 3032 262274 3088
rect 256698 584 256754 640
rect 257434 584 257490 640
rect 259182 584 259238 640
rect 259918 584 259974 640
rect 260470 584 260526 640
rect 261758 584 261814 640
rect 263046 5888 263102 5944
rect 262954 5752 263010 5808
rect 263138 5636 263194 5672
rect 263138 5616 263140 5636
rect 263140 5616 263192 5636
rect 263192 5616 263194 5636
rect 263230 5208 263286 5264
rect 264426 10376 264482 10432
rect 264334 10240 264390 10296
rect 263414 6604 263416 6624
rect 263416 6604 263468 6624
rect 263468 6604 263470 6624
rect 263414 6568 263470 6604
rect 263414 6452 263470 6488
rect 263414 6432 263416 6452
rect 263416 6432 263468 6452
rect 263468 6432 263470 6452
rect 263782 7520 263838 7576
rect 264150 6704 264206 6760
rect 265714 10240 265770 10296
rect 264058 5344 264114 5400
rect 264886 4528 264942 4584
rect 265346 6840 265402 6896
rect 265806 7656 265862 7712
rect 265990 7520 266046 7576
rect 265438 3576 265494 3632
rect 265254 2760 265310 2816
rect 264978 1400 265034 1456
rect 266174 7520 266230 7576
rect 266450 8336 266506 8392
rect 265898 3168 265954 3224
rect 267646 9460 267648 9480
rect 267648 9460 267700 9480
rect 267700 9460 267702 9480
rect 267646 9424 267702 9460
rect 267094 6840 267150 6896
rect 266910 5616 266966 5672
rect 266450 4256 266506 4312
rect 266634 2624 266690 2680
rect 267278 7812 267334 7848
rect 267278 7792 267280 7812
rect 267280 7792 267332 7812
rect 267332 7792 267334 7812
rect 267278 6160 267334 6216
rect 267186 5480 267242 5536
rect 267278 5344 267334 5400
rect 267278 4392 267334 4448
rect 266818 2896 266874 2952
rect 267186 2624 267242 2680
rect 267370 3712 267426 3768
rect 268014 9152 268070 9208
rect 268474 9560 268530 9616
rect 268106 9016 268162 9072
rect 267922 8880 267978 8936
rect 267830 7792 267886 7848
rect 268014 7792 268070 7848
rect 267646 7656 267702 7712
rect 267646 7520 267702 7576
rect 267738 7268 267794 7304
rect 267738 7248 267740 7268
rect 267740 7248 267792 7268
rect 267792 7248 267794 7268
rect 268014 7420 268016 7440
rect 268016 7420 268068 7440
rect 268068 7420 268070 7440
rect 268014 7384 268070 7420
rect 268014 7284 268016 7304
rect 268016 7284 268068 7304
rect 268068 7284 268070 7304
rect 268014 7248 268070 7284
rect 268014 6976 268070 7032
rect 268106 6840 268162 6896
rect 267738 5788 267740 5808
rect 267740 5788 267792 5808
rect 267792 5788 267794 5808
rect 267738 5752 267794 5788
rect 267738 5616 267794 5672
rect 268198 6432 268254 6488
rect 268382 6296 268438 6352
rect 268198 5888 268254 5944
rect 268474 5888 268530 5944
rect 268014 5752 268070 5808
rect 267922 5616 267978 5672
rect 267738 4684 267794 4720
rect 267738 4664 267740 4684
rect 267740 4664 267792 4684
rect 267792 4664 267794 4684
rect 268106 4936 268162 4992
rect 268014 3984 268070 4040
rect 268014 3712 268070 3768
rect 267738 3576 267794 3632
rect 267922 3576 267978 3632
rect 267738 3340 267740 3360
rect 267740 3340 267792 3360
rect 267792 3340 267794 3360
rect 267738 3304 267794 3340
rect 268106 3168 268162 3224
rect 268382 5072 268438 5128
rect 269026 10004 269028 10024
rect 269028 10004 269080 10024
rect 269080 10004 269082 10024
rect 269026 9968 269082 10004
rect 268934 9288 268990 9344
rect 271343 9818 271399 9820
rect 271423 9818 271479 9820
rect 271503 9818 271559 9820
rect 271583 9818 271639 9820
rect 271343 9766 271389 9818
rect 271389 9766 271399 9818
rect 271423 9766 271453 9818
rect 271453 9766 271465 9818
rect 271465 9766 271479 9818
rect 271503 9766 271517 9818
rect 271517 9766 271529 9818
rect 271529 9766 271559 9818
rect 271583 9766 271593 9818
rect 271593 9766 271639 9818
rect 271343 9764 271399 9766
rect 271423 9764 271479 9766
rect 271503 9764 271559 9766
rect 271583 9764 271639 9766
rect 268842 8472 268898 8528
rect 268750 7928 268806 7984
rect 268750 6432 268806 6488
rect 268566 4256 268622 4312
rect 268014 2896 268070 2952
rect 268198 2760 268254 2816
rect 268474 3984 268530 4040
rect 268290 2488 268346 2544
rect 268474 2488 268530 2544
rect 268934 8064 268990 8120
rect 269026 6568 269082 6624
rect 269118 6296 269174 6352
rect 268934 6160 268990 6216
rect 269026 6060 269028 6080
rect 269028 6060 269080 6080
rect 269080 6060 269082 6080
rect 269026 6024 269082 6060
rect 268934 5480 268990 5536
rect 268842 5344 268898 5400
rect 269394 5616 269450 5672
rect 268934 5208 268990 5264
rect 268842 4800 268898 4856
rect 269578 5616 269634 5672
rect 270130 7928 270186 7984
rect 268750 2216 268806 2272
rect 267646 1672 267702 1728
rect 268842 2080 268898 2136
rect 269026 2080 269082 2136
rect 269026 1536 269082 1592
rect 268842 1400 268898 1456
rect 270590 8472 270646 8528
rect 270498 8200 270554 8256
rect 270314 8064 270370 8120
rect 270314 5752 270370 5808
rect 270590 5752 270646 5808
rect 270498 5616 270554 5672
rect 270774 3168 270830 3224
rect 270498 2796 270500 2816
rect 270500 2796 270552 2816
rect 270552 2796 270554 2816
rect 270498 2760 270554 2796
rect 270774 2760 270830 2816
rect 271786 9424 271842 9480
rect 271970 8880 272026 8936
rect 271343 8730 271399 8732
rect 271423 8730 271479 8732
rect 271503 8730 271559 8732
rect 271583 8730 271639 8732
rect 271343 8678 271389 8730
rect 271389 8678 271399 8730
rect 271423 8678 271453 8730
rect 271453 8678 271465 8730
rect 271465 8678 271479 8730
rect 271503 8678 271517 8730
rect 271517 8678 271529 8730
rect 271529 8678 271559 8730
rect 271583 8678 271593 8730
rect 271593 8678 271639 8730
rect 271343 8676 271399 8678
rect 271423 8676 271479 8678
rect 271503 8676 271559 8678
rect 271583 8676 271639 8678
rect 271234 8336 271290 8392
rect 271786 7656 271842 7712
rect 271343 7642 271399 7644
rect 271423 7642 271479 7644
rect 271503 7642 271559 7644
rect 271583 7642 271639 7644
rect 271343 7590 271389 7642
rect 271389 7590 271399 7642
rect 271423 7590 271453 7642
rect 271453 7590 271465 7642
rect 271465 7590 271479 7642
rect 271503 7590 271517 7642
rect 271517 7590 271529 7642
rect 271529 7590 271559 7642
rect 271583 7590 271593 7642
rect 271593 7590 271639 7642
rect 271343 7588 271399 7590
rect 271423 7588 271479 7590
rect 271503 7588 271559 7590
rect 271583 7588 271639 7590
rect 271142 7520 271198 7576
rect 271786 7520 271842 7576
rect 271786 7248 271842 7304
rect 271970 7284 271972 7304
rect 271972 7284 272024 7304
rect 272024 7284 272026 7304
rect 271970 7248 272026 7284
rect 271694 6704 271750 6760
rect 272062 6704 272118 6760
rect 271343 6554 271399 6556
rect 271423 6554 271479 6556
rect 271503 6554 271559 6556
rect 271583 6554 271639 6556
rect 271343 6502 271389 6554
rect 271389 6502 271399 6554
rect 271423 6502 271453 6554
rect 271453 6502 271465 6554
rect 271465 6502 271479 6554
rect 271503 6502 271517 6554
rect 271517 6502 271529 6554
rect 271529 6502 271559 6554
rect 271583 6502 271593 6554
rect 271593 6502 271639 6554
rect 271343 6500 271399 6502
rect 271423 6500 271479 6502
rect 271503 6500 271559 6502
rect 271583 6500 271639 6502
rect 271878 6568 271934 6624
rect 271786 6024 271842 6080
rect 271694 5888 271750 5944
rect 271343 5466 271399 5468
rect 271423 5466 271479 5468
rect 271503 5466 271559 5468
rect 271583 5466 271639 5468
rect 271343 5414 271389 5466
rect 271389 5414 271399 5466
rect 271423 5414 271453 5466
rect 271453 5414 271465 5466
rect 271465 5414 271479 5466
rect 271503 5414 271517 5466
rect 271517 5414 271529 5466
rect 271529 5414 271559 5466
rect 271583 5414 271593 5466
rect 271593 5414 271639 5466
rect 271343 5412 271399 5414
rect 271423 5412 271479 5414
rect 271503 5412 271559 5414
rect 271583 5412 271639 5414
rect 271142 5364 271198 5400
rect 271142 5344 271144 5364
rect 271144 5344 271196 5364
rect 271196 5344 271198 5364
rect 271142 4392 271198 4448
rect 271343 4378 271399 4380
rect 271423 4378 271479 4380
rect 271503 4378 271559 4380
rect 271583 4378 271639 4380
rect 271343 4326 271389 4378
rect 271389 4326 271399 4378
rect 271423 4326 271453 4378
rect 271453 4326 271465 4378
rect 271465 4326 271479 4378
rect 271503 4326 271517 4378
rect 271517 4326 271529 4378
rect 271529 4326 271559 4378
rect 271583 4326 271593 4378
rect 271593 4326 271639 4378
rect 271343 4324 271399 4326
rect 271423 4324 271479 4326
rect 271503 4324 271559 4326
rect 271583 4324 271639 4326
rect 271786 5480 271842 5536
rect 271786 5072 271842 5128
rect 271142 3984 271198 4040
rect 271602 3712 271658 3768
rect 271142 3304 271198 3360
rect 271343 3290 271399 3292
rect 271423 3290 271479 3292
rect 271503 3290 271559 3292
rect 271583 3290 271639 3292
rect 271343 3238 271389 3290
rect 271389 3238 271399 3290
rect 271423 3238 271453 3290
rect 271453 3238 271465 3290
rect 271465 3238 271479 3290
rect 271503 3238 271517 3290
rect 271517 3238 271529 3290
rect 271529 3238 271559 3290
rect 271583 3238 271593 3290
rect 271593 3238 271639 3290
rect 271343 3236 271399 3238
rect 271423 3236 271479 3238
rect 271503 3236 271559 3238
rect 271583 3236 271639 3238
rect 271786 3168 271842 3224
rect 271970 6296 272026 6352
rect 271970 5364 272026 5400
rect 271970 5344 271972 5364
rect 271972 5344 272024 5364
rect 272024 5344 272026 5364
rect 271970 5072 272026 5128
rect 271970 3460 272026 3496
rect 271970 3440 271972 3460
rect 271972 3440 272024 3460
rect 272024 3440 272026 3460
rect 272154 4664 272210 4720
rect 271786 2896 271842 2952
rect 271970 2896 272026 2952
rect 268750 992 268806 1048
rect 262494 584 262550 640
rect 263230 584 263286 640
rect 264334 584 264390 640
rect 265346 584 265402 640
rect 266082 584 266138 640
rect 266910 584 266966 640
rect 267646 584 267702 640
rect 268382 584 268438 640
rect 261850 448 261906 504
rect 269026 856 269082 912
rect 270314 584 270370 640
rect 270038 448 270094 504
rect 255134 312 255190 368
rect 271970 2352 272026 2408
rect 271142 2216 271198 2272
rect 271343 2202 271399 2204
rect 271423 2202 271479 2204
rect 271503 2202 271559 2204
rect 271583 2202 271639 2204
rect 271343 2150 271389 2202
rect 271389 2150 271399 2202
rect 271423 2150 271453 2202
rect 271453 2150 271465 2202
rect 271465 2150 271479 2202
rect 271503 2150 271517 2202
rect 271517 2150 271529 2202
rect 271529 2150 271559 2202
rect 271583 2150 271593 2202
rect 271593 2150 271639 2202
rect 271343 2148 271399 2150
rect 271423 2148 271479 2150
rect 271503 2148 271559 2150
rect 271583 2148 271639 2150
rect 271786 2080 271842 2136
rect 271970 1944 272026 2000
rect 272154 1980 272156 2000
rect 272156 1980 272208 2000
rect 272208 1980 272210 2000
rect 272154 1944 272210 1980
rect 271786 1128 271842 1184
rect 271343 1114 271399 1116
rect 271423 1114 271479 1116
rect 271503 1114 271559 1116
rect 271583 1114 271639 1116
rect 271343 1062 271389 1114
rect 271389 1062 271399 1114
rect 271423 1062 271453 1114
rect 271453 1062 271465 1114
rect 271465 1062 271479 1114
rect 271503 1062 271517 1114
rect 271517 1062 271529 1114
rect 271529 1062 271559 1114
rect 271583 1062 271593 1114
rect 271593 1062 271639 1114
rect 271343 1060 271399 1062
rect 271423 1060 271479 1062
rect 271503 1060 271559 1062
rect 271583 1060 271639 1062
rect 270774 312 270830 368
rect 180890 40 180946 96
rect 224774 40 224830 96
rect 224958 40 225014 96
rect 239586 40 239642 96
rect 271786 40 271842 96
<< metal3 >>
rect 227437 10842 227503 10845
rect 231853 10842 231919 10845
rect 233693 10842 233759 10845
rect 227437 10840 233759 10842
rect 227437 10784 227442 10840
rect 227498 10784 231858 10840
rect 231914 10784 233698 10840
rect 233754 10784 233759 10840
rect 227437 10782 233759 10784
rect 227437 10779 227503 10782
rect 231853 10779 231919 10782
rect 233693 10779 233759 10782
rect 9673 10572 9739 10573
rect 20713 10572 20779 10573
rect 71313 10572 71379 10573
rect 74257 10572 74323 10573
rect 84561 10572 84627 10573
rect 86769 10572 86835 10573
rect 9622 10570 9628 10572
rect 9582 10510 9628 10570
rect 9692 10568 9739 10572
rect 20662 10570 20668 10572
rect 9734 10512 9739 10568
rect 9622 10508 9628 10510
rect 9692 10508 9739 10512
rect 20622 10510 20668 10570
rect 20732 10568 20779 10572
rect 71262 10570 71268 10572
rect 20774 10512 20779 10568
rect 20662 10508 20668 10510
rect 20732 10508 20779 10512
rect 71222 10510 71268 10570
rect 71332 10568 71379 10572
rect 74206 10570 74212 10572
rect 71374 10512 71379 10568
rect 71262 10508 71268 10510
rect 71332 10508 71379 10512
rect 74166 10510 74212 10570
rect 74276 10568 74323 10572
rect 84510 10570 84516 10572
rect 74318 10512 74323 10568
rect 74206 10508 74212 10510
rect 74276 10508 74323 10512
rect 84470 10510 84516 10570
rect 84580 10568 84627 10572
rect 86718 10570 86724 10572
rect 84622 10512 84627 10568
rect 84510 10508 84516 10510
rect 84580 10508 84627 10512
rect 86678 10510 86724 10570
rect 86788 10568 86835 10572
rect 86830 10512 86835 10568
rect 86718 10508 86724 10510
rect 86788 10508 86835 10512
rect 207790 10508 207796 10572
rect 207860 10570 207866 10572
rect 208301 10570 208367 10573
rect 207860 10568 208367 10570
rect 207860 10512 208306 10568
rect 208362 10512 208367 10568
rect 207860 10510 208367 10512
rect 207860 10508 207866 10510
rect 9673 10507 9739 10508
rect 20713 10507 20779 10508
rect 71313 10507 71379 10508
rect 74257 10507 74323 10508
rect 84561 10507 84627 10508
rect 86769 10507 86835 10508
rect 208301 10507 208367 10510
rect 218094 10508 218100 10572
rect 218164 10570 218170 10572
rect 218605 10570 218671 10573
rect 218164 10568 218671 10570
rect 218164 10512 218610 10568
rect 218666 10512 218671 10568
rect 218164 10510 218671 10512
rect 218164 10508 218170 10510
rect 218605 10507 218671 10510
rect 258349 10570 258415 10573
rect 260281 10570 260347 10573
rect 258349 10568 260347 10570
rect 258349 10512 258354 10568
rect 258410 10512 260286 10568
rect 260342 10512 260347 10568
rect 258349 10510 260347 10512
rect 258349 10507 258415 10510
rect 260281 10507 260347 10510
rect 54058 10372 54064 10436
rect 54128 10434 54134 10436
rect 54661 10434 54727 10437
rect 72049 10436 72115 10437
rect 77201 10436 77267 10437
rect 82353 10436 82419 10437
rect 83825 10436 83891 10437
rect 125317 10436 125383 10437
rect 71998 10434 72004 10436
rect 54128 10432 54727 10434
rect 54128 10376 54666 10432
rect 54722 10376 54727 10432
rect 54128 10374 54727 10376
rect 71958 10374 72004 10434
rect 72068 10432 72115 10436
rect 77150 10434 77156 10436
rect 72110 10376 72115 10432
rect 54128 10372 54134 10374
rect 54661 10371 54727 10374
rect 71998 10372 72004 10374
rect 72068 10372 72115 10376
rect 77110 10374 77156 10434
rect 77220 10432 77267 10436
rect 82302 10434 82308 10436
rect 77262 10376 77267 10432
rect 77150 10372 77156 10374
rect 77220 10372 77267 10376
rect 82262 10374 82308 10434
rect 82372 10432 82419 10436
rect 83774 10434 83780 10436
rect 82414 10376 82419 10432
rect 82302 10372 82308 10374
rect 82372 10372 82419 10376
rect 83734 10374 83780 10434
rect 83844 10432 83891 10436
rect 83886 10376 83891 10432
rect 83774 10372 83780 10374
rect 83844 10372 83891 10376
rect 125266 10372 125272 10436
rect 125336 10434 125383 10436
rect 127801 10434 127867 10437
rect 128210 10434 128216 10436
rect 125336 10432 125428 10434
rect 125378 10376 125428 10432
rect 125336 10374 125428 10376
rect 127801 10432 128216 10434
rect 127801 10376 127806 10432
rect 127862 10376 128216 10432
rect 127801 10374 128216 10376
rect 125336 10372 125383 10374
rect 72049 10371 72115 10372
rect 77201 10371 77267 10372
rect 82353 10371 82419 10372
rect 83825 10371 83891 10372
rect 125317 10371 125383 10372
rect 127801 10371 127867 10374
rect 128210 10372 128216 10374
rect 128280 10372 128286 10436
rect 147622 10372 147628 10436
rect 147692 10434 147698 10436
rect 148409 10434 148475 10437
rect 181805 10436 181871 10437
rect 181754 10434 181760 10436
rect 147692 10432 148475 10434
rect 147692 10376 148414 10432
rect 148470 10376 148475 10432
rect 147692 10374 148475 10376
rect 181714 10374 181760 10434
rect 181824 10432 181871 10436
rect 181866 10376 181871 10432
rect 147692 10372 147698 10374
rect 148409 10371 148475 10374
rect 181754 10372 181760 10374
rect 181824 10372 181871 10376
rect 190586 10372 190592 10436
rect 190656 10434 190662 10436
rect 191281 10434 191347 10437
rect 190656 10432 191347 10434
rect 190656 10376 191286 10432
rect 191342 10376 191347 10432
rect 190656 10374 191347 10376
rect 190656 10372 190662 10374
rect 181805 10371 181871 10372
rect 191281 10371 191347 10374
rect 193530 10372 193536 10436
rect 193600 10434 193606 10436
rect 194225 10434 194291 10437
rect 193600 10432 194291 10434
rect 193600 10376 194230 10432
rect 194286 10376 194291 10432
rect 193600 10374 194291 10376
rect 193600 10372 193606 10374
rect 194225 10371 194291 10374
rect 198682 10372 198688 10436
rect 198752 10434 198758 10436
rect 199469 10434 199535 10437
rect 200941 10436 201007 10437
rect 198752 10432 199535 10434
rect 198752 10376 199474 10432
rect 199530 10376 199535 10432
rect 198752 10374 199535 10376
rect 198752 10372 198758 10374
rect 199469 10371 199535 10374
rect 200890 10372 200896 10436
rect 200960 10434 201007 10436
rect 200960 10432 201052 10434
rect 201002 10376 201052 10432
rect 200960 10374 201052 10376
rect 200960 10372 201007 10374
rect 202362 10372 202368 10436
rect 202432 10434 202438 10436
rect 202597 10434 202663 10437
rect 202432 10432 202663 10434
rect 202432 10376 202602 10432
rect 202658 10376 202663 10432
rect 202432 10374 202663 10376
rect 202432 10372 202438 10374
rect 200941 10371 201007 10372
rect 202597 10371 202663 10374
rect 209998 10372 210004 10436
rect 210068 10434 210074 10436
rect 210877 10434 210943 10437
rect 210068 10432 210943 10434
rect 210068 10376 210882 10432
rect 210938 10376 210943 10432
rect 210068 10374 210943 10376
rect 210068 10372 210074 10374
rect 210877 10371 210943 10374
rect 211470 10372 211476 10436
rect 211540 10434 211546 10436
rect 211705 10434 211771 10437
rect 211540 10432 211771 10434
rect 211540 10376 211710 10432
rect 211766 10376 211771 10432
rect 211540 10374 211771 10376
rect 211540 10372 211546 10374
rect 211705 10371 211771 10374
rect 221038 10372 221044 10436
rect 221108 10434 221114 10436
rect 221825 10434 221891 10437
rect 221108 10432 221891 10434
rect 221108 10376 221830 10432
rect 221886 10376 221891 10432
rect 221108 10374 221891 10376
rect 221108 10372 221114 10374
rect 221825 10371 221891 10374
rect 261058 10372 261064 10436
rect 261128 10434 261134 10436
rect 262213 10434 262279 10437
rect 261128 10432 262279 10434
rect 261128 10376 262218 10432
rect 262274 10376 262279 10432
rect 261128 10374 262279 10376
rect 261128 10372 261134 10374
rect 262213 10371 262279 10374
rect 264421 10434 264487 10437
rect 264738 10434 264744 10436
rect 264421 10432 264744 10434
rect 264421 10376 264426 10432
rect 264482 10376 264744 10432
rect 264421 10374 264744 10376
rect 264421 10371 264487 10374
rect 264738 10372 264744 10374
rect 264808 10372 264814 10436
rect 31753 10300 31819 10301
rect 31702 10298 31708 10300
rect 31666 10238 31708 10298
rect 31772 10298 31819 10300
rect 31772 10296 31864 10298
rect 31814 10240 31864 10296
rect 31702 10236 31708 10238
rect 31772 10238 31864 10240
rect 31772 10236 31819 10238
rect 34922 10236 34928 10300
rect 34992 10298 34998 10300
rect 35157 10298 35223 10301
rect 34992 10296 35223 10298
rect 34992 10240 35162 10296
rect 35218 10240 35223 10296
rect 34992 10238 35223 10240
rect 34992 10236 34998 10238
rect 31753 10235 31819 10236
rect 35157 10235 35223 10238
rect 35617 10300 35683 10301
rect 35617 10296 35664 10300
rect 35728 10298 35734 10300
rect 36261 10298 36327 10301
rect 36394 10298 36400 10300
rect 35617 10240 35622 10296
rect 35617 10236 35664 10240
rect 35728 10238 35774 10298
rect 36261 10296 36400 10298
rect 36261 10240 36266 10296
rect 36322 10240 36400 10296
rect 36261 10238 36400 10240
rect 35728 10236 35734 10238
rect 35617 10235 35683 10236
rect 36261 10235 36327 10238
rect 36394 10236 36400 10238
rect 36464 10236 36470 10300
rect 36905 10298 36971 10301
rect 37130 10298 37136 10300
rect 36905 10296 37136 10298
rect 36905 10240 36910 10296
rect 36966 10240 37136 10296
rect 36905 10238 37136 10240
rect 36905 10235 36971 10238
rect 37130 10236 37136 10238
rect 37200 10236 37206 10300
rect 37866 10236 37872 10300
rect 37936 10298 37942 10300
rect 38101 10298 38167 10301
rect 37936 10296 38167 10298
rect 37936 10240 38106 10296
rect 38162 10240 38167 10296
rect 37936 10238 38167 10240
rect 37936 10236 37942 10238
rect 38101 10235 38167 10238
rect 38602 10236 38608 10300
rect 38672 10298 38678 10300
rect 38837 10298 38903 10301
rect 38672 10296 38903 10298
rect 38672 10240 38842 10296
rect 38898 10240 38903 10296
rect 38672 10238 38903 10240
rect 38672 10236 38678 10238
rect 38837 10235 38903 10238
rect 39338 10236 39344 10300
rect 39408 10298 39414 10300
rect 39481 10298 39547 10301
rect 39408 10296 39547 10298
rect 39408 10240 39486 10296
rect 39542 10240 39547 10296
rect 39408 10238 39547 10240
rect 39408 10236 39414 10238
rect 39481 10235 39547 10238
rect 40074 10236 40080 10300
rect 40144 10298 40150 10300
rect 40309 10298 40375 10301
rect 40144 10296 40375 10298
rect 40144 10240 40314 10296
rect 40370 10240 40375 10296
rect 40144 10238 40375 10240
rect 40144 10236 40150 10238
rect 40309 10235 40375 10238
rect 40769 10300 40835 10301
rect 40769 10296 40816 10300
rect 40880 10298 40886 10300
rect 41413 10298 41479 10301
rect 41546 10298 41552 10300
rect 40769 10240 40774 10296
rect 40769 10236 40816 10240
rect 40880 10238 40926 10298
rect 41413 10296 41552 10298
rect 41413 10240 41418 10296
rect 41474 10240 41552 10296
rect 41413 10238 41552 10240
rect 40880 10236 40886 10238
rect 40769 10235 40835 10236
rect 41413 10235 41479 10238
rect 41546 10236 41552 10238
rect 41616 10236 41622 10300
rect 42057 10298 42123 10301
rect 42282 10298 42288 10300
rect 42057 10296 42288 10298
rect 42057 10240 42062 10296
rect 42118 10240 42288 10296
rect 42057 10238 42288 10240
rect 42057 10235 42123 10238
rect 42282 10236 42288 10238
rect 42352 10236 42358 10300
rect 43018 10236 43024 10300
rect 43088 10298 43094 10300
rect 43253 10298 43319 10301
rect 43088 10296 43319 10298
rect 43088 10240 43258 10296
rect 43314 10240 43319 10296
rect 43088 10238 43319 10240
rect 43088 10236 43094 10238
rect 43253 10235 43319 10238
rect 43754 10236 43760 10300
rect 43824 10298 43830 10300
rect 43989 10298 44055 10301
rect 43824 10296 44055 10298
rect 43824 10240 43994 10296
rect 44050 10240 44055 10296
rect 43824 10238 44055 10240
rect 43824 10236 43830 10238
rect 43989 10235 44055 10238
rect 44490 10236 44496 10300
rect 44560 10298 44566 10300
rect 44633 10298 44699 10301
rect 44560 10296 44699 10298
rect 44560 10240 44638 10296
rect 44694 10240 44699 10296
rect 44560 10238 44699 10240
rect 44560 10236 44566 10238
rect 44633 10235 44699 10238
rect 45226 10236 45232 10300
rect 45296 10298 45302 10300
rect 45461 10298 45527 10301
rect 45296 10296 45527 10298
rect 45296 10240 45466 10296
rect 45522 10240 45527 10296
rect 45296 10238 45527 10240
rect 45296 10236 45302 10238
rect 45461 10235 45527 10238
rect 45921 10300 45987 10301
rect 45921 10296 45968 10300
rect 46032 10298 46038 10300
rect 46565 10298 46631 10301
rect 46698 10298 46704 10300
rect 45921 10240 45926 10296
rect 45921 10236 45968 10240
rect 46032 10238 46078 10298
rect 46565 10296 46704 10298
rect 46565 10240 46570 10296
rect 46626 10240 46704 10296
rect 46565 10238 46704 10240
rect 46032 10236 46038 10238
rect 45921 10235 45987 10236
rect 46565 10235 46631 10238
rect 46698 10236 46704 10238
rect 46768 10236 46774 10300
rect 47209 10298 47275 10301
rect 48221 10300 48287 10301
rect 47434 10298 47440 10300
rect 47209 10296 47440 10298
rect 47209 10240 47214 10296
rect 47270 10240 47440 10296
rect 47209 10238 47440 10240
rect 47209 10235 47275 10238
rect 47434 10236 47440 10238
rect 47504 10236 47510 10300
rect 48170 10298 48176 10300
rect 48130 10238 48176 10298
rect 48240 10296 48287 10300
rect 48282 10240 48287 10296
rect 48170 10236 48176 10238
rect 48240 10236 48287 10240
rect 48906 10236 48912 10300
rect 48976 10298 48982 10300
rect 49141 10298 49207 10301
rect 48976 10296 49207 10298
rect 48976 10240 49146 10296
rect 49202 10240 49207 10296
rect 48976 10238 49207 10240
rect 48976 10236 48982 10238
rect 48221 10235 48287 10236
rect 49141 10235 49207 10238
rect 49642 10236 49648 10300
rect 49712 10298 49718 10300
rect 49785 10298 49851 10301
rect 49712 10296 49851 10298
rect 49712 10240 49790 10296
rect 49846 10240 49851 10296
rect 49712 10238 49851 10240
rect 49712 10236 49718 10238
rect 49785 10235 49851 10238
rect 50378 10236 50384 10300
rect 50448 10298 50454 10300
rect 50613 10298 50679 10301
rect 50448 10296 50679 10298
rect 50448 10240 50618 10296
rect 50674 10240 50679 10296
rect 50448 10238 50679 10240
rect 50448 10236 50454 10238
rect 50613 10235 50679 10238
rect 51114 10236 51120 10300
rect 51184 10298 51190 10300
rect 51349 10298 51415 10301
rect 51184 10296 51415 10298
rect 51184 10240 51354 10296
rect 51410 10240 51415 10296
rect 51184 10238 51415 10240
rect 51184 10236 51190 10238
rect 51349 10235 51415 10238
rect 51850 10236 51856 10300
rect 51920 10298 51926 10300
rect 52085 10298 52151 10301
rect 51920 10296 52151 10298
rect 51920 10240 52090 10296
rect 52146 10240 52151 10296
rect 51920 10238 52151 10240
rect 51920 10236 51926 10238
rect 52085 10235 52151 10238
rect 52586 10236 52592 10300
rect 52656 10298 52662 10300
rect 53005 10298 53071 10301
rect 52656 10296 53071 10298
rect 52656 10240 53010 10296
rect 53066 10240 53071 10296
rect 52656 10238 53071 10240
rect 52656 10236 52662 10238
rect 53005 10235 53071 10238
rect 53189 10298 53255 10301
rect 54753 10300 54819 10301
rect 55489 10300 55555 10301
rect 56225 10300 56291 10301
rect 57053 10300 57119 10301
rect 57789 10300 57855 10301
rect 53322 10298 53328 10300
rect 53189 10296 53328 10298
rect 53189 10240 53194 10296
rect 53250 10240 53328 10296
rect 53189 10238 53328 10240
rect 53189 10235 53255 10238
rect 53322 10236 53328 10238
rect 53392 10236 53398 10300
rect 54753 10298 54800 10300
rect 54708 10296 54800 10298
rect 54708 10240 54758 10296
rect 54708 10238 54800 10240
rect 54753 10236 54800 10238
rect 54864 10236 54870 10300
rect 55489 10298 55536 10300
rect 55444 10296 55536 10298
rect 55444 10240 55494 10296
rect 55444 10238 55536 10240
rect 55489 10236 55536 10238
rect 55600 10236 55606 10300
rect 56225 10298 56272 10300
rect 56180 10296 56272 10298
rect 56180 10240 56230 10296
rect 56180 10238 56272 10240
rect 56225 10236 56272 10238
rect 56336 10236 56342 10300
rect 57002 10236 57008 10300
rect 57072 10298 57119 10300
rect 57072 10296 57164 10298
rect 57114 10240 57164 10296
rect 57072 10238 57164 10240
rect 57072 10236 57119 10238
rect 57738 10236 57744 10300
rect 57808 10298 57855 10300
rect 57808 10296 57900 10298
rect 57850 10240 57900 10296
rect 57808 10238 57900 10240
rect 57808 10236 57855 10238
rect 58474 10236 58480 10300
rect 58544 10298 58550 10300
rect 58617 10298 58683 10301
rect 59261 10300 59327 10301
rect 59997 10300 60063 10301
rect 58544 10296 58683 10298
rect 58544 10240 58622 10296
rect 58678 10240 58683 10296
rect 58544 10238 58683 10240
rect 58544 10236 58550 10238
rect 54753 10235 54819 10236
rect 55489 10235 55555 10236
rect 56225 10235 56291 10236
rect 57053 10235 57119 10236
rect 57789 10235 57855 10236
rect 58617 10235 58683 10238
rect 59210 10236 59216 10300
rect 59280 10298 59327 10300
rect 59280 10296 59372 10298
rect 59322 10240 59372 10296
rect 59280 10238 59372 10240
rect 59280 10236 59327 10238
rect 59946 10236 59952 10300
rect 60016 10298 60063 10300
rect 60016 10296 60108 10298
rect 60058 10240 60108 10296
rect 60016 10238 60108 10240
rect 60016 10236 60063 10238
rect 60682 10236 60688 10300
rect 60752 10298 60758 10300
rect 60825 10298 60891 10301
rect 60752 10296 60891 10298
rect 60752 10240 60830 10296
rect 60886 10240 60891 10296
rect 60752 10238 60891 10240
rect 60752 10236 60758 10238
rect 59261 10235 59327 10236
rect 59997 10235 60063 10236
rect 60825 10235 60891 10238
rect 61418 10236 61424 10300
rect 61488 10298 61494 10300
rect 61561 10298 61627 10301
rect 61488 10296 61627 10298
rect 61488 10240 61566 10296
rect 61622 10240 61627 10296
rect 61488 10238 61627 10240
rect 61488 10236 61494 10238
rect 61561 10235 61627 10238
rect 62154 10236 62160 10300
rect 62224 10298 62230 10300
rect 62297 10298 62363 10301
rect 62224 10296 62363 10298
rect 62224 10240 62302 10296
rect 62358 10240 62363 10296
rect 62224 10238 62363 10240
rect 62224 10236 62230 10238
rect 62297 10235 62363 10238
rect 62890 10236 62896 10300
rect 62960 10298 62966 10300
rect 63401 10298 63467 10301
rect 62960 10296 63467 10298
rect 62960 10240 63406 10296
rect 63462 10240 63467 10296
rect 62960 10238 63467 10240
rect 62960 10236 62966 10238
rect 63401 10235 63467 10238
rect 63626 10236 63632 10300
rect 63696 10298 63702 10300
rect 63769 10298 63835 10301
rect 63696 10296 63835 10298
rect 63696 10240 63774 10296
rect 63830 10240 63835 10296
rect 63696 10238 63835 10240
rect 63696 10236 63702 10238
rect 63769 10235 63835 10238
rect 64362 10236 64368 10300
rect 64432 10298 64438 10300
rect 64597 10298 64663 10301
rect 64432 10296 64663 10298
rect 64432 10240 64602 10296
rect 64658 10240 64663 10296
rect 64432 10238 64663 10240
rect 64432 10236 64438 10238
rect 64597 10235 64663 10238
rect 65098 10236 65104 10300
rect 65168 10298 65174 10300
rect 65425 10298 65491 10301
rect 65168 10296 65491 10298
rect 65168 10240 65430 10296
rect 65486 10240 65491 10296
rect 65168 10238 65491 10240
rect 65168 10236 65174 10238
rect 65425 10235 65491 10238
rect 65834 10236 65840 10300
rect 65904 10298 65910 10300
rect 66161 10298 66227 10301
rect 65904 10296 66227 10298
rect 65904 10240 66166 10296
rect 66222 10240 66227 10296
rect 65904 10238 66227 10240
rect 65904 10236 65910 10238
rect 66161 10235 66227 10238
rect 66570 10236 66576 10300
rect 66640 10298 66646 10300
rect 66897 10298 66963 10301
rect 66640 10296 66963 10298
rect 66640 10240 66902 10296
rect 66958 10240 66963 10296
rect 66640 10238 66963 10240
rect 66640 10236 66646 10238
rect 66897 10235 66963 10238
rect 89662 10236 89668 10300
rect 89732 10298 89738 10300
rect 90357 10298 90423 10301
rect 103237 10300 103303 10301
rect 89732 10296 90423 10298
rect 89732 10240 90362 10296
rect 90418 10240 90423 10296
rect 89732 10238 90423 10240
rect 89732 10236 89738 10238
rect 90357 10235 90423 10238
rect 103186 10236 103192 10300
rect 103256 10298 103303 10300
rect 103881 10300 103947 10301
rect 103256 10296 103348 10298
rect 103298 10240 103348 10296
rect 103256 10238 103348 10240
rect 103881 10296 103928 10300
rect 103992 10298 103998 10300
rect 103881 10240 103886 10296
rect 103256 10236 103303 10238
rect 103237 10235 103303 10236
rect 103881 10236 103928 10240
rect 103992 10238 104038 10298
rect 103992 10236 103998 10238
rect 104658 10236 104664 10300
rect 104728 10298 104734 10300
rect 104893 10298 104959 10301
rect 104728 10296 104959 10298
rect 104728 10240 104898 10296
rect 104954 10240 104959 10296
rect 104728 10238 104959 10240
rect 104728 10236 104734 10238
rect 103881 10235 103947 10236
rect 104893 10235 104959 10238
rect 105394 10236 105400 10300
rect 105464 10298 105470 10300
rect 105629 10298 105695 10301
rect 105464 10296 105695 10298
rect 105464 10240 105634 10296
rect 105690 10240 105695 10296
rect 105464 10238 105695 10240
rect 105464 10236 105470 10238
rect 105629 10235 105695 10238
rect 106130 10236 106136 10300
rect 106200 10298 106206 10300
rect 106273 10298 106339 10301
rect 106200 10296 106339 10298
rect 106200 10240 106278 10296
rect 106334 10240 106339 10296
rect 106200 10238 106339 10240
rect 106200 10236 106206 10238
rect 106273 10235 106339 10238
rect 106866 10236 106872 10300
rect 106936 10298 106942 10300
rect 107193 10298 107259 10301
rect 106936 10296 107259 10298
rect 106936 10240 107198 10296
rect 107254 10240 107259 10296
rect 106936 10238 107259 10240
rect 106936 10236 106942 10238
rect 107193 10235 107259 10238
rect 107602 10236 107608 10300
rect 107672 10298 107678 10300
rect 107745 10298 107811 10301
rect 108389 10300 108455 10301
rect 108338 10298 108344 10300
rect 107672 10296 107811 10298
rect 107672 10240 107750 10296
rect 107806 10240 107811 10296
rect 107672 10238 107811 10240
rect 108298 10238 108344 10298
rect 108408 10296 108455 10300
rect 108450 10240 108455 10296
rect 107672 10236 107678 10238
rect 107745 10235 107811 10238
rect 108338 10236 108344 10238
rect 108408 10236 108455 10240
rect 108389 10235 108455 10236
rect 109033 10300 109099 10301
rect 109033 10296 109080 10300
rect 109144 10298 109150 10300
rect 109033 10240 109038 10296
rect 109033 10236 109080 10240
rect 109144 10238 109190 10298
rect 109144 10236 109150 10238
rect 109810 10236 109816 10300
rect 109880 10298 109886 10300
rect 110045 10298 110111 10301
rect 109880 10296 110111 10298
rect 109880 10240 110050 10296
rect 110106 10240 110111 10296
rect 109880 10238 110111 10240
rect 109880 10236 109886 10238
rect 109033 10235 109099 10236
rect 110045 10235 110111 10238
rect 110546 10236 110552 10300
rect 110616 10298 110622 10300
rect 110781 10298 110847 10301
rect 110616 10296 110847 10298
rect 110616 10240 110786 10296
rect 110842 10240 110847 10296
rect 110616 10238 110847 10240
rect 110616 10236 110622 10238
rect 110781 10235 110847 10238
rect 111282 10236 111288 10300
rect 111352 10298 111358 10300
rect 111517 10298 111583 10301
rect 111352 10296 111583 10298
rect 111352 10240 111522 10296
rect 111578 10240 111583 10296
rect 111352 10238 111583 10240
rect 111352 10236 111358 10238
rect 111517 10235 111583 10238
rect 112018 10236 112024 10300
rect 112088 10298 112094 10300
rect 112345 10298 112411 10301
rect 112088 10296 112411 10298
rect 112088 10240 112350 10296
rect 112406 10240 112411 10296
rect 112088 10238 112411 10240
rect 112088 10236 112094 10238
rect 112345 10235 112411 10238
rect 112754 10236 112760 10300
rect 112824 10298 112830 10300
rect 112897 10298 112963 10301
rect 113541 10300 113607 10301
rect 113490 10298 113496 10300
rect 112824 10296 112963 10298
rect 112824 10240 112902 10296
rect 112958 10240 112963 10296
rect 112824 10238 112963 10240
rect 113450 10238 113496 10298
rect 113560 10296 113607 10300
rect 113602 10240 113607 10296
rect 112824 10236 112830 10238
rect 112897 10235 112963 10238
rect 113490 10236 113496 10238
rect 113560 10236 113607 10240
rect 113541 10235 113607 10236
rect 114185 10300 114251 10301
rect 114185 10296 114232 10300
rect 114296 10298 114302 10300
rect 114185 10240 114190 10296
rect 114185 10236 114232 10240
rect 114296 10238 114342 10298
rect 114296 10236 114302 10238
rect 114962 10236 114968 10300
rect 115032 10298 115038 10300
rect 115197 10298 115263 10301
rect 115032 10296 115263 10298
rect 115032 10240 115202 10296
rect 115258 10240 115263 10296
rect 115032 10238 115263 10240
rect 115032 10236 115038 10238
rect 114185 10235 114251 10236
rect 115197 10235 115263 10238
rect 115698 10236 115704 10300
rect 115768 10298 115774 10300
rect 115933 10298 115999 10301
rect 115768 10296 115999 10298
rect 115768 10240 115938 10296
rect 115994 10240 115999 10296
rect 115768 10238 115999 10240
rect 115768 10236 115774 10238
rect 115933 10235 115999 10238
rect 116434 10236 116440 10300
rect 116504 10298 116510 10300
rect 116669 10298 116735 10301
rect 116504 10296 116735 10298
rect 116504 10240 116674 10296
rect 116730 10240 116735 10296
rect 116504 10238 116735 10240
rect 116504 10236 116510 10238
rect 116669 10235 116735 10238
rect 117170 10236 117176 10300
rect 117240 10298 117246 10300
rect 117313 10298 117379 10301
rect 117240 10296 117379 10298
rect 117240 10240 117318 10296
rect 117374 10240 117379 10296
rect 117240 10238 117379 10240
rect 117240 10236 117246 10238
rect 117313 10235 117379 10238
rect 117906 10236 117912 10300
rect 117976 10298 117982 10300
rect 118049 10298 118115 10301
rect 118693 10300 118759 10301
rect 117976 10296 118115 10298
rect 117976 10240 118054 10296
rect 118110 10240 118115 10296
rect 117976 10238 118115 10240
rect 117976 10236 117982 10238
rect 118049 10235 118115 10238
rect 118642 10236 118648 10300
rect 118712 10298 118759 10300
rect 119337 10300 119403 10301
rect 118712 10296 118804 10298
rect 118754 10240 118804 10296
rect 118712 10238 118804 10240
rect 119337 10296 119384 10300
rect 119448 10298 119454 10300
rect 119337 10240 119342 10296
rect 118712 10236 118759 10238
rect 118693 10235 118759 10236
rect 119337 10236 119384 10240
rect 119448 10238 119494 10298
rect 119448 10236 119454 10238
rect 120114 10236 120120 10300
rect 120184 10298 120190 10300
rect 120349 10298 120415 10301
rect 120184 10296 120415 10298
rect 120184 10240 120354 10296
rect 120410 10240 120415 10296
rect 120184 10238 120415 10240
rect 120184 10236 120190 10238
rect 119337 10235 119403 10236
rect 120349 10235 120415 10238
rect 120850 10236 120856 10300
rect 120920 10298 120926 10300
rect 121085 10298 121151 10301
rect 120920 10296 121151 10298
rect 120920 10240 121090 10296
rect 121146 10240 121151 10296
rect 120920 10238 121151 10240
rect 120920 10236 120926 10238
rect 121085 10235 121151 10238
rect 121361 10298 121427 10301
rect 121586 10298 121592 10300
rect 121361 10296 121592 10298
rect 121361 10240 121366 10296
rect 121422 10240 121592 10296
rect 121361 10238 121592 10240
rect 121361 10235 121427 10238
rect 121586 10236 121592 10238
rect 121656 10236 121662 10300
rect 122322 10236 122328 10300
rect 122392 10298 122398 10300
rect 122649 10298 122715 10301
rect 122392 10296 122715 10298
rect 122392 10240 122654 10296
rect 122710 10240 122715 10296
rect 122392 10238 122715 10240
rect 122392 10236 122398 10238
rect 122649 10235 122715 10238
rect 123058 10236 123064 10300
rect 123128 10298 123134 10300
rect 123201 10298 123267 10301
rect 123128 10296 123267 10298
rect 123128 10240 123206 10296
rect 123262 10240 123267 10296
rect 123128 10238 123267 10240
rect 123128 10236 123134 10238
rect 123201 10235 123267 10238
rect 123794 10236 123800 10300
rect 123864 10298 123870 10300
rect 123937 10298 124003 10301
rect 123864 10296 124003 10298
rect 123864 10240 123942 10296
rect 123998 10240 124003 10296
rect 123864 10238 124003 10240
rect 123864 10236 123870 10238
rect 123937 10235 124003 10238
rect 124530 10236 124536 10300
rect 124600 10298 124606 10300
rect 125225 10298 125291 10301
rect 124600 10296 125291 10298
rect 124600 10240 125230 10296
rect 125286 10240 125291 10296
rect 124600 10238 125291 10240
rect 124600 10236 124606 10238
rect 125225 10235 125291 10238
rect 126002 10236 126008 10300
rect 126072 10298 126078 10300
rect 126329 10298 126395 10301
rect 126789 10300 126855 10301
rect 126072 10296 126395 10298
rect 126072 10240 126334 10296
rect 126390 10240 126395 10296
rect 126072 10238 126395 10240
rect 126072 10236 126078 10238
rect 126329 10235 126395 10238
rect 126738 10236 126744 10300
rect 126808 10298 126855 10300
rect 126808 10296 126900 10298
rect 126850 10240 126900 10296
rect 126808 10238 126900 10240
rect 126808 10236 126855 10238
rect 127474 10236 127480 10300
rect 127544 10298 127550 10300
rect 127893 10298 127959 10301
rect 127544 10296 127959 10298
rect 127544 10240 127898 10296
rect 127954 10240 127959 10296
rect 127544 10238 127959 10240
rect 127544 10236 127550 10238
rect 126789 10235 126855 10236
rect 127893 10235 127959 10238
rect 128813 10298 128879 10301
rect 129641 10300 129707 10301
rect 130469 10300 130535 10301
rect 128946 10298 128952 10300
rect 128813 10296 128952 10298
rect 128813 10240 128818 10296
rect 128874 10240 128952 10296
rect 128813 10238 128952 10240
rect 128813 10235 128879 10238
rect 128946 10236 128952 10238
rect 129016 10236 129022 10300
rect 129641 10298 129688 10300
rect 129596 10296 129688 10298
rect 129596 10240 129646 10296
rect 129596 10238 129688 10240
rect 129641 10236 129688 10238
rect 129752 10236 129758 10300
rect 130418 10236 130424 10300
rect 130488 10298 130535 10300
rect 130488 10296 130580 10298
rect 130530 10240 130580 10296
rect 130488 10238 130580 10240
rect 130488 10236 130535 10238
rect 131154 10236 131160 10300
rect 131224 10298 131230 10300
rect 131481 10298 131547 10301
rect 131224 10296 131547 10298
rect 131224 10240 131486 10296
rect 131542 10240 131547 10296
rect 131224 10238 131547 10240
rect 131224 10236 131230 10238
rect 129641 10235 129707 10236
rect 130469 10235 130535 10236
rect 131481 10235 131547 10238
rect 131890 10236 131896 10300
rect 131960 10298 131966 10300
rect 132309 10298 132375 10301
rect 131960 10296 132375 10298
rect 131960 10240 132314 10296
rect 132370 10240 132375 10296
rect 131960 10238 132375 10240
rect 131960 10236 131966 10238
rect 132309 10235 132375 10238
rect 132626 10236 132632 10300
rect 132696 10298 132702 10300
rect 133045 10298 133111 10301
rect 132696 10296 133111 10298
rect 132696 10240 133050 10296
rect 133106 10240 133111 10296
rect 132696 10238 133111 10240
rect 132696 10236 132702 10238
rect 133045 10235 133111 10238
rect 133362 10236 133368 10300
rect 133432 10298 133438 10300
rect 133505 10298 133571 10301
rect 133432 10296 133571 10298
rect 133432 10240 133510 10296
rect 133566 10240 133571 10296
rect 133432 10238 133571 10240
rect 133432 10236 133438 10238
rect 133505 10235 133571 10238
rect 134098 10236 134104 10300
rect 134168 10298 134174 10300
rect 134241 10298 134307 10301
rect 134885 10300 134951 10301
rect 134168 10296 134307 10298
rect 134168 10240 134246 10296
rect 134302 10240 134307 10296
rect 134168 10238 134307 10240
rect 134168 10236 134174 10238
rect 134241 10235 134307 10238
rect 134834 10236 134840 10300
rect 134904 10298 134951 10300
rect 134904 10296 134996 10298
rect 134946 10240 134996 10296
rect 134904 10238 134996 10240
rect 134904 10236 134951 10238
rect 138054 10236 138060 10300
rect 138124 10298 138130 10300
rect 138749 10298 138815 10301
rect 138124 10296 138815 10298
rect 138124 10240 138754 10296
rect 138810 10240 138815 10296
rect 138124 10238 138815 10240
rect 138124 10236 138130 10238
rect 134885 10235 134951 10236
rect 138749 10235 138815 10238
rect 142470 10236 142476 10300
rect 142540 10298 142546 10300
rect 143257 10298 143323 10301
rect 142540 10296 143323 10298
rect 142540 10240 143262 10296
rect 143318 10240 143323 10296
rect 142540 10238 143323 10240
rect 142540 10236 142546 10238
rect 143257 10235 143323 10238
rect 153510 10236 153516 10300
rect 153580 10298 153586 10300
rect 154205 10298 154271 10301
rect 157241 10300 157307 10301
rect 157190 10298 157196 10300
rect 153580 10296 154271 10298
rect 153580 10240 154210 10296
rect 154266 10240 154271 10296
rect 153580 10238 154271 10240
rect 157150 10238 157196 10298
rect 157260 10296 157307 10300
rect 157302 10240 157307 10296
rect 153580 10236 153586 10238
rect 154205 10235 154271 10238
rect 157190 10236 157196 10238
rect 157260 10236 157307 10240
rect 171450 10236 171456 10300
rect 171520 10298 171526 10300
rect 171685 10298 171751 10301
rect 171520 10296 171751 10298
rect 171520 10240 171690 10296
rect 171746 10240 171751 10296
rect 171520 10238 171751 10240
rect 171520 10236 171526 10238
rect 157241 10235 157307 10236
rect 171685 10235 171751 10238
rect 172186 10236 172192 10300
rect 172256 10298 172262 10300
rect 172329 10298 172395 10301
rect 172256 10296 172395 10298
rect 172256 10240 172334 10296
rect 172390 10240 172395 10296
rect 172256 10238 172395 10240
rect 172256 10236 172262 10238
rect 172329 10235 172395 10238
rect 172922 10236 172928 10300
rect 172992 10298 172998 10300
rect 173065 10298 173131 10301
rect 173709 10300 173775 10301
rect 174445 10300 174511 10301
rect 175181 10300 175247 10301
rect 175917 10300 175983 10301
rect 173658 10298 173664 10300
rect 172992 10296 173131 10298
rect 172992 10240 173070 10296
rect 173126 10240 173131 10296
rect 172992 10238 173131 10240
rect 173618 10238 173664 10298
rect 173728 10296 173775 10300
rect 174394 10298 174400 10300
rect 173770 10240 173775 10296
rect 172992 10236 172998 10238
rect 173065 10235 173131 10238
rect 173658 10236 173664 10238
rect 173728 10236 173775 10240
rect 174354 10238 174400 10298
rect 174464 10296 174511 10300
rect 175130 10298 175136 10300
rect 174506 10240 174511 10296
rect 174394 10236 174400 10238
rect 174464 10236 174511 10240
rect 175090 10238 175136 10298
rect 175200 10296 175247 10300
rect 175866 10298 175872 10300
rect 175242 10240 175247 10296
rect 175130 10236 175136 10238
rect 175200 10236 175247 10240
rect 175826 10238 175872 10298
rect 175936 10296 175983 10300
rect 175978 10240 175983 10296
rect 175866 10236 175872 10238
rect 175936 10236 175983 10240
rect 176602 10236 176608 10300
rect 176672 10298 176678 10300
rect 176745 10298 176811 10301
rect 176672 10296 176811 10298
rect 176672 10240 176750 10296
rect 176806 10240 176811 10296
rect 176672 10238 176811 10240
rect 176672 10236 176678 10238
rect 173709 10235 173775 10236
rect 174445 10235 174511 10236
rect 175181 10235 175247 10236
rect 175917 10235 175983 10236
rect 176745 10235 176811 10238
rect 177338 10236 177344 10300
rect 177408 10298 177414 10300
rect 177481 10298 177547 10301
rect 177408 10296 177547 10298
rect 177408 10240 177486 10296
rect 177542 10240 177547 10296
rect 177408 10238 177547 10240
rect 177408 10236 177414 10238
rect 177481 10235 177547 10238
rect 177941 10298 178007 10301
rect 178074 10298 178080 10300
rect 177941 10296 178080 10298
rect 177941 10240 177946 10296
rect 178002 10240 178080 10296
rect 177941 10238 178080 10240
rect 177941 10235 178007 10238
rect 178074 10236 178080 10238
rect 178144 10236 178150 10300
rect 178810 10236 178816 10300
rect 178880 10298 178886 10300
rect 179137 10298 179203 10301
rect 179597 10300 179663 10301
rect 180333 10300 180399 10301
rect 179546 10298 179552 10300
rect 178880 10296 179203 10298
rect 178880 10240 179142 10296
rect 179198 10240 179203 10296
rect 178880 10238 179203 10240
rect 179506 10238 179552 10298
rect 179616 10296 179663 10300
rect 180282 10298 180288 10300
rect 179658 10240 179663 10296
rect 178880 10236 178886 10238
rect 179137 10235 179203 10238
rect 179546 10236 179552 10238
rect 179616 10236 179663 10240
rect 180242 10238 180288 10298
rect 180352 10296 180399 10300
rect 180394 10240 180399 10296
rect 180282 10236 180288 10238
rect 180352 10236 180399 10240
rect 181018 10236 181024 10300
rect 181088 10298 181094 10300
rect 181713 10298 181779 10301
rect 182541 10300 182607 10301
rect 183277 10300 183343 10301
rect 182490 10298 182496 10300
rect 181088 10296 181779 10298
rect 181088 10240 181718 10296
rect 181774 10240 181779 10296
rect 181088 10238 181779 10240
rect 182450 10238 182496 10298
rect 182560 10296 182607 10300
rect 183226 10298 183232 10300
rect 182602 10240 182607 10296
rect 181088 10236 181094 10238
rect 179597 10235 179663 10236
rect 180333 10235 180399 10236
rect 181713 10235 181779 10238
rect 182490 10236 182496 10238
rect 182560 10236 182607 10240
rect 183186 10238 183232 10298
rect 183296 10296 183343 10300
rect 183338 10240 183343 10296
rect 183226 10236 183232 10238
rect 183296 10236 183343 10240
rect 183962 10236 183968 10300
rect 184032 10298 184038 10300
rect 184289 10298 184355 10301
rect 184749 10300 184815 10301
rect 185485 10300 185551 10301
rect 186221 10300 186287 10301
rect 186957 10300 187023 10301
rect 187693 10300 187759 10301
rect 188429 10300 188495 10301
rect 184698 10298 184704 10300
rect 184032 10296 184355 10298
rect 184032 10240 184294 10296
rect 184350 10240 184355 10296
rect 184032 10238 184355 10240
rect 184658 10238 184704 10298
rect 184768 10296 184815 10300
rect 185434 10298 185440 10300
rect 184810 10240 184815 10296
rect 184032 10236 184038 10238
rect 182541 10235 182607 10236
rect 183277 10235 183343 10236
rect 184289 10235 184355 10238
rect 184698 10236 184704 10238
rect 184768 10236 184815 10240
rect 185394 10238 185440 10298
rect 185504 10296 185551 10300
rect 186170 10298 186176 10300
rect 185546 10240 185551 10296
rect 185434 10236 185440 10238
rect 185504 10236 185551 10240
rect 186130 10238 186176 10298
rect 186240 10296 186287 10300
rect 186906 10298 186912 10300
rect 186282 10240 186287 10296
rect 186170 10236 186176 10238
rect 186240 10236 186287 10240
rect 186866 10238 186912 10298
rect 186976 10296 187023 10300
rect 187642 10298 187648 10300
rect 187018 10240 187023 10296
rect 186906 10236 186912 10238
rect 186976 10236 187023 10240
rect 187602 10238 187648 10298
rect 187712 10296 187759 10300
rect 188378 10298 188384 10300
rect 187754 10240 187759 10296
rect 187642 10236 187648 10238
rect 187712 10236 187759 10240
rect 188338 10238 188384 10298
rect 188448 10296 188495 10300
rect 188490 10240 188495 10296
rect 188378 10236 188384 10238
rect 188448 10236 188495 10240
rect 189114 10236 189120 10300
rect 189184 10298 189190 10300
rect 189441 10298 189507 10301
rect 189901 10300 189967 10301
rect 191373 10300 191439 10301
rect 189850 10298 189856 10300
rect 189184 10296 189507 10298
rect 189184 10240 189446 10296
rect 189502 10240 189507 10296
rect 189184 10238 189507 10240
rect 189810 10238 189856 10298
rect 189920 10296 189967 10300
rect 189962 10240 189967 10296
rect 189184 10236 189190 10238
rect 184749 10235 184815 10236
rect 185485 10235 185551 10236
rect 186221 10235 186287 10236
rect 186957 10235 187023 10236
rect 187693 10235 187759 10236
rect 188429 10235 188495 10236
rect 189441 10235 189507 10238
rect 189850 10236 189856 10238
rect 189920 10236 189967 10240
rect 191322 10236 191328 10300
rect 191392 10298 191439 10300
rect 191392 10296 191484 10298
rect 191434 10240 191484 10296
rect 191392 10238 191484 10240
rect 191392 10236 191439 10238
rect 192058 10236 192064 10300
rect 192128 10298 192134 10300
rect 192569 10298 192635 10301
rect 192845 10300 192911 10301
rect 194317 10300 194383 10301
rect 192128 10296 192635 10298
rect 192128 10240 192574 10296
rect 192630 10240 192635 10296
rect 192128 10238 192635 10240
rect 192128 10236 192134 10238
rect 189901 10235 189967 10236
rect 191373 10235 191439 10236
rect 192569 10235 192635 10238
rect 192794 10236 192800 10300
rect 192864 10298 192911 10300
rect 192864 10296 192956 10298
rect 192906 10240 192956 10296
rect 192864 10238 192956 10240
rect 192864 10236 192911 10238
rect 194266 10236 194272 10300
rect 194336 10298 194383 10300
rect 194336 10296 194428 10298
rect 194378 10240 194428 10296
rect 194336 10238 194428 10240
rect 194336 10236 194383 10238
rect 195002 10236 195008 10300
rect 195072 10298 195078 10300
rect 195605 10298 195671 10301
rect 195789 10300 195855 10301
rect 196525 10300 196591 10301
rect 197261 10300 197327 10301
rect 197997 10300 198063 10301
rect 195072 10296 195671 10298
rect 195072 10240 195610 10296
rect 195666 10240 195671 10296
rect 195072 10238 195671 10240
rect 195072 10236 195078 10238
rect 192845 10235 192911 10236
rect 194317 10235 194383 10236
rect 195605 10235 195671 10238
rect 195738 10236 195744 10300
rect 195808 10298 195855 10300
rect 195808 10296 195900 10298
rect 195850 10240 195900 10296
rect 195808 10238 195900 10240
rect 195808 10236 195855 10238
rect 196474 10236 196480 10300
rect 196544 10298 196591 10300
rect 196544 10296 196636 10298
rect 196586 10240 196636 10296
rect 196544 10238 196636 10240
rect 196544 10236 196591 10238
rect 197210 10236 197216 10300
rect 197280 10298 197327 10300
rect 197280 10296 197372 10298
rect 197322 10240 197372 10296
rect 197280 10238 197372 10240
rect 197280 10236 197327 10238
rect 197946 10236 197952 10300
rect 198016 10298 198063 10300
rect 198016 10296 198108 10298
rect 198058 10240 198108 10296
rect 198016 10238 198108 10240
rect 198016 10236 198063 10238
rect 199418 10236 199424 10300
rect 199488 10298 199494 10300
rect 200021 10298 200087 10301
rect 199488 10296 200087 10298
rect 199488 10240 200026 10296
rect 200082 10240 200087 10296
rect 199488 10238 200087 10240
rect 199488 10236 199494 10238
rect 195789 10235 195855 10236
rect 196525 10235 196591 10236
rect 197261 10235 197327 10236
rect 197997 10235 198063 10236
rect 200021 10235 200087 10238
rect 200154 10236 200160 10300
rect 200224 10298 200230 10300
rect 200849 10298 200915 10301
rect 200224 10296 200915 10298
rect 200224 10240 200854 10296
rect 200910 10240 200915 10296
rect 200224 10238 200915 10240
rect 200224 10236 200230 10238
rect 200849 10235 200915 10238
rect 201626 10236 201632 10300
rect 201696 10298 201702 10300
rect 202505 10298 202571 10301
rect 201696 10296 202571 10298
rect 201696 10240 202510 10296
rect 202566 10240 202571 10296
rect 201696 10238 202571 10240
rect 201696 10236 201702 10238
rect 202505 10235 202571 10238
rect 203098 10236 203104 10300
rect 203168 10298 203174 10300
rect 204069 10298 204135 10301
rect 203168 10296 204135 10298
rect 203168 10240 204074 10296
rect 204130 10240 204135 10296
rect 203168 10238 204135 10240
rect 203168 10236 203174 10238
rect 204069 10235 204135 10238
rect 215150 10236 215156 10300
rect 215220 10298 215226 10300
rect 215477 10298 215543 10301
rect 215220 10296 215543 10298
rect 215220 10240 215482 10296
rect 215538 10240 215543 10296
rect 215220 10238 215543 10240
rect 215220 10236 215226 10238
rect 215477 10235 215543 10238
rect 220302 10236 220308 10300
rect 220372 10298 220378 10300
rect 220813 10298 220879 10301
rect 220372 10296 220879 10298
rect 220372 10240 220818 10296
rect 220874 10240 220879 10296
rect 220372 10238 220879 10240
rect 220372 10236 220378 10238
rect 220813 10235 220879 10238
rect 221774 10236 221780 10300
rect 221844 10298 221850 10300
rect 222009 10298 222075 10301
rect 221844 10296 222075 10298
rect 221844 10240 222014 10296
rect 222070 10240 222075 10296
rect 221844 10238 222075 10240
rect 221844 10236 221850 10238
rect 222009 10235 222075 10238
rect 222510 10236 222516 10300
rect 222580 10298 222586 10300
rect 223113 10298 223179 10301
rect 239673 10300 239739 10301
rect 239673 10298 239720 10300
rect 222580 10296 223179 10298
rect 222580 10240 223118 10296
rect 223174 10240 223179 10296
rect 222580 10238 223179 10240
rect 239628 10296 239720 10298
rect 239628 10240 239678 10296
rect 239628 10238 239720 10240
rect 222580 10236 222586 10238
rect 223113 10235 223179 10238
rect 239673 10236 239720 10238
rect 239784 10236 239790 10300
rect 240225 10298 240291 10301
rect 241237 10300 241303 10301
rect 241973 10300 242039 10301
rect 242709 10300 242775 10301
rect 243445 10300 243511 10301
rect 244181 10300 244247 10301
rect 244917 10300 244983 10301
rect 240450 10298 240456 10300
rect 240225 10296 240456 10298
rect 240225 10240 240230 10296
rect 240286 10240 240456 10296
rect 240225 10238 240456 10240
rect 239673 10235 239739 10236
rect 240225 10235 240291 10238
rect 240450 10236 240456 10238
rect 240520 10236 240526 10300
rect 241186 10298 241192 10300
rect 241146 10238 241192 10298
rect 241256 10296 241303 10300
rect 241922 10298 241928 10300
rect 241298 10240 241303 10296
rect 241186 10236 241192 10238
rect 241256 10236 241303 10240
rect 241882 10238 241928 10298
rect 241992 10296 242039 10300
rect 242658 10298 242664 10300
rect 242034 10240 242039 10296
rect 241922 10236 241928 10238
rect 241992 10236 242039 10240
rect 242618 10238 242664 10298
rect 242728 10296 242775 10300
rect 243394 10298 243400 10300
rect 242770 10240 242775 10296
rect 242658 10236 242664 10238
rect 242728 10236 242775 10240
rect 243354 10238 243400 10298
rect 243464 10296 243511 10300
rect 244130 10298 244136 10300
rect 243506 10240 243511 10296
rect 243394 10236 243400 10238
rect 243464 10236 243511 10240
rect 244090 10238 244136 10298
rect 244200 10296 244247 10300
rect 244866 10298 244872 10300
rect 244242 10240 244247 10296
rect 244130 10236 244136 10238
rect 244200 10236 244247 10240
rect 244826 10238 244872 10298
rect 244936 10296 244983 10300
rect 244978 10240 244983 10296
rect 244866 10236 244872 10238
rect 244936 10236 244983 10240
rect 245602 10236 245608 10300
rect 245672 10298 245678 10300
rect 246113 10298 246179 10301
rect 246389 10300 246455 10301
rect 246338 10298 246344 10300
rect 245672 10296 246179 10298
rect 245672 10240 246118 10296
rect 246174 10240 246179 10296
rect 245672 10238 246179 10240
rect 246298 10238 246344 10298
rect 246408 10296 246455 10300
rect 246450 10240 246455 10296
rect 245672 10236 245678 10238
rect 241237 10235 241303 10236
rect 241973 10235 242039 10236
rect 242709 10235 242775 10236
rect 243445 10235 243511 10236
rect 244181 10235 244247 10236
rect 244917 10235 244983 10236
rect 246113 10235 246179 10238
rect 246338 10236 246344 10238
rect 246408 10236 246455 10240
rect 247074 10236 247080 10300
rect 247144 10298 247150 10300
rect 247401 10298 247467 10301
rect 247861 10300 247927 10301
rect 247810 10298 247816 10300
rect 247144 10296 247467 10298
rect 247144 10240 247406 10296
rect 247462 10240 247467 10296
rect 247144 10238 247467 10240
rect 247770 10238 247816 10298
rect 247880 10296 247927 10300
rect 247922 10240 247927 10296
rect 247144 10236 247150 10238
rect 246389 10235 246455 10236
rect 247401 10235 247467 10238
rect 247810 10236 247816 10238
rect 247880 10236 247927 10240
rect 248546 10236 248552 10300
rect 248616 10298 248622 10300
rect 248689 10298 248755 10301
rect 249333 10300 249399 10301
rect 250069 10300 250135 10301
rect 250805 10300 250871 10301
rect 251541 10300 251607 10301
rect 252277 10300 252343 10301
rect 249282 10298 249288 10300
rect 248616 10296 248755 10298
rect 248616 10240 248694 10296
rect 248750 10240 248755 10296
rect 248616 10238 248755 10240
rect 249242 10238 249288 10298
rect 249352 10296 249399 10300
rect 250018 10298 250024 10300
rect 249394 10240 249399 10296
rect 248616 10236 248622 10238
rect 247861 10235 247927 10236
rect 248689 10235 248755 10238
rect 249282 10236 249288 10238
rect 249352 10236 249399 10240
rect 249978 10238 250024 10298
rect 250088 10296 250135 10300
rect 250754 10298 250760 10300
rect 250130 10240 250135 10296
rect 250018 10236 250024 10238
rect 250088 10236 250135 10240
rect 250714 10238 250760 10298
rect 250824 10296 250871 10300
rect 251490 10298 251496 10300
rect 250866 10240 250871 10296
rect 250754 10236 250760 10238
rect 250824 10236 250871 10240
rect 251450 10238 251496 10298
rect 251560 10296 251607 10300
rect 252226 10298 252232 10300
rect 251602 10240 251607 10296
rect 251490 10236 251496 10238
rect 251560 10236 251607 10240
rect 252186 10238 252232 10298
rect 252296 10296 252343 10300
rect 252338 10240 252343 10296
rect 252226 10236 252232 10238
rect 252296 10236 252343 10240
rect 252962 10236 252968 10300
rect 253032 10298 253038 10300
rect 253105 10298 253171 10301
rect 253032 10296 253171 10298
rect 253032 10240 253110 10296
rect 253166 10240 253171 10296
rect 253032 10238 253171 10240
rect 253032 10236 253038 10238
rect 249333 10235 249399 10236
rect 250069 10235 250135 10236
rect 250805 10235 250871 10236
rect 251541 10235 251607 10236
rect 252277 10235 252343 10236
rect 253105 10235 253171 10238
rect 253698 10236 253704 10300
rect 253768 10298 253774 10300
rect 253841 10298 253907 10301
rect 254485 10300 254551 10301
rect 255221 10300 255287 10301
rect 254434 10298 254440 10300
rect 253768 10296 253907 10298
rect 253768 10240 253846 10296
rect 253902 10240 253907 10296
rect 253768 10238 253907 10240
rect 254394 10238 254440 10298
rect 254504 10296 254551 10300
rect 255170 10298 255176 10300
rect 254546 10240 254551 10296
rect 253768 10236 253774 10238
rect 253841 10235 253907 10238
rect 254434 10236 254440 10238
rect 254504 10236 254551 10240
rect 255130 10238 255176 10298
rect 255240 10296 255287 10300
rect 255282 10240 255287 10296
rect 255170 10236 255176 10238
rect 255240 10236 255287 10240
rect 255906 10236 255912 10300
rect 255976 10298 255982 10300
rect 256417 10298 256483 10301
rect 256693 10300 256759 10301
rect 256642 10298 256648 10300
rect 255976 10296 256483 10298
rect 255976 10240 256422 10296
rect 256478 10240 256483 10296
rect 255976 10238 256483 10240
rect 256602 10238 256648 10298
rect 256712 10296 256759 10300
rect 256754 10240 256759 10296
rect 255976 10236 255982 10238
rect 254485 10235 254551 10236
rect 255221 10235 255287 10236
rect 256417 10235 256483 10238
rect 256642 10236 256648 10238
rect 256712 10236 256759 10240
rect 257378 10236 257384 10300
rect 257448 10298 257454 10300
rect 257705 10298 257771 10301
rect 257448 10296 257771 10298
rect 257448 10240 257710 10296
rect 257766 10240 257771 10296
rect 257448 10238 257771 10240
rect 257448 10236 257454 10238
rect 256693 10235 256759 10236
rect 257705 10235 257771 10238
rect 258114 10236 258120 10300
rect 258184 10298 258190 10300
rect 258257 10298 258323 10301
rect 258184 10296 258323 10298
rect 258184 10240 258262 10296
rect 258318 10240 258323 10296
rect 258184 10238 258323 10240
rect 258184 10236 258190 10238
rect 258257 10235 258323 10238
rect 258850 10236 258856 10300
rect 258920 10298 258926 10300
rect 258993 10298 259059 10301
rect 258920 10296 259059 10298
rect 258920 10240 258998 10296
rect 259054 10240 259059 10296
rect 258920 10238 259059 10240
rect 258920 10236 258926 10238
rect 258993 10235 259059 10238
rect 259586 10236 259592 10300
rect 259656 10298 259662 10300
rect 260005 10298 260071 10301
rect 259656 10296 260071 10298
rect 259656 10240 260010 10296
rect 260066 10240 260071 10296
rect 259656 10238 260071 10240
rect 259656 10236 259662 10238
rect 260005 10235 260071 10238
rect 260322 10236 260328 10300
rect 260392 10298 260398 10300
rect 260465 10298 260531 10301
rect 261753 10300 261819 10301
rect 262489 10300 262555 10301
rect 263225 10300 263291 10301
rect 261753 10298 261800 10300
rect 260392 10296 260531 10298
rect 260392 10240 260470 10296
rect 260526 10240 260531 10296
rect 260392 10238 260531 10240
rect 261708 10296 261800 10298
rect 261708 10240 261758 10296
rect 261708 10238 261800 10240
rect 260392 10236 260398 10238
rect 260465 10235 260531 10238
rect 261753 10236 261800 10238
rect 261864 10236 261870 10300
rect 262489 10298 262536 10300
rect 262444 10296 262536 10298
rect 262444 10240 262494 10296
rect 262444 10238 262536 10240
rect 262489 10236 262536 10238
rect 262600 10236 262606 10300
rect 263225 10298 263272 10300
rect 263180 10296 263272 10298
rect 263180 10240 263230 10296
rect 263180 10238 263272 10240
rect 263225 10236 263272 10238
rect 263336 10236 263342 10300
rect 264002 10236 264008 10300
rect 264072 10298 264078 10300
rect 264329 10298 264395 10301
rect 264072 10296 264395 10298
rect 264072 10240 264334 10296
rect 264390 10240 264395 10296
rect 264072 10238 264395 10240
rect 264072 10236 264078 10238
rect 261753 10235 261819 10236
rect 262489 10235 262555 10236
rect 263225 10235 263291 10236
rect 264329 10235 264395 10238
rect 265474 10236 265480 10300
rect 265544 10298 265550 10300
rect 265709 10298 265775 10301
rect 265544 10296 265775 10298
rect 265544 10240 265714 10296
rect 265770 10240 265775 10296
rect 265544 10238 265775 10240
rect 265544 10236 265550 10238
rect 265709 10235 265775 10238
rect 1526 10100 1532 10164
rect 1596 10162 1602 10164
rect 1669 10162 1735 10165
rect 1596 10160 1735 10162
rect 1596 10104 1674 10160
rect 1730 10104 1735 10160
rect 1596 10102 1735 10104
rect 1596 10100 1602 10102
rect 1669 10099 1735 10102
rect 2262 10100 2268 10164
rect 2332 10162 2338 10164
rect 2405 10162 2471 10165
rect 2332 10160 2471 10162
rect 2332 10104 2410 10160
rect 2466 10104 2471 10160
rect 2332 10102 2471 10104
rect 2332 10100 2338 10102
rect 2405 10099 2471 10102
rect 3233 10162 3299 10165
rect 3734 10162 3740 10164
rect 3233 10160 3740 10162
rect 3233 10104 3238 10160
rect 3294 10104 3740 10160
rect 3233 10102 3740 10104
rect 3233 10099 3299 10102
rect 3734 10100 3740 10102
rect 3804 10100 3810 10164
rect 4337 10162 4403 10165
rect 4470 10162 4476 10164
rect 4337 10160 4476 10162
rect 4337 10104 4342 10160
rect 4398 10104 4476 10160
rect 4337 10102 4476 10104
rect 4337 10099 4403 10102
rect 4470 10100 4476 10102
rect 4540 10100 4546 10164
rect 5073 10162 5139 10165
rect 5206 10162 5212 10164
rect 5073 10160 5212 10162
rect 5073 10104 5078 10160
rect 5134 10104 5212 10160
rect 5073 10102 5212 10104
rect 5073 10099 5139 10102
rect 5206 10100 5212 10102
rect 5276 10100 5282 10164
rect 5809 10162 5875 10165
rect 5942 10162 5948 10164
rect 5809 10160 5948 10162
rect 5809 10104 5814 10160
rect 5870 10104 5948 10160
rect 5809 10102 5948 10104
rect 5809 10099 5875 10102
rect 5942 10100 5948 10102
rect 6012 10100 6018 10164
rect 6678 10100 6684 10164
rect 6748 10162 6754 10164
rect 6821 10162 6887 10165
rect 6748 10160 6887 10162
rect 6748 10104 6826 10160
rect 6882 10104 6887 10160
rect 6748 10102 6887 10104
rect 6748 10100 6754 10102
rect 6821 10099 6887 10102
rect 7414 10100 7420 10164
rect 7484 10162 7490 10164
rect 7557 10162 7623 10165
rect 7484 10160 7623 10162
rect 7484 10104 7562 10160
rect 7618 10104 7623 10160
rect 7484 10102 7623 10104
rect 7484 10100 7490 10102
rect 7557 10099 7623 10102
rect 8385 10162 8451 10165
rect 8886 10162 8892 10164
rect 8385 10160 8892 10162
rect 8385 10104 8390 10160
rect 8446 10104 8892 10160
rect 8385 10102 8892 10104
rect 8385 10099 8451 10102
rect 8886 10100 8892 10102
rect 8956 10100 8962 10164
rect 11830 10100 11836 10164
rect 11900 10162 11906 10164
rect 11973 10162 12039 10165
rect 11900 10160 12039 10162
rect 11900 10104 11978 10160
rect 12034 10104 12039 10160
rect 11900 10102 12039 10104
rect 11900 10100 11906 10102
rect 11973 10099 12039 10102
rect 12566 10100 12572 10164
rect 12636 10162 12642 10164
rect 12709 10162 12775 10165
rect 12636 10160 12775 10162
rect 12636 10104 12714 10160
rect 12770 10104 12775 10160
rect 12636 10102 12775 10104
rect 12636 10100 12642 10102
rect 12709 10099 12775 10102
rect 13721 10162 13787 10165
rect 14038 10162 14044 10164
rect 13721 10160 14044 10162
rect 13721 10104 13726 10160
rect 13782 10104 14044 10160
rect 13721 10102 14044 10104
rect 13721 10099 13787 10102
rect 14038 10100 14044 10102
rect 14108 10100 14114 10164
rect 14641 10162 14707 10165
rect 14774 10162 14780 10164
rect 14641 10160 14780 10162
rect 14641 10104 14646 10160
rect 14702 10104 14780 10160
rect 14641 10102 14780 10104
rect 14641 10099 14707 10102
rect 14774 10100 14780 10102
rect 14844 10100 14850 10164
rect 15377 10162 15443 10165
rect 15510 10162 15516 10164
rect 15377 10160 15516 10162
rect 15377 10104 15382 10160
rect 15438 10104 15516 10160
rect 15377 10102 15516 10104
rect 15377 10099 15443 10102
rect 15510 10100 15516 10102
rect 15580 10100 15586 10164
rect 16113 10162 16179 10165
rect 16246 10162 16252 10164
rect 16113 10160 16252 10162
rect 16113 10104 16118 10160
rect 16174 10104 16252 10160
rect 16113 10102 16252 10104
rect 16113 10099 16179 10102
rect 16246 10100 16252 10102
rect 16316 10100 16322 10164
rect 16982 10100 16988 10164
rect 17052 10162 17058 10164
rect 17125 10162 17191 10165
rect 17052 10160 17191 10162
rect 17052 10104 17130 10160
rect 17186 10104 17191 10160
rect 17052 10102 17191 10104
rect 17052 10100 17058 10102
rect 17125 10099 17191 10102
rect 17718 10100 17724 10164
rect 17788 10162 17794 10164
rect 17861 10162 17927 10165
rect 17788 10160 17927 10162
rect 17788 10104 17866 10160
rect 17922 10104 17927 10160
rect 17788 10102 17927 10104
rect 17788 10100 17794 10102
rect 17861 10099 17927 10102
rect 18454 10100 18460 10164
rect 18524 10162 18530 10164
rect 18597 10162 18663 10165
rect 18524 10160 18663 10162
rect 18524 10104 18602 10160
rect 18658 10104 18663 10160
rect 18524 10102 18663 10104
rect 18524 10100 18530 10102
rect 18597 10099 18663 10102
rect 22134 10100 22140 10164
rect 22204 10162 22210 10164
rect 22369 10162 22435 10165
rect 138841 10164 138907 10165
rect 138790 10162 138796 10164
rect 22204 10160 22435 10162
rect 22204 10104 22374 10160
rect 22430 10104 22435 10160
rect 22204 10102 22435 10104
rect 138750 10102 138796 10162
rect 138860 10160 138907 10164
rect 138902 10104 138907 10160
rect 22204 10100 22210 10102
rect 22369 10099 22435 10102
rect 138790 10100 138796 10102
rect 138860 10100 138907 10104
rect 140262 10100 140268 10164
rect 140332 10162 140338 10164
rect 140681 10162 140747 10165
rect 140332 10160 140747 10162
rect 140332 10104 140686 10160
rect 140742 10104 140747 10160
rect 140332 10102 140747 10104
rect 140332 10100 140338 10102
rect 138841 10099 138907 10100
rect 140681 10099 140747 10102
rect 140998 10100 141004 10164
rect 141068 10162 141074 10164
rect 141325 10162 141391 10165
rect 141068 10160 141391 10162
rect 141068 10104 141330 10160
rect 141386 10104 141391 10160
rect 141068 10102 141391 10104
rect 141068 10100 141074 10102
rect 141325 10099 141391 10102
rect 141734 10100 141740 10164
rect 141804 10162 141810 10164
rect 141969 10162 142035 10165
rect 141804 10160 142035 10162
rect 141804 10104 141974 10160
rect 142030 10104 142035 10160
rect 141804 10102 142035 10104
rect 141804 10100 141810 10102
rect 141969 10099 142035 10102
rect 143206 10100 143212 10164
rect 143276 10162 143282 10164
rect 143349 10162 143415 10165
rect 143276 10160 143415 10162
rect 143276 10104 143354 10160
rect 143410 10104 143415 10160
rect 143276 10102 143415 10104
rect 143276 10100 143282 10102
rect 143349 10099 143415 10102
rect 143942 10100 143948 10164
rect 144012 10162 144018 10164
rect 144545 10162 144611 10165
rect 144012 10160 144611 10162
rect 144012 10104 144550 10160
rect 144606 10104 144611 10160
rect 144012 10102 144611 10104
rect 144012 10100 144018 10102
rect 144545 10099 144611 10102
rect 145414 10100 145420 10164
rect 145484 10162 145490 10164
rect 145833 10162 145899 10165
rect 146201 10164 146267 10165
rect 146150 10162 146156 10164
rect 145484 10160 145899 10162
rect 145484 10104 145838 10160
rect 145894 10104 145899 10160
rect 145484 10102 145899 10104
rect 146110 10102 146156 10162
rect 146220 10160 146267 10164
rect 146262 10104 146267 10160
rect 145484 10100 145490 10102
rect 145833 10099 145899 10102
rect 146150 10100 146156 10102
rect 146220 10100 146267 10104
rect 146886 10100 146892 10164
rect 146956 10162 146962 10164
rect 147121 10162 147187 10165
rect 146956 10160 147187 10162
rect 146956 10104 147126 10160
rect 147182 10104 147187 10160
rect 146956 10102 147187 10104
rect 146956 10100 146962 10102
rect 146201 10099 146267 10100
rect 147121 10099 147187 10102
rect 148358 10100 148364 10164
rect 148428 10162 148434 10164
rect 148501 10162 148567 10165
rect 148428 10160 148567 10162
rect 148428 10104 148506 10160
rect 148562 10104 148567 10160
rect 148428 10102 148567 10104
rect 148428 10100 148434 10102
rect 148501 10099 148567 10102
rect 149094 10100 149100 10164
rect 149164 10162 149170 10164
rect 149697 10162 149763 10165
rect 149164 10160 149763 10162
rect 149164 10104 149702 10160
rect 149758 10104 149763 10160
rect 149164 10102 149763 10104
rect 149164 10100 149170 10102
rect 149697 10099 149763 10102
rect 150566 10100 150572 10164
rect 150636 10162 150642 10164
rect 150985 10162 151051 10165
rect 150636 10160 151051 10162
rect 150636 10104 150990 10160
rect 151046 10104 151051 10160
rect 150636 10102 151051 10104
rect 150636 10100 150642 10102
rect 150985 10099 151051 10102
rect 151302 10100 151308 10164
rect 151372 10162 151378 10164
rect 151629 10162 151695 10165
rect 151372 10160 151695 10162
rect 151372 10104 151634 10160
rect 151690 10104 151695 10160
rect 151372 10102 151695 10104
rect 151372 10100 151378 10102
rect 151629 10099 151695 10102
rect 152038 10100 152044 10164
rect 152108 10162 152114 10164
rect 152273 10162 152339 10165
rect 152108 10160 152339 10162
rect 152108 10104 152278 10160
rect 152334 10104 152339 10160
rect 152108 10102 152339 10104
rect 152108 10100 152114 10102
rect 152273 10099 152339 10102
rect 152774 10100 152780 10164
rect 152844 10162 152850 10164
rect 153193 10162 153259 10165
rect 152844 10160 153259 10162
rect 152844 10104 153198 10160
rect 153254 10104 153259 10160
rect 152844 10102 153259 10104
rect 152844 10100 152850 10102
rect 153193 10099 153259 10102
rect 154246 10100 154252 10164
rect 154316 10162 154322 10164
rect 154573 10162 154639 10165
rect 154316 10160 154639 10162
rect 154316 10104 154578 10160
rect 154634 10104 154639 10160
rect 154316 10102 154639 10104
rect 154316 10100 154322 10102
rect 154573 10099 154639 10102
rect 206318 10100 206324 10164
rect 206388 10162 206394 10164
rect 206553 10162 206619 10165
rect 206388 10160 206619 10162
rect 206388 10104 206558 10160
rect 206614 10104 206619 10160
rect 206388 10102 206619 10104
rect 206388 10100 206394 10102
rect 206553 10099 206619 10102
rect 207054 10100 207060 10164
rect 207124 10162 207130 10164
rect 207657 10162 207723 10165
rect 207124 10160 207723 10162
rect 207124 10104 207662 10160
rect 207718 10104 207723 10160
rect 207124 10102 207723 10104
rect 207124 10100 207130 10102
rect 207657 10099 207723 10102
rect 208526 10100 208532 10164
rect 208596 10162 208602 10164
rect 208945 10162 209011 10165
rect 209313 10164 209379 10165
rect 210785 10164 210851 10165
rect 209262 10162 209268 10164
rect 208596 10160 209011 10162
rect 208596 10104 208950 10160
rect 209006 10104 209011 10160
rect 208596 10102 209011 10104
rect 209222 10102 209268 10162
rect 209332 10160 209379 10164
rect 210734 10162 210740 10164
rect 209374 10104 209379 10160
rect 208596 10100 208602 10102
rect 208945 10099 209011 10102
rect 209262 10100 209268 10102
rect 209332 10100 209379 10104
rect 210694 10102 210740 10162
rect 210804 10160 210851 10164
rect 210846 10104 210851 10160
rect 210734 10100 210740 10102
rect 210804 10100 210851 10104
rect 212942 10100 212948 10164
rect 213012 10162 213018 10164
rect 213453 10162 213519 10165
rect 213012 10160 213519 10162
rect 213012 10104 213458 10160
rect 213514 10104 213519 10160
rect 213012 10102 213519 10104
rect 213012 10100 213018 10102
rect 209313 10099 209379 10100
rect 210785 10099 210851 10100
rect 213453 10099 213519 10102
rect 213678 10100 213684 10164
rect 213748 10162 213754 10164
rect 213913 10162 213979 10165
rect 213748 10160 213979 10162
rect 213748 10104 213918 10160
rect 213974 10104 213979 10160
rect 213748 10102 213979 10104
rect 213748 10100 213754 10102
rect 213913 10099 213979 10102
rect 214414 10100 214420 10164
rect 214484 10162 214490 10164
rect 215293 10162 215359 10165
rect 214484 10160 215359 10162
rect 214484 10104 215298 10160
rect 215354 10104 215359 10160
rect 214484 10102 215359 10104
rect 214484 10100 214490 10102
rect 215293 10099 215359 10102
rect 215886 10100 215892 10164
rect 215956 10162 215962 10164
rect 216673 10162 216739 10165
rect 215956 10160 216739 10162
rect 215956 10104 216678 10160
rect 216734 10104 216739 10160
rect 215956 10102 216739 10104
rect 215956 10100 215962 10102
rect 216673 10099 216739 10102
rect 217358 10100 217364 10164
rect 217428 10162 217434 10164
rect 217961 10162 218027 10165
rect 217428 10160 218027 10162
rect 217428 10104 217966 10160
rect 218022 10104 218027 10160
rect 217428 10102 218027 10104
rect 217428 10100 217434 10102
rect 217961 10099 218027 10102
rect 218830 10100 218836 10164
rect 218900 10162 218906 10164
rect 219249 10162 219315 10165
rect 218900 10160 219315 10162
rect 218900 10104 219254 10160
rect 219310 10104 219315 10160
rect 218900 10102 219315 10104
rect 218900 10100 218906 10102
rect 219249 10099 219315 10102
rect 219566 10100 219572 10164
rect 219636 10162 219642 10164
rect 220537 10162 220603 10165
rect 223297 10164 223363 10165
rect 223246 10162 223252 10164
rect 219636 10160 220603 10162
rect 219636 10104 220542 10160
rect 220598 10104 220603 10160
rect 219636 10102 220603 10104
rect 223206 10102 223252 10162
rect 223316 10160 223363 10164
rect 223358 10104 223363 10160
rect 219636 10100 219642 10102
rect 220537 10099 220603 10102
rect 223246 10100 223252 10102
rect 223316 10100 223363 10104
rect 223297 10099 223363 10100
rect 269021 10026 269087 10029
rect 269021 10024 272442 10026
rect 269021 9968 269026 10024
rect 269082 9968 272442 10024
rect 269021 9966 272442 9968
rect 269021 9963 269087 9966
rect 2998 9828 3004 9892
rect 3068 9890 3074 9892
rect 3141 9890 3207 9893
rect 8201 9892 8267 9893
rect 8150 9890 8156 9892
rect 3068 9888 3207 9890
rect 3068 9832 3146 9888
rect 3202 9832 3207 9888
rect 3068 9830 3207 9832
rect 8110 9830 8156 9890
rect 8220 9888 8267 9892
rect 8262 9832 8267 9888
rect 3068 9828 3074 9830
rect 3141 9827 3207 9830
rect 8150 9828 8156 9830
rect 8220 9828 8267 9832
rect 10358 9828 10364 9892
rect 10428 9890 10434 9892
rect 10501 9890 10567 9893
rect 10428 9888 10567 9890
rect 10428 9832 10506 9888
rect 10562 9832 10567 9888
rect 10428 9830 10567 9832
rect 10428 9828 10434 9830
rect 8201 9827 8267 9828
rect 10501 9827 10567 9830
rect 11094 9828 11100 9892
rect 11164 9890 11170 9892
rect 11237 9890 11303 9893
rect 11164 9888 11303 9890
rect 11164 9832 11242 9888
rect 11298 9832 11303 9888
rect 11164 9830 11303 9832
rect 11164 9828 11170 9830
rect 11237 9827 11303 9830
rect 13302 9828 13308 9892
rect 13372 9890 13378 9892
rect 13445 9890 13511 9893
rect 21449 9892 21515 9893
rect 21398 9890 21404 9892
rect 13372 9888 13511 9890
rect 13372 9832 13450 9888
rect 13506 9832 13511 9888
rect 13372 9830 13511 9832
rect 21358 9830 21404 9890
rect 21468 9888 21515 9892
rect 21510 9832 21515 9888
rect 13372 9828 13378 9830
rect 13445 9827 13511 9830
rect 21398 9828 21404 9830
rect 21468 9828 21515 9832
rect 85246 9828 85252 9892
rect 85316 9890 85322 9892
rect 85389 9890 85455 9893
rect 85316 9888 85455 9890
rect 85316 9832 85394 9888
rect 85450 9832 85455 9888
rect 85316 9830 85455 9832
rect 85316 9828 85322 9830
rect 21449 9827 21515 9828
rect 85389 9827 85455 9830
rect 85982 9828 85988 9892
rect 86052 9890 86058 9892
rect 86493 9890 86559 9893
rect 86052 9888 86559 9890
rect 86052 9832 86498 9888
rect 86554 9832 86559 9888
rect 86052 9830 86559 9832
rect 86052 9828 86058 9830
rect 86493 9827 86559 9830
rect 139526 9828 139532 9892
rect 139596 9890 139602 9892
rect 139761 9890 139827 9893
rect 144729 9892 144795 9893
rect 144678 9890 144684 9892
rect 139596 9888 139827 9890
rect 139596 9832 139766 9888
rect 139822 9832 139827 9888
rect 139596 9830 139827 9832
rect 144638 9830 144684 9890
rect 144748 9888 144795 9892
rect 144790 9832 144795 9888
rect 139596 9828 139602 9830
rect 139761 9827 139827 9830
rect 144678 9828 144684 9830
rect 144748 9828 144795 9832
rect 149830 9828 149836 9892
rect 149900 9890 149906 9892
rect 150065 9890 150131 9893
rect 149900 9888 150131 9890
rect 149900 9832 150070 9888
rect 150126 9832 150131 9888
rect 149900 9830 150131 9832
rect 149900 9828 149906 9830
rect 144729 9827 144795 9828
rect 150065 9827 150131 9830
rect 154982 9828 154988 9892
rect 155052 9890 155058 9892
rect 155125 9890 155191 9893
rect 155052 9888 155191 9890
rect 155052 9832 155130 9888
rect 155186 9832 155191 9888
rect 155052 9830 155191 9832
rect 155052 9828 155058 9830
rect 155125 9827 155191 9830
rect 216622 9828 216628 9892
rect 216692 9890 216698 9892
rect 216857 9890 216923 9893
rect 216692 9888 216923 9890
rect 216692 9832 216862 9888
rect 216918 9832 216923 9888
rect 216692 9830 216923 9832
rect 216692 9828 216698 9830
rect 216857 9827 216923 9830
rect 68542 9824 68858 9825
rect 68542 9760 68548 9824
rect 68612 9760 68628 9824
rect 68692 9760 68708 9824
rect 68772 9760 68788 9824
rect 68852 9760 68858 9824
rect 68542 9759 68858 9760
rect 136139 9824 136455 9825
rect 136139 9760 136145 9824
rect 136209 9760 136225 9824
rect 136289 9760 136305 9824
rect 136369 9760 136385 9824
rect 136449 9760 136455 9824
rect 136139 9759 136455 9760
rect 203736 9824 204052 9825
rect 203736 9760 203742 9824
rect 203806 9760 203822 9824
rect 203886 9760 203902 9824
rect 203966 9760 203982 9824
rect 204046 9760 204052 9824
rect 203736 9759 204052 9760
rect 271333 9824 271649 9825
rect 271333 9760 271339 9824
rect 271403 9760 271419 9824
rect 271483 9760 271499 9824
rect 271563 9760 271579 9824
rect 271643 9760 271649 9824
rect 271333 9759 271649 9760
rect 76465 9756 76531 9757
rect 79409 9756 79475 9757
rect 81617 9756 81683 9757
rect 76414 9754 76420 9756
rect 76374 9694 76420 9754
rect 76484 9752 76531 9756
rect 79358 9754 79364 9756
rect 76526 9696 76531 9752
rect 76414 9692 76420 9694
rect 76484 9692 76531 9696
rect 79318 9694 79364 9754
rect 79428 9752 79475 9756
rect 81566 9754 81572 9756
rect 79470 9696 79475 9752
rect 79358 9692 79364 9694
rect 79428 9692 79475 9696
rect 81526 9694 81572 9754
rect 81636 9752 81683 9756
rect 81678 9696 81683 9752
rect 81566 9692 81572 9694
rect 81636 9692 81683 9696
rect 93342 9692 93348 9756
rect 93412 9754 93418 9756
rect 93485 9754 93551 9757
rect 93412 9752 93551 9754
rect 93412 9696 93490 9752
rect 93546 9696 93551 9752
rect 93412 9694 93551 9696
rect 93412 9692 93418 9694
rect 76465 9691 76531 9692
rect 79409 9691 79475 9692
rect 81617 9691 81683 9692
rect 93485 9691 93551 9694
rect 95550 9692 95556 9756
rect 95620 9754 95626 9756
rect 95969 9754 96035 9757
rect 96337 9756 96403 9757
rect 95620 9752 96035 9754
rect 95620 9696 95974 9752
rect 96030 9696 96035 9752
rect 95620 9694 96035 9696
rect 95620 9692 95626 9694
rect 95969 9691 96035 9694
rect 96286 9692 96292 9756
rect 96356 9754 96403 9756
rect 96356 9752 96448 9754
rect 96398 9696 96448 9752
rect 96356 9694 96448 9696
rect 96356 9692 96403 9694
rect 97758 9692 97764 9756
rect 97828 9754 97834 9756
rect 97993 9754 98059 9757
rect 100661 9756 100727 9757
rect 100661 9754 100708 9756
rect 97828 9752 98059 9754
rect 97828 9696 97998 9752
rect 98054 9696 98059 9752
rect 97828 9694 98059 9696
rect 100616 9752 100708 9754
rect 100616 9696 100666 9752
rect 100616 9694 100708 9696
rect 97828 9692 97834 9694
rect 96337 9691 96403 9692
rect 97993 9691 98059 9694
rect 100661 9692 100708 9694
rect 100772 9692 100778 9756
rect 155718 9692 155724 9756
rect 155788 9754 155794 9756
rect 155953 9754 156019 9757
rect 155788 9752 156019 9754
rect 155788 9696 155958 9752
rect 156014 9696 156019 9752
rect 155788 9694 156019 9696
rect 155788 9692 155794 9694
rect 100661 9691 100727 9692
rect 155953 9691 156019 9694
rect 156454 9692 156460 9756
rect 156524 9754 156530 9756
rect 156873 9754 156939 9757
rect 157977 9756 158043 9757
rect 159449 9756 159515 9757
rect 163865 9756 163931 9757
rect 156524 9752 156939 9754
rect 156524 9696 156878 9752
rect 156934 9696 156939 9752
rect 156524 9694 156939 9696
rect 156524 9692 156530 9694
rect 156873 9691 156939 9694
rect 157926 9692 157932 9756
rect 157996 9754 158043 9756
rect 157996 9752 158088 9754
rect 158038 9696 158088 9752
rect 157996 9694 158088 9696
rect 157996 9692 158043 9694
rect 159398 9692 159404 9756
rect 159468 9754 159515 9756
rect 159468 9752 159560 9754
rect 159510 9696 159560 9752
rect 159468 9694 159560 9696
rect 159468 9692 159515 9694
rect 163814 9692 163820 9756
rect 163884 9754 163931 9756
rect 163884 9752 163976 9754
rect 163926 9696 163976 9752
rect 163884 9694 163976 9696
rect 163884 9692 163931 9694
rect 225454 9692 225460 9756
rect 225524 9754 225530 9756
rect 225689 9754 225755 9757
rect 229829 9756 229895 9757
rect 229829 9754 229876 9756
rect 225524 9752 225755 9754
rect 225524 9696 225694 9752
rect 225750 9696 225755 9752
rect 225524 9694 225755 9696
rect 229784 9752 229876 9754
rect 229784 9696 229834 9752
rect 229784 9694 229876 9696
rect 225524 9692 225530 9694
rect 157977 9691 158043 9692
rect 159449 9691 159515 9692
rect 163865 9691 163931 9692
rect 225689 9691 225755 9694
rect 229829 9692 229876 9694
rect 229940 9692 229946 9756
rect 231342 9692 231348 9756
rect 231412 9754 231418 9756
rect 231577 9754 231643 9757
rect 233509 9756 233575 9757
rect 234337 9756 234403 9757
rect 235073 9756 235139 9757
rect 233509 9754 233556 9756
rect 231412 9752 231643 9754
rect 231412 9696 231582 9752
rect 231638 9696 231643 9752
rect 231412 9694 231643 9696
rect 233464 9752 233556 9754
rect 233464 9696 233514 9752
rect 233464 9694 233556 9696
rect 231412 9692 231418 9694
rect 229829 9691 229895 9692
rect 231577 9691 231643 9694
rect 233509 9692 233556 9694
rect 233620 9692 233626 9756
rect 234286 9692 234292 9756
rect 234356 9754 234403 9756
rect 234356 9752 234448 9754
rect 234398 9696 234448 9752
rect 234356 9694 234448 9696
rect 234356 9692 234403 9694
rect 235022 9692 235028 9756
rect 235092 9754 235139 9756
rect 272382 9754 272442 9966
rect 235092 9752 235184 9754
rect 235134 9696 235184 9752
rect 235092 9694 235184 9696
rect 272198 9694 272442 9754
rect 235092 9692 235139 9694
rect 233509 9691 233575 9692
rect 234337 9691 234403 9692
rect 235073 9691 235139 9692
rect 25865 9620 25931 9621
rect 25814 9556 25820 9620
rect 25884 9618 25931 9620
rect 25884 9616 25976 9618
rect 25926 9560 25976 9616
rect 25884 9558 25976 9560
rect 25884 9556 25931 9558
rect 32438 9556 32444 9620
rect 32508 9618 32514 9620
rect 32581 9618 32647 9621
rect 69105 9620 69171 9621
rect 32508 9616 32647 9618
rect 32508 9560 32586 9616
rect 32642 9560 32647 9616
rect 32508 9558 32647 9560
rect 32508 9556 32514 9558
rect 25865 9555 25931 9556
rect 32581 9555 32647 9558
rect 69054 9556 69060 9620
rect 69124 9618 69171 9620
rect 70301 9618 70367 9621
rect 70526 9618 70532 9620
rect 69124 9616 69216 9618
rect 69166 9560 69216 9616
rect 69124 9558 69216 9560
rect 70301 9616 70532 9618
rect 70301 9560 70306 9616
rect 70362 9560 70532 9616
rect 70301 9558 70532 9560
rect 69124 9556 69171 9558
rect 69105 9555 69171 9556
rect 70301 9555 70367 9558
rect 70526 9556 70532 9558
rect 70596 9556 70602 9620
rect 72141 9618 72207 9621
rect 72734 9618 72740 9620
rect 72141 9616 72740 9618
rect 72141 9560 72146 9616
rect 72202 9560 72740 9616
rect 72141 9558 72740 9560
rect 72141 9555 72207 9558
rect 72734 9556 72740 9558
rect 72804 9556 72810 9620
rect 74717 9618 74783 9621
rect 75678 9618 75684 9620
rect 74717 9616 75684 9618
rect 74717 9560 74722 9616
rect 74778 9560 75684 9616
rect 74717 9558 75684 9560
rect 74717 9555 74783 9558
rect 75678 9556 75684 9558
rect 75748 9556 75754 9620
rect 77293 9618 77359 9621
rect 77886 9618 77892 9620
rect 77293 9616 77892 9618
rect 77293 9560 77298 9616
rect 77354 9560 77892 9616
rect 77293 9558 77892 9560
rect 77293 9555 77359 9558
rect 77886 9556 77892 9558
rect 77956 9556 77962 9620
rect 79961 9618 80027 9621
rect 80830 9618 80836 9620
rect 79961 9616 80836 9618
rect 79961 9560 79966 9616
rect 80022 9560 80836 9616
rect 79961 9558 80836 9560
rect 79961 9555 80027 9558
rect 80830 9556 80836 9558
rect 80900 9556 80906 9620
rect 82629 9618 82695 9621
rect 137369 9620 137435 9621
rect 83038 9618 83044 9620
rect 82629 9616 83044 9618
rect 82629 9560 82634 9616
rect 82690 9560 83044 9616
rect 82629 9558 83044 9560
rect 82629 9555 82695 9558
rect 83038 9556 83044 9558
rect 83108 9556 83114 9620
rect 137318 9556 137324 9620
rect 137388 9618 137435 9620
rect 137388 9616 137480 9618
rect 137430 9560 137480 9616
rect 137388 9558 137480 9560
rect 137388 9556 137435 9558
rect 205582 9556 205588 9620
rect 205652 9618 205658 9620
rect 205817 9618 205883 9621
rect 205652 9616 205883 9618
rect 205652 9560 205822 9616
rect 205878 9560 205883 9616
rect 205652 9558 205883 9560
rect 205652 9556 205658 9558
rect 137369 9555 137435 9556
rect 205817 9555 205883 9558
rect 268469 9618 268535 9621
rect 272198 9618 272258 9694
rect 268469 9616 272074 9618
rect 268469 9560 268474 9616
rect 268530 9560 272074 9616
rect 268469 9558 272074 9560
rect 272198 9558 272504 9618
rect 268469 9555 268535 9558
rect 28809 9484 28875 9485
rect 28758 9420 28764 9484
rect 28828 9482 28875 9484
rect 28828 9480 28920 9482
rect 28870 9424 28920 9480
rect 28828 9422 28920 9424
rect 28828 9420 28875 9422
rect 158662 9420 158668 9484
rect 158732 9482 158738 9484
rect 159449 9482 159515 9485
rect 158732 9480 159515 9482
rect 158732 9424 159454 9480
rect 159510 9424 159515 9480
rect 158732 9422 159515 9424
rect 158732 9420 158738 9422
rect 28809 9419 28875 9420
rect 159449 9419 159515 9422
rect 224769 9482 224835 9485
rect 225965 9482 226031 9485
rect 224769 9480 226031 9482
rect 224769 9424 224774 9480
rect 224830 9424 225970 9480
rect 226026 9424 226031 9480
rect 224769 9422 226031 9424
rect 224769 9419 224835 9422
rect 225965 9419 226031 9422
rect 228265 9482 228331 9485
rect 228398 9482 228404 9484
rect 228265 9480 228404 9482
rect 228265 9424 228270 9480
rect 228326 9424 228404 9480
rect 228265 9422 228404 9424
rect 228265 9419 228331 9422
rect 228398 9420 228404 9422
rect 228468 9420 228474 9484
rect 267641 9482 267707 9485
rect 271781 9482 271847 9485
rect 267641 9480 271847 9482
rect 267641 9424 267646 9480
rect 267702 9424 271786 9480
rect 271842 9424 271847 9480
rect 267641 9422 271847 9424
rect 272014 9482 272074 9558
rect 272014 9422 272504 9482
rect 267641 9419 267707 9422
rect 271781 9419 271847 9422
rect 268929 9346 268995 9349
rect 268929 9344 272504 9346
rect 268929 9288 268934 9344
rect 268990 9288 272504 9344
rect 268929 9286 272504 9288
rect 268929 9283 268995 9286
rect 34744 9280 35060 9281
rect 34744 9216 34750 9280
rect 34814 9216 34830 9280
rect 34894 9216 34910 9280
rect 34974 9216 34990 9280
rect 35054 9216 35060 9280
rect 34744 9215 35060 9216
rect 102341 9280 102657 9281
rect 102341 9216 102347 9280
rect 102411 9216 102427 9280
rect 102491 9216 102507 9280
rect 102571 9216 102587 9280
rect 102651 9216 102657 9280
rect 102341 9215 102657 9216
rect 169938 9280 170254 9281
rect 169938 9216 169944 9280
rect 170008 9216 170024 9280
rect 170088 9216 170104 9280
rect 170168 9216 170184 9280
rect 170248 9216 170254 9280
rect 169938 9215 170254 9216
rect 237535 9280 237851 9281
rect 237535 9216 237541 9280
rect 237605 9216 237621 9280
rect 237685 9216 237701 9280
rect 237765 9216 237781 9280
rect 237845 9216 237851 9280
rect 237535 9215 237851 9216
rect 790 9148 796 9212
rect 860 9210 866 9212
rect 1393 9210 1459 9213
rect 860 9208 1459 9210
rect 860 9152 1398 9208
rect 1454 9152 1459 9208
rect 860 9150 1459 9152
rect 860 9148 866 9150
rect 1393 9147 1459 9150
rect 88190 9148 88196 9212
rect 88260 9210 88266 9212
rect 88333 9210 88399 9213
rect 169017 9212 169083 9213
rect 88260 9208 88399 9210
rect 88260 9152 88338 9208
rect 88394 9152 88399 9208
rect 88260 9150 88399 9152
rect 88260 9148 88266 9150
rect 88333 9147 88399 9150
rect 168966 9148 168972 9212
rect 169036 9210 169083 9212
rect 223481 9210 223547 9213
rect 223982 9210 223988 9212
rect 169036 9208 169128 9210
rect 169078 9152 169128 9208
rect 169036 9150 169128 9152
rect 223481 9208 223988 9210
rect 223481 9152 223486 9208
rect 223542 9152 223988 9208
rect 223481 9150 223988 9152
rect 169036 9148 169083 9150
rect 169017 9147 169083 9148
rect 223481 9147 223547 9150
rect 223982 9148 223988 9150
rect 224052 9148 224058 9212
rect 235758 9148 235764 9212
rect 235828 9210 235834 9212
rect 235993 9210 236059 9213
rect 237281 9212 237347 9213
rect 235828 9208 236059 9210
rect 235828 9152 235998 9208
rect 236054 9152 236059 9208
rect 235828 9150 236059 9152
rect 235828 9148 235834 9150
rect 235993 9147 236059 9150
rect 237230 9148 237236 9212
rect 237300 9210 237347 9212
rect 268009 9210 268075 9213
rect 237300 9208 237392 9210
rect 237342 9152 237392 9208
rect 237300 9150 237392 9152
rect 268009 9208 272504 9210
rect 268009 9152 268014 9208
rect 268070 9152 272504 9208
rect 268009 9150 272504 9152
rect 237300 9148 237347 9150
rect 237281 9147 237347 9148
rect 268009 9147 268075 9150
rect 69565 9074 69631 9077
rect 73429 9076 73495 9077
rect 69790 9074 69796 9076
rect 69565 9072 69796 9074
rect 69565 9016 69570 9072
rect 69626 9016 69796 9072
rect 69565 9014 69796 9016
rect 69565 9011 69631 9014
rect 69790 9012 69796 9014
rect 69860 9012 69866 9076
rect 73429 9074 73476 9076
rect 73384 9072 73476 9074
rect 73384 9016 73434 9072
rect 73384 9014 73476 9016
rect 73429 9012 73476 9014
rect 73540 9012 73546 9076
rect 74717 9074 74783 9077
rect 78581 9076 78647 9077
rect 74942 9074 74948 9076
rect 74717 9072 74948 9074
rect 74717 9016 74722 9072
rect 74778 9016 74948 9072
rect 74717 9014 74948 9016
rect 73429 9011 73495 9012
rect 74717 9011 74783 9014
rect 74942 9012 74948 9014
rect 75012 9012 75018 9076
rect 78581 9074 78628 9076
rect 78536 9072 78628 9074
rect 78536 9016 78586 9072
rect 78536 9014 78628 9016
rect 78581 9012 78628 9014
rect 78692 9012 78698 9076
rect 79961 9074 80027 9077
rect 80094 9074 80100 9076
rect 79961 9072 80100 9074
rect 79961 9016 79966 9072
rect 80022 9016 80100 9072
rect 79961 9014 80100 9016
rect 78581 9011 78647 9012
rect 79961 9011 80027 9014
rect 80094 9012 80100 9014
rect 80164 9012 80170 9076
rect 193305 9074 193371 9077
rect 198181 9074 198247 9077
rect 193305 9072 198247 9074
rect 193305 9016 193310 9072
rect 193366 9016 198186 9072
rect 198242 9016 198247 9072
rect 193305 9014 198247 9016
rect 193305 9011 193371 9014
rect 198181 9011 198247 9014
rect 268101 9074 268167 9077
rect 268101 9072 272504 9074
rect 268101 9016 268106 9072
rect 268162 9016 272504 9072
rect 268101 9014 272504 9016
rect 268101 9011 268167 9014
rect 225597 8938 225663 8941
rect 227161 8938 227227 8941
rect 228449 8938 228515 8941
rect 225597 8936 228515 8938
rect 225597 8880 225602 8936
rect 225658 8880 227166 8936
rect 227222 8880 228454 8936
rect 228510 8880 228515 8936
rect 225597 8878 228515 8880
rect 225597 8875 225663 8878
rect 227161 8875 227227 8878
rect 228449 8875 228515 8878
rect 267917 8938 267983 8941
rect 271965 8938 272031 8941
rect 267917 8936 271890 8938
rect 267917 8880 267922 8936
rect 267978 8880 271890 8936
rect 267917 8878 271890 8880
rect 267917 8875 267983 8878
rect 24025 8802 24091 8805
rect 25681 8802 25747 8805
rect 24025 8800 25747 8802
rect 24025 8744 24030 8800
rect 24086 8744 25686 8800
rect 25742 8744 25747 8800
rect 24025 8742 25747 8744
rect 24025 8739 24091 8742
rect 25681 8739 25747 8742
rect 91134 8740 91140 8804
rect 91204 8802 91210 8804
rect 91829 8802 91895 8805
rect 91204 8800 91895 8802
rect 91204 8744 91834 8800
rect 91890 8744 91895 8800
rect 91204 8742 91895 8744
rect 91204 8740 91210 8742
rect 91829 8739 91895 8742
rect 223941 8802 224007 8805
rect 228817 8802 228883 8805
rect 230105 8802 230171 8805
rect 223941 8800 230171 8802
rect 223941 8744 223946 8800
rect 224002 8744 228822 8800
rect 228878 8744 230110 8800
rect 230166 8744 230171 8800
rect 223941 8742 230171 8744
rect 223941 8739 224007 8742
rect 228817 8739 228883 8742
rect 230105 8739 230171 8742
rect 262070 8740 262076 8804
rect 262140 8802 262146 8804
rect 262581 8802 262647 8805
rect 262140 8800 262647 8802
rect 262140 8744 262586 8800
rect 262642 8744 262647 8800
rect 262140 8742 262647 8744
rect 271830 8802 271890 8878
rect 271965 8936 272504 8938
rect 271965 8880 271970 8936
rect 272026 8880 272504 8936
rect 271965 8878 272504 8880
rect 271965 8875 272031 8878
rect 271830 8742 272504 8802
rect 262140 8740 262146 8742
rect 262581 8739 262647 8742
rect 68542 8736 68858 8737
rect 68542 8672 68548 8736
rect 68612 8672 68628 8736
rect 68692 8672 68708 8736
rect 68772 8672 68788 8736
rect 68852 8672 68858 8736
rect 68542 8671 68858 8672
rect 136139 8736 136455 8737
rect 136139 8672 136145 8736
rect 136209 8672 136225 8736
rect 136289 8672 136305 8736
rect 136369 8672 136385 8736
rect 136449 8672 136455 8736
rect 136139 8671 136455 8672
rect 203736 8736 204052 8737
rect 203736 8672 203742 8736
rect 203806 8672 203822 8736
rect 203886 8672 203902 8736
rect 203966 8672 203982 8736
rect 204046 8672 204052 8736
rect 203736 8671 204052 8672
rect 271333 8736 271649 8737
rect 271333 8672 271339 8736
rect 271403 8672 271419 8736
rect 271483 8672 271499 8736
rect 271563 8672 271579 8736
rect 271643 8672 271649 8736
rect 271333 8671 271649 8672
rect 23473 8666 23539 8669
rect 24342 8666 24348 8668
rect 23473 8664 24348 8666
rect 23473 8608 23478 8664
rect 23534 8608 24348 8664
rect 23473 8606 24348 8608
rect 23473 8603 23539 8606
rect 24342 8604 24348 8606
rect 24412 8604 24418 8668
rect 29494 8604 29500 8668
rect 29564 8666 29570 8668
rect 29637 8666 29703 8669
rect 30189 8668 30255 8669
rect 30189 8666 30236 8668
rect 29564 8664 29703 8666
rect 29564 8608 29642 8664
rect 29698 8608 29703 8664
rect 29564 8606 29703 8608
rect 30144 8664 30236 8666
rect 30144 8608 30194 8664
rect 30144 8606 30236 8608
rect 29564 8604 29570 8606
rect 29637 8603 29703 8606
rect 30189 8604 30236 8606
rect 30300 8604 30306 8668
rect 30966 8604 30972 8668
rect 31036 8666 31042 8668
rect 31293 8666 31359 8669
rect 31036 8664 31359 8666
rect 31036 8608 31298 8664
rect 31354 8608 31359 8664
rect 31036 8606 31359 8608
rect 31036 8604 31042 8606
rect 30189 8603 30255 8604
rect 31293 8603 31359 8606
rect 87454 8604 87460 8668
rect 87524 8666 87530 8668
rect 88333 8666 88399 8669
rect 90449 8668 90515 8669
rect 91921 8668 91987 8669
rect 87524 8664 88399 8666
rect 87524 8608 88338 8664
rect 88394 8608 88399 8664
rect 87524 8606 88399 8608
rect 87524 8604 87530 8606
rect 88333 8603 88399 8606
rect 90398 8604 90404 8668
rect 90468 8666 90515 8668
rect 90468 8664 90560 8666
rect 90510 8608 90560 8664
rect 90468 8606 90560 8608
rect 90468 8604 90515 8606
rect 91870 8604 91876 8668
rect 91940 8666 91987 8668
rect 91940 8664 92032 8666
rect 91982 8608 92032 8664
rect 91940 8606 92032 8608
rect 91940 8604 91987 8606
rect 94078 8604 94084 8668
rect 94148 8666 94154 8668
rect 94589 8666 94655 8669
rect 94865 8668 94931 8669
rect 94148 8664 94655 8666
rect 94148 8608 94594 8664
rect 94650 8608 94655 8664
rect 94148 8606 94655 8608
rect 94148 8604 94154 8606
rect 90449 8603 90515 8604
rect 91921 8603 91987 8604
rect 94589 8603 94655 8606
rect 94814 8604 94820 8668
rect 94884 8666 94931 8668
rect 94884 8664 94976 8666
rect 94926 8608 94976 8664
rect 94884 8606 94976 8608
rect 94884 8604 94931 8606
rect 97022 8604 97028 8668
rect 97092 8666 97098 8668
rect 97441 8666 97507 8669
rect 97092 8664 97507 8666
rect 97092 8608 97446 8664
rect 97502 8608 97507 8664
rect 97092 8606 97507 8608
rect 97092 8604 97098 8606
rect 94865 8603 94931 8604
rect 97441 8603 97507 8606
rect 98494 8604 98500 8668
rect 98564 8666 98570 8668
rect 98637 8666 98703 8669
rect 98564 8664 98703 8666
rect 98564 8608 98642 8664
rect 98698 8608 98703 8664
rect 98564 8606 98703 8608
rect 98564 8604 98570 8606
rect 98637 8603 98703 8606
rect 99966 8604 99972 8668
rect 100036 8666 100042 8668
rect 100293 8666 100359 8669
rect 100036 8664 100359 8666
rect 100036 8608 100298 8664
rect 100354 8608 100359 8664
rect 100036 8606 100359 8608
rect 100036 8604 100042 8606
rect 100293 8603 100359 8606
rect 225965 8666 226031 8669
rect 226190 8666 226196 8668
rect 225965 8664 226196 8666
rect 225965 8608 225970 8664
rect 226026 8608 226196 8664
rect 225965 8606 226196 8608
rect 225965 8603 226031 8606
rect 226190 8604 226196 8606
rect 226260 8604 226266 8668
rect 226701 8666 226767 8669
rect 226926 8666 226932 8668
rect 226701 8664 226932 8666
rect 226701 8608 226706 8664
rect 226762 8608 226932 8664
rect 226701 8606 226932 8608
rect 226701 8603 226767 8606
rect 226926 8604 226932 8606
rect 226996 8604 227002 8668
rect 227662 8604 227668 8668
rect 227732 8666 227738 8668
rect 228265 8666 228331 8669
rect 229093 8668 229159 8669
rect 229093 8666 229140 8668
rect 227732 8664 228331 8666
rect 227732 8608 228270 8664
rect 228326 8608 228331 8664
rect 227732 8606 228331 8608
rect 229048 8664 229140 8666
rect 229048 8608 229098 8664
rect 229048 8606 229140 8608
rect 227732 8604 227738 8606
rect 228265 8603 228331 8606
rect 229093 8604 229140 8606
rect 229204 8604 229210 8668
rect 231945 8666 232011 8669
rect 232865 8668 232931 8669
rect 232078 8666 232084 8668
rect 231945 8664 232084 8666
rect 231945 8608 231950 8664
rect 232006 8608 232084 8664
rect 231945 8606 232084 8608
rect 229093 8603 229159 8604
rect 231945 8603 232011 8606
rect 232078 8604 232084 8606
rect 232148 8604 232154 8668
rect 232814 8604 232820 8668
rect 232884 8666 232931 8668
rect 232884 8664 232976 8666
rect 232926 8608 232976 8664
rect 232884 8606 232976 8608
rect 232884 8604 232931 8606
rect 236494 8604 236500 8668
rect 236564 8666 236570 8668
rect 236637 8666 236703 8669
rect 236564 8664 236703 8666
rect 236564 8608 236642 8664
rect 236698 8608 236703 8664
rect 236564 8606 236703 8608
rect 272304 8606 272504 8666
rect 236564 8604 236570 8606
rect 232865 8603 232931 8604
rect 236637 8603 236703 8606
rect 161606 8468 161612 8532
rect 161676 8530 161682 8532
rect 162301 8530 162367 8533
rect 268837 8530 268903 8533
rect 161676 8528 162367 8530
rect 161676 8472 162306 8528
rect 162362 8472 162367 8528
rect 161676 8470 162367 8472
rect 161676 8468 161682 8470
rect 162301 8467 162367 8470
rect 263550 8528 268903 8530
rect 263550 8472 268842 8528
rect 268898 8472 268903 8528
rect 263550 8470 268903 8472
rect 26550 8332 26556 8396
rect 26620 8394 26626 8396
rect 26693 8394 26759 8397
rect 26620 8392 26759 8394
rect 26620 8336 26698 8392
rect 26754 8336 26759 8392
rect 26620 8334 26759 8336
rect 26620 8332 26626 8334
rect 26693 8331 26759 8334
rect 28022 8332 28028 8396
rect 28092 8394 28098 8396
rect 28349 8394 28415 8397
rect 28092 8392 28415 8394
rect 28092 8336 28354 8392
rect 28410 8336 28415 8392
rect 28092 8334 28415 8336
rect 28092 8332 28098 8334
rect 28349 8331 28415 8334
rect 92606 8332 92612 8396
rect 92676 8394 92682 8396
rect 93301 8394 93367 8397
rect 92676 8392 93367 8394
rect 92676 8336 93306 8392
rect 93362 8336 93367 8392
rect 92676 8334 93367 8336
rect 92676 8332 92682 8334
rect 93301 8331 93367 8334
rect 160134 8332 160140 8396
rect 160204 8394 160210 8396
rect 160277 8394 160343 8397
rect 160204 8392 160343 8394
rect 160204 8336 160282 8392
rect 160338 8336 160343 8392
rect 160204 8334 160343 8336
rect 160204 8332 160210 8334
rect 160277 8331 160343 8334
rect 160870 8332 160876 8396
rect 160940 8394 160946 8396
rect 161289 8394 161355 8397
rect 160940 8392 161355 8394
rect 160940 8336 161294 8392
rect 161350 8336 161355 8392
rect 160940 8334 161355 8336
rect 160940 8332 160946 8334
rect 161289 8331 161355 8334
rect 162342 8332 162348 8396
rect 162412 8394 162418 8396
rect 162577 8394 162643 8397
rect 162412 8392 162643 8394
rect 162412 8336 162582 8392
rect 162638 8336 162643 8392
rect 162412 8334 162643 8336
rect 162412 8332 162418 8334
rect 162577 8331 162643 8334
rect 163078 8332 163084 8396
rect 163148 8394 163154 8396
rect 164049 8394 164115 8397
rect 163148 8392 164115 8394
rect 163148 8336 164054 8392
rect 164110 8336 164115 8392
rect 163148 8334 164115 8336
rect 163148 8332 163154 8334
rect 164049 8331 164115 8334
rect 164550 8332 164556 8396
rect 164620 8394 164626 8396
rect 164785 8394 164851 8397
rect 164620 8392 164851 8394
rect 164620 8336 164790 8392
rect 164846 8336 164851 8392
rect 164620 8334 164851 8336
rect 164620 8332 164626 8334
rect 164785 8331 164851 8334
rect 165286 8332 165292 8396
rect 165356 8394 165362 8396
rect 165521 8394 165587 8397
rect 165356 8392 165587 8394
rect 165356 8336 165526 8392
rect 165582 8336 165587 8392
rect 165356 8334 165587 8336
rect 165356 8332 165362 8334
rect 165521 8331 165587 8334
rect 166022 8332 166028 8396
rect 166092 8394 166098 8396
rect 166349 8394 166415 8397
rect 166092 8392 166415 8394
rect 166092 8336 166354 8392
rect 166410 8336 166415 8392
rect 166092 8334 166415 8336
rect 166092 8332 166098 8334
rect 166349 8331 166415 8334
rect 167494 8332 167500 8396
rect 167564 8394 167570 8396
rect 167821 8394 167887 8397
rect 224769 8396 224835 8397
rect 224718 8394 224724 8396
rect 167564 8392 167887 8394
rect 167564 8336 167826 8392
rect 167882 8336 167887 8392
rect 167564 8334 167887 8336
rect 224678 8334 224724 8394
rect 224788 8392 224835 8396
rect 224830 8336 224835 8392
rect 167564 8332 167570 8334
rect 167821 8331 167887 8334
rect 224718 8332 224724 8334
rect 224788 8332 224835 8336
rect 230606 8332 230612 8396
rect 230676 8394 230682 8396
rect 230841 8394 230907 8397
rect 230676 8392 230907 8394
rect 230676 8336 230846 8392
rect 230902 8336 230907 8392
rect 230676 8334 230907 8336
rect 230676 8332 230682 8334
rect 224769 8331 224835 8332
rect 230841 8331 230907 8334
rect 235257 8394 235323 8397
rect 258165 8394 258231 8397
rect 235257 8392 258231 8394
rect 235257 8336 235262 8392
rect 235318 8336 258170 8392
rect 258226 8336 258231 8392
rect 235257 8334 258231 8336
rect 235257 8331 235323 8334
rect 258165 8331 258231 8334
rect 262857 8394 262923 8397
rect 263174 8394 263180 8396
rect 262857 8392 263180 8394
rect 262857 8336 262862 8392
rect 262918 8336 263180 8392
rect 262857 8334 263180 8336
rect 262857 8331 262923 8334
rect 263174 8332 263180 8334
rect 263244 8332 263250 8396
rect 99281 8260 99347 8261
rect 166809 8260 166875 8261
rect 99230 8258 99236 8260
rect 99190 8198 99236 8258
rect 99300 8256 99347 8260
rect 166758 8258 166764 8260
rect 99342 8200 99347 8256
rect 99230 8196 99236 8198
rect 99300 8196 99347 8200
rect 166718 8198 166764 8258
rect 166828 8256 166875 8260
rect 166870 8200 166875 8256
rect 166758 8196 166764 8198
rect 166828 8196 166875 8200
rect 99281 8195 99347 8196
rect 166809 8195 166875 8196
rect 226333 8258 226399 8261
rect 237097 8258 237163 8261
rect 226333 8256 237163 8258
rect 226333 8200 226338 8256
rect 226394 8200 237102 8256
rect 237158 8200 237163 8256
rect 226333 8198 237163 8200
rect 226333 8195 226399 8198
rect 237097 8195 237163 8198
rect 262305 8258 262371 8261
rect 263550 8258 263610 8470
rect 268837 8467 268903 8470
rect 270585 8530 270651 8533
rect 270585 8528 272504 8530
rect 270585 8472 270590 8528
rect 270646 8472 272504 8528
rect 270585 8470 272504 8472
rect 270585 8467 270651 8470
rect 266445 8396 266511 8397
rect 266445 8394 266492 8396
rect 266400 8392 266492 8394
rect 266400 8336 266450 8392
rect 266400 8334 266492 8336
rect 266445 8332 266492 8334
rect 266556 8332 266562 8396
rect 271229 8394 271295 8397
rect 271229 8392 272504 8394
rect 271229 8336 271234 8392
rect 271290 8336 272504 8392
rect 271229 8334 272504 8336
rect 266445 8331 266511 8332
rect 271229 8331 271295 8334
rect 262305 8256 263610 8258
rect 262305 8200 262310 8256
rect 262366 8200 263610 8256
rect 262305 8198 263610 8200
rect 270493 8258 270559 8261
rect 270493 8256 272504 8258
rect 270493 8200 270498 8256
rect 270554 8200 272504 8256
rect 270493 8198 272504 8200
rect 262305 8195 262371 8198
rect 270493 8195 270559 8198
rect 34744 8192 35060 8193
rect 34744 8128 34750 8192
rect 34814 8128 34830 8192
rect 34894 8128 34910 8192
rect 34974 8128 34990 8192
rect 35054 8128 35060 8192
rect 34744 8127 35060 8128
rect 102341 8192 102657 8193
rect 102341 8128 102347 8192
rect 102411 8128 102427 8192
rect 102491 8128 102507 8192
rect 102571 8128 102587 8192
rect 102651 8128 102657 8192
rect 102341 8127 102657 8128
rect 169938 8192 170254 8193
rect 169938 8128 169944 8192
rect 170008 8128 170024 8192
rect 170088 8128 170104 8192
rect 170168 8128 170184 8192
rect 170248 8128 170254 8192
rect 169938 8127 170254 8128
rect 237535 8192 237851 8193
rect 237535 8128 237541 8192
rect 237605 8128 237621 8192
rect 237685 8128 237701 8192
rect 237765 8128 237781 8192
rect 237845 8128 237851 8192
rect 237535 8127 237851 8128
rect 88926 8060 88932 8124
rect 88996 8122 89002 8124
rect 89713 8122 89779 8125
rect 88996 8120 89779 8122
rect 88996 8064 89718 8120
rect 89774 8064 89779 8120
rect 88996 8062 89779 8064
rect 88996 8060 89002 8062
rect 89713 8059 89779 8062
rect 168230 8060 168236 8124
rect 168300 8122 168306 8124
rect 168373 8122 168439 8125
rect 168300 8120 168439 8122
rect 168300 8064 168378 8120
rect 168434 8064 168439 8120
rect 168300 8062 168439 8064
rect 168300 8060 168306 8062
rect 168373 8059 168439 8062
rect 187693 8122 187759 8125
rect 227621 8122 227687 8125
rect 187693 8120 227687 8122
rect 187693 8064 187698 8120
rect 187754 8064 227626 8120
rect 227682 8064 227687 8120
rect 187693 8062 227687 8064
rect 187693 8059 187759 8062
rect 227621 8059 227687 8062
rect 237925 8122 237991 8125
rect 268929 8122 268995 8125
rect 237925 8120 268995 8122
rect 237925 8064 237930 8120
rect 237986 8064 268934 8120
rect 268990 8064 268995 8120
rect 237925 8062 268995 8064
rect 237925 8059 237991 8062
rect 268929 8059 268995 8062
rect 270309 8122 270375 8125
rect 270309 8120 272504 8122
rect 270309 8064 270314 8120
rect 270370 8064 272504 8120
rect 270309 8062 272504 8064
rect 270309 8059 270375 8062
rect 84101 7986 84167 7989
rect 114829 7986 114895 7989
rect 84101 7984 114895 7986
rect 84101 7928 84106 7984
rect 84162 7928 114834 7984
rect 114890 7928 114895 7984
rect 84101 7926 114895 7928
rect 84101 7923 84167 7926
rect 114829 7923 114895 7926
rect 151353 7986 151419 7989
rect 173433 7986 173499 7989
rect 151353 7984 173499 7986
rect 151353 7928 151358 7984
rect 151414 7928 173438 7984
rect 173494 7928 173499 7984
rect 151353 7926 173499 7928
rect 151353 7923 151419 7926
rect 173433 7923 173499 7926
rect 194409 7986 194475 7989
rect 237649 7986 237715 7989
rect 194409 7984 237715 7986
rect 194409 7928 194414 7984
rect 194470 7928 237654 7984
rect 237710 7928 237715 7984
rect 194409 7926 237715 7928
rect 194409 7923 194475 7926
rect 237649 7923 237715 7926
rect 237833 7986 237899 7989
rect 268745 7986 268811 7989
rect 237833 7984 268811 7986
rect 237833 7928 237838 7984
rect 237894 7928 268750 7984
rect 268806 7928 268811 7984
rect 237833 7926 268811 7928
rect 237833 7923 237899 7926
rect 268745 7923 268811 7926
rect 270125 7986 270191 7989
rect 270125 7984 272504 7986
rect 270125 7928 270130 7984
rect 270186 7928 272504 7984
rect 270125 7926 272504 7928
rect 270125 7923 270191 7926
rect 27286 7788 27292 7852
rect 27356 7850 27362 7852
rect 27889 7850 27955 7853
rect 27356 7848 27955 7850
rect 27356 7792 27894 7848
rect 27950 7792 27955 7848
rect 27356 7790 27955 7792
rect 27356 7788 27362 7790
rect 27889 7787 27955 7790
rect 82721 7850 82787 7853
rect 114737 7850 114803 7853
rect 82721 7848 114803 7850
rect 82721 7792 82726 7848
rect 82782 7792 114742 7848
rect 114798 7792 114803 7848
rect 82721 7790 114803 7792
rect 82721 7787 82787 7790
rect 114737 7787 114803 7790
rect 154113 7850 154179 7853
rect 177941 7850 178007 7853
rect 154113 7848 178007 7850
rect 154113 7792 154118 7848
rect 154174 7792 177946 7848
rect 178002 7792 178007 7848
rect 154113 7790 178007 7792
rect 154113 7787 154179 7790
rect 177941 7787 178007 7790
rect 197169 7850 197235 7853
rect 220629 7850 220695 7853
rect 197169 7848 220695 7850
rect 197169 7792 197174 7848
rect 197230 7792 220634 7848
rect 220690 7792 220695 7848
rect 197169 7790 220695 7792
rect 197169 7787 197235 7790
rect 220629 7787 220695 7790
rect 224309 7850 224375 7853
rect 229737 7850 229803 7853
rect 224309 7848 229803 7850
rect 224309 7792 224314 7848
rect 224370 7792 229742 7848
rect 229798 7792 229803 7848
rect 224309 7790 229803 7792
rect 224309 7787 224375 7790
rect 229737 7787 229803 7790
rect 237005 7850 237071 7853
rect 237925 7850 237991 7853
rect 237005 7848 237991 7850
rect 237005 7792 237010 7848
rect 237066 7792 237930 7848
rect 237986 7792 237991 7848
rect 237005 7790 237991 7792
rect 237005 7787 237071 7790
rect 237925 7787 237991 7790
rect 238937 7850 239003 7853
rect 267273 7850 267339 7853
rect 267825 7850 267891 7853
rect 238937 7848 267891 7850
rect 238937 7792 238942 7848
rect 238998 7792 267278 7848
rect 267334 7792 267830 7848
rect 267886 7792 267891 7848
rect 238937 7790 267891 7792
rect 238937 7787 239003 7790
rect 267273 7787 267339 7790
rect 267825 7787 267891 7790
rect 268009 7850 268075 7853
rect 268009 7848 272504 7850
rect 268009 7792 268014 7848
rect 268070 7792 272504 7848
rect 268009 7790 272504 7792
rect 268009 7787 268075 7790
rect 86585 7714 86651 7717
rect 118969 7714 119035 7717
rect 86585 7712 119035 7714
rect 86585 7656 86590 7712
rect 86646 7656 118974 7712
rect 119030 7656 119035 7712
rect 86585 7654 119035 7656
rect 86585 7651 86651 7654
rect 118969 7651 119035 7654
rect 146569 7714 146635 7717
rect 178033 7714 178099 7717
rect 146569 7712 178099 7714
rect 146569 7656 146574 7712
rect 146630 7656 178038 7712
rect 178094 7656 178099 7712
rect 146569 7654 178099 7656
rect 146569 7651 146635 7654
rect 178033 7651 178099 7654
rect 214833 7714 214899 7717
rect 242985 7714 243051 7717
rect 265801 7714 265867 7717
rect 267406 7714 267412 7716
rect 214833 7712 243051 7714
rect 214833 7656 214838 7712
rect 214894 7656 242990 7712
rect 243046 7656 243051 7712
rect 214833 7654 243051 7656
rect 214833 7651 214899 7654
rect 242985 7651 243051 7654
rect 244230 7654 248430 7714
rect 68542 7648 68858 7649
rect 68542 7584 68548 7648
rect 68612 7584 68628 7648
rect 68692 7584 68708 7648
rect 68772 7584 68788 7648
rect 68852 7584 68858 7648
rect 68542 7583 68858 7584
rect 136139 7648 136455 7649
rect 136139 7584 136145 7648
rect 136209 7584 136225 7648
rect 136289 7584 136305 7648
rect 136369 7584 136385 7648
rect 136449 7584 136455 7648
rect 136139 7583 136455 7584
rect 203736 7648 204052 7649
rect 203736 7584 203742 7648
rect 203806 7584 203822 7648
rect 203886 7584 203902 7648
rect 203966 7584 203982 7648
rect 204046 7584 204052 7648
rect 203736 7583 204052 7584
rect 87045 7578 87111 7581
rect 120349 7578 120415 7581
rect 87045 7576 120415 7578
rect 87045 7520 87050 7576
rect 87106 7520 120354 7576
rect 120410 7520 120415 7576
rect 87045 7518 120415 7520
rect 87045 7515 87111 7518
rect 120349 7515 120415 7518
rect 144545 7578 144611 7581
rect 176837 7578 176903 7581
rect 144545 7576 176903 7578
rect 144545 7520 144550 7576
rect 144606 7520 176842 7576
rect 176898 7520 176903 7576
rect 144545 7518 176903 7520
rect 144545 7515 144611 7518
rect 176837 7515 176903 7518
rect 223849 7578 223915 7581
rect 224953 7578 225019 7581
rect 223849 7576 225019 7578
rect 223849 7520 223854 7576
rect 223910 7520 224958 7576
rect 225014 7520 225019 7576
rect 223849 7518 225019 7520
rect 223849 7515 223915 7518
rect 224953 7515 225019 7518
rect 229737 7578 229803 7581
rect 238753 7578 238819 7581
rect 229737 7576 238819 7578
rect 229737 7520 229742 7576
rect 229798 7520 238758 7576
rect 238814 7520 238819 7576
rect 229737 7518 238819 7520
rect 229737 7515 229803 7518
rect 238753 7515 238819 7518
rect 239029 7578 239095 7581
rect 244230 7578 244290 7654
rect 239029 7576 244290 7578
rect 239029 7520 239034 7576
rect 239090 7520 244290 7576
rect 239029 7518 244290 7520
rect 248370 7578 248430 7654
rect 253890 7712 267412 7714
rect 253890 7656 265806 7712
rect 265862 7656 267412 7712
rect 253890 7654 267412 7656
rect 253890 7578 253950 7654
rect 265801 7651 265867 7654
rect 267406 7652 267412 7654
rect 267476 7714 267482 7716
rect 267641 7714 267707 7717
rect 267476 7712 267707 7714
rect 267476 7656 267646 7712
rect 267702 7656 267707 7712
rect 267476 7654 267707 7656
rect 267476 7652 267482 7654
rect 267641 7651 267707 7654
rect 271781 7714 271847 7717
rect 271781 7712 272504 7714
rect 271781 7656 271786 7712
rect 271842 7656 272504 7712
rect 271781 7654 272504 7656
rect 271781 7651 271847 7654
rect 271333 7648 271649 7649
rect 271333 7584 271339 7648
rect 271403 7584 271419 7648
rect 271483 7584 271499 7648
rect 271563 7584 271579 7648
rect 271643 7584 271649 7648
rect 271333 7583 271649 7584
rect 248370 7518 253950 7578
rect 263777 7578 263843 7581
rect 265985 7578 266051 7581
rect 263777 7576 266051 7578
rect 263777 7520 263782 7576
rect 263838 7520 265990 7576
rect 266046 7520 266051 7576
rect 263777 7518 266051 7520
rect 239029 7515 239095 7518
rect 263777 7515 263843 7518
rect 265985 7515 266051 7518
rect 266169 7578 266235 7581
rect 267641 7578 267707 7581
rect 266169 7576 267707 7578
rect 266169 7520 266174 7576
rect 266230 7520 267646 7576
rect 267702 7520 267707 7576
rect 266169 7518 267707 7520
rect 266169 7515 266235 7518
rect 267641 7515 267707 7518
rect 267958 7516 267964 7580
rect 268028 7578 268034 7580
rect 271137 7578 271203 7581
rect 268028 7576 271203 7578
rect 268028 7520 271142 7576
rect 271198 7520 271203 7576
rect 268028 7518 271203 7520
rect 268028 7516 268034 7518
rect 271137 7515 271203 7518
rect 271781 7578 271847 7581
rect 271781 7576 272504 7578
rect 271781 7520 271786 7576
rect 271842 7520 272504 7576
rect 271781 7518 272504 7520
rect 271781 7515 271847 7518
rect 82629 7442 82695 7445
rect 112345 7442 112411 7445
rect 82629 7440 112411 7442
rect 82629 7384 82634 7440
rect 82690 7384 112350 7440
rect 112406 7384 112411 7440
rect 82629 7382 112411 7384
rect 82629 7379 82695 7382
rect 112345 7379 112411 7382
rect 130285 7442 130351 7445
rect 230289 7442 230355 7445
rect 130285 7440 230355 7442
rect 130285 7384 130290 7440
rect 130346 7384 230294 7440
rect 230350 7384 230355 7440
rect 130285 7382 230355 7384
rect 130285 7379 130351 7382
rect 230289 7379 230355 7382
rect 237281 7442 237347 7445
rect 268009 7442 268075 7445
rect 237281 7440 253950 7442
rect 237281 7384 237286 7440
rect 237342 7384 253950 7440
rect 237281 7382 253950 7384
rect 237281 7379 237347 7382
rect 163681 7306 163747 7309
rect 220813 7306 220879 7309
rect 163681 7304 220879 7306
rect 163681 7248 163686 7304
rect 163742 7248 220818 7304
rect 220874 7248 220879 7304
rect 163681 7246 220879 7248
rect 163681 7243 163747 7246
rect 220813 7243 220879 7246
rect 221365 7306 221431 7309
rect 221917 7306 221983 7309
rect 221365 7304 221983 7306
rect 221365 7248 221370 7304
rect 221426 7248 221922 7304
rect 221978 7248 221983 7304
rect 221365 7246 221983 7248
rect 221365 7243 221431 7246
rect 221917 7243 221983 7246
rect 222193 7306 222259 7309
rect 248965 7306 249031 7309
rect 222193 7304 249031 7306
rect 222193 7248 222198 7304
rect 222254 7248 248970 7304
rect 249026 7248 249031 7304
rect 222193 7246 249031 7248
rect 253890 7306 253950 7382
rect 268009 7440 272504 7442
rect 268009 7384 268014 7440
rect 268070 7384 272504 7440
rect 268009 7382 272504 7384
rect 268009 7379 268075 7382
rect 267733 7306 267799 7309
rect 253890 7304 267799 7306
rect 253890 7248 267738 7304
rect 267794 7248 267799 7304
rect 253890 7246 267799 7248
rect 222193 7243 222259 7246
rect 248965 7243 249031 7246
rect 267733 7243 267799 7246
rect 268009 7306 268075 7309
rect 271781 7306 271847 7309
rect 268009 7304 271847 7306
rect 268009 7248 268014 7304
rect 268070 7248 271786 7304
rect 271842 7248 271847 7304
rect 268009 7246 271847 7248
rect 268009 7243 268075 7246
rect 271781 7243 271847 7246
rect 271965 7306 272031 7309
rect 271965 7304 272504 7306
rect 271965 7248 271970 7304
rect 272026 7248 272504 7304
rect 271965 7246 272504 7248
rect 271965 7243 272031 7246
rect 177941 7170 178007 7173
rect 215569 7170 215635 7173
rect 218513 7170 218579 7173
rect 177941 7168 195990 7170
rect 177941 7112 177946 7168
rect 178002 7112 195990 7168
rect 177941 7110 195990 7112
rect 177941 7107 178007 7110
rect 34744 7104 35060 7105
rect 34744 7040 34750 7104
rect 34814 7040 34830 7104
rect 34894 7040 34910 7104
rect 34974 7040 34990 7104
rect 35054 7040 35060 7104
rect 34744 7039 35060 7040
rect 102341 7104 102657 7105
rect 102341 7040 102347 7104
rect 102411 7040 102427 7104
rect 102491 7040 102507 7104
rect 102571 7040 102587 7104
rect 102651 7040 102657 7104
rect 102341 7039 102657 7040
rect 169938 7104 170254 7105
rect 169938 7040 169944 7104
rect 170008 7040 170024 7104
rect 170088 7040 170104 7104
rect 170168 7040 170184 7104
rect 170248 7040 170254 7104
rect 169938 7039 170254 7040
rect 195930 7034 195990 7110
rect 215569 7168 218579 7170
rect 215569 7112 215574 7168
rect 215630 7112 218518 7168
rect 218574 7112 218579 7168
rect 215569 7110 218579 7112
rect 215569 7107 215635 7110
rect 218513 7107 218579 7110
rect 218697 7170 218763 7173
rect 219709 7170 219775 7173
rect 218697 7168 219775 7170
rect 218697 7112 218702 7168
rect 218758 7112 219714 7168
rect 219770 7112 219775 7168
rect 218697 7110 219775 7112
rect 218697 7107 218763 7110
rect 219709 7107 219775 7110
rect 220905 7170 220971 7173
rect 237189 7170 237255 7173
rect 220905 7168 237255 7170
rect 220905 7112 220910 7168
rect 220966 7112 237194 7168
rect 237250 7112 237255 7168
rect 220905 7110 237255 7112
rect 220905 7107 220971 7110
rect 237189 7107 237255 7110
rect 262489 7170 262555 7173
rect 262489 7168 272504 7170
rect 262489 7112 262494 7168
rect 262550 7112 272504 7168
rect 262489 7110 272504 7112
rect 262489 7107 262555 7110
rect 237535 7104 237851 7105
rect 237535 7040 237541 7104
rect 237605 7040 237621 7104
rect 237685 7040 237701 7104
rect 237765 7040 237781 7104
rect 237845 7040 237851 7104
rect 237535 7039 237851 7040
rect 215293 7034 215359 7037
rect 224861 7034 224927 7037
rect 195930 7032 215359 7034
rect 195930 6976 215298 7032
rect 215354 6976 215359 7032
rect 195930 6974 215359 6976
rect 215293 6971 215359 6974
rect 216584 7032 224927 7034
rect 216584 6976 224866 7032
rect 224922 6976 224927 7032
rect 216584 6974 224927 6976
rect 19241 6900 19307 6901
rect 19977 6900 20043 6901
rect 19190 6898 19196 6900
rect 19150 6838 19196 6898
rect 19260 6896 19307 6900
rect 19926 6898 19932 6900
rect 19302 6840 19307 6896
rect 19190 6836 19196 6838
rect 19260 6836 19307 6840
rect 19886 6838 19932 6898
rect 19996 6896 20043 6900
rect 20038 6840 20043 6896
rect 19926 6836 19932 6838
rect 19996 6836 20043 6840
rect 22870 6836 22876 6900
rect 22940 6898 22946 6900
rect 23473 6898 23539 6901
rect 22940 6896 23539 6898
rect 22940 6840 23478 6896
rect 23534 6840 23539 6896
rect 22940 6838 23539 6840
rect 22940 6836 22946 6838
rect 19241 6835 19307 6836
rect 19977 6835 20043 6836
rect 23473 6835 23539 6838
rect 23606 6836 23612 6900
rect 23676 6898 23682 6900
rect 24761 6898 24827 6901
rect 23676 6896 24827 6898
rect 23676 6840 24766 6896
rect 24822 6840 24827 6896
rect 23676 6838 24827 6840
rect 23676 6836 23682 6838
rect 24761 6835 24827 6838
rect 25078 6836 25084 6900
rect 25148 6898 25154 6900
rect 26233 6898 26299 6901
rect 25148 6896 26299 6898
rect 25148 6840 26238 6896
rect 26294 6840 26299 6896
rect 25148 6838 26299 6840
rect 25148 6836 25154 6838
rect 26233 6835 26299 6838
rect 101857 6898 101923 6901
rect 101857 6896 109050 6898
rect 101857 6840 101862 6896
rect 101918 6840 109050 6896
rect 101857 6838 109050 6840
rect 101857 6835 101923 6838
rect 79317 6762 79383 6765
rect 100109 6762 100175 6765
rect 108990 6762 109050 6838
rect 212206 6836 212212 6900
rect 212276 6898 212282 6900
rect 212441 6898 212507 6901
rect 212276 6896 212507 6898
rect 212276 6840 212446 6896
rect 212502 6840 212507 6896
rect 212276 6838 212507 6840
rect 212276 6836 212282 6838
rect 212441 6835 212507 6838
rect 215017 6898 215083 6901
rect 216584 6898 216644 6974
rect 224861 6971 224927 6974
rect 268009 7034 268075 7037
rect 268009 7032 272504 7034
rect 268009 6976 268014 7032
rect 268070 6976 272504 7032
rect 268009 6974 272504 6976
rect 268009 6971 268075 6974
rect 215017 6896 216644 6898
rect 215017 6840 215022 6896
rect 215078 6840 216644 6896
rect 215017 6838 216644 6840
rect 216765 6898 216831 6901
rect 219617 6898 219683 6901
rect 216765 6896 219683 6898
rect 216765 6840 216770 6896
rect 216826 6840 219622 6896
rect 219678 6840 219683 6896
rect 216765 6838 219683 6840
rect 215017 6835 215083 6838
rect 216765 6835 216831 6838
rect 219617 6835 219683 6838
rect 220629 6898 220695 6901
rect 224953 6898 225019 6901
rect 220629 6896 225019 6898
rect 220629 6840 220634 6896
rect 220690 6840 224958 6896
rect 225014 6840 225019 6896
rect 220629 6838 225019 6840
rect 220629 6835 220695 6838
rect 224953 6835 225019 6838
rect 237005 6898 237071 6901
rect 243813 6898 243879 6901
rect 237005 6896 243879 6898
rect 237005 6840 237010 6896
rect 237066 6840 243818 6896
rect 243874 6840 243879 6896
rect 237005 6838 243879 6840
rect 237005 6835 237071 6838
rect 243813 6835 243879 6838
rect 265341 6898 265407 6901
rect 267089 6898 267155 6901
rect 265341 6896 267155 6898
rect 265341 6840 265346 6896
rect 265402 6840 267094 6896
rect 267150 6840 267155 6896
rect 265341 6838 267155 6840
rect 265341 6835 265407 6838
rect 267089 6835 267155 6838
rect 268101 6898 268167 6901
rect 268101 6896 272504 6898
rect 268101 6840 268106 6896
rect 268162 6840 272504 6896
rect 268101 6838 272504 6840
rect 268101 6835 268167 6838
rect 113173 6762 113239 6765
rect 79317 6760 102794 6762
rect 79317 6704 79322 6760
rect 79378 6704 100114 6760
rect 100170 6704 102794 6760
rect 79317 6702 102794 6704
rect 108990 6760 113239 6762
rect 108990 6704 113178 6760
rect 113234 6704 113239 6760
rect 108990 6702 113239 6704
rect 79317 6699 79383 6702
rect 100109 6699 100175 6702
rect 86585 6626 86651 6629
rect 102225 6626 102291 6629
rect 86585 6624 102291 6626
rect 86585 6568 86590 6624
rect 86646 6568 102230 6624
rect 102286 6568 102291 6624
rect 86585 6566 102291 6568
rect 102734 6626 102794 6702
rect 113173 6699 113239 6702
rect 156045 6762 156111 6765
rect 215569 6762 215635 6765
rect 156045 6760 215635 6762
rect 156045 6704 156050 6760
rect 156106 6704 215574 6760
rect 215630 6704 215635 6760
rect 156045 6702 215635 6704
rect 156045 6699 156111 6702
rect 215569 6699 215635 6702
rect 218881 6762 218947 6765
rect 251449 6762 251515 6765
rect 218881 6760 251515 6762
rect 218881 6704 218886 6760
rect 218942 6704 251454 6760
rect 251510 6704 251515 6760
rect 218881 6702 251515 6704
rect 218881 6699 218947 6702
rect 251449 6699 251515 6702
rect 264145 6762 264211 6765
rect 266118 6762 266124 6764
rect 264145 6760 266124 6762
rect 264145 6704 264150 6760
rect 264206 6704 266124 6760
rect 264145 6702 266124 6704
rect 264145 6699 264211 6702
rect 266118 6700 266124 6702
rect 266188 6700 266194 6764
rect 267590 6700 267596 6764
rect 267660 6762 267666 6764
rect 271689 6762 271755 6765
rect 267660 6760 271755 6762
rect 267660 6704 271694 6760
rect 271750 6704 271755 6760
rect 267660 6702 271755 6704
rect 267660 6700 267666 6702
rect 271689 6699 271755 6702
rect 272057 6762 272123 6765
rect 272057 6760 272504 6762
rect 272057 6704 272062 6760
rect 272118 6704 272504 6760
rect 272057 6702 272504 6704
rect 272057 6699 272123 6702
rect 152641 6626 152707 6629
rect 177941 6626 178007 6629
rect 102734 6566 109050 6626
rect 86585 6563 86651 6566
rect 102225 6563 102291 6566
rect 68542 6560 68858 6561
rect 68542 6496 68548 6560
rect 68612 6496 68628 6560
rect 68692 6496 68708 6560
rect 68772 6496 68788 6560
rect 68852 6496 68858 6560
rect 68542 6495 68858 6496
rect 35893 6490 35959 6493
rect 46013 6490 46079 6493
rect 35893 6488 46079 6490
rect 35893 6432 35898 6488
rect 35954 6432 46018 6488
rect 46074 6432 46079 6488
rect 35893 6430 46079 6432
rect 108990 6490 109050 6566
rect 152641 6624 178007 6626
rect 152641 6568 152646 6624
rect 152702 6568 177946 6624
rect 178002 6568 178007 6624
rect 152641 6566 178007 6568
rect 152641 6563 152707 6566
rect 177941 6563 178007 6566
rect 216622 6564 216628 6628
rect 216692 6626 216698 6628
rect 231485 6626 231551 6629
rect 231761 6626 231827 6629
rect 216692 6624 231827 6626
rect 216692 6568 231490 6624
rect 231546 6568 231766 6624
rect 231822 6568 231827 6624
rect 216692 6566 231827 6568
rect 216692 6564 216698 6566
rect 231485 6563 231551 6566
rect 231761 6563 231827 6566
rect 242893 6626 242959 6629
rect 263409 6626 263475 6629
rect 269021 6626 269087 6629
rect 242893 6624 258826 6626
rect 242893 6568 242898 6624
rect 242954 6568 258826 6624
rect 242893 6566 258826 6568
rect 242893 6563 242959 6566
rect 136139 6560 136455 6561
rect 136139 6496 136145 6560
rect 136209 6496 136225 6560
rect 136289 6496 136305 6560
rect 136369 6496 136385 6560
rect 136449 6496 136455 6560
rect 136139 6495 136455 6496
rect 203736 6560 204052 6561
rect 203736 6496 203742 6560
rect 203806 6496 203822 6560
rect 203886 6496 203902 6560
rect 203966 6496 203982 6560
rect 204046 6496 204052 6560
rect 203736 6495 204052 6496
rect 115933 6490 115999 6493
rect 180057 6490 180123 6493
rect 108990 6488 115999 6490
rect 108990 6432 115938 6488
rect 115994 6432 115999 6488
rect 108990 6430 115999 6432
rect 35893 6427 35959 6430
rect 46013 6427 46079 6430
rect 115933 6427 115999 6430
rect 152782 6488 180123 6490
rect 152782 6432 180062 6488
rect 180118 6432 180123 6488
rect 152782 6430 180123 6432
rect 95233 6354 95299 6357
rect 112713 6354 112779 6357
rect 152641 6354 152707 6357
rect 95233 6352 152707 6354
rect 95233 6296 95238 6352
rect 95294 6296 112718 6352
rect 112774 6296 152646 6352
rect 152702 6296 152707 6352
rect 95233 6294 152707 6296
rect 95233 6291 95299 6294
rect 112713 6291 112779 6294
rect 152641 6291 152707 6294
rect 44081 6218 44147 6221
rect 92657 6218 92723 6221
rect 44081 6216 92723 6218
rect 44081 6160 44086 6216
rect 44142 6160 92662 6216
rect 92718 6160 92723 6216
rect 44081 6158 92723 6160
rect 44081 6155 44147 6158
rect 92657 6155 92723 6158
rect 94497 6218 94563 6221
rect 108665 6218 108731 6221
rect 148133 6218 148199 6221
rect 152782 6218 152842 6430
rect 180057 6427 180123 6430
rect 219985 6490 220051 6493
rect 226241 6490 226307 6493
rect 219985 6488 226307 6490
rect 219985 6432 219990 6488
rect 220046 6432 226246 6488
rect 226302 6432 226307 6488
rect 219985 6430 226307 6432
rect 219985 6427 220051 6430
rect 226241 6427 226307 6430
rect 230381 6490 230447 6493
rect 230381 6488 253950 6490
rect 230381 6432 230386 6488
rect 230442 6432 253950 6488
rect 230381 6430 253950 6432
rect 230381 6427 230447 6430
rect 162761 6354 162827 6357
rect 170581 6354 170647 6357
rect 162761 6352 170647 6354
rect 162761 6296 162766 6352
rect 162822 6296 170586 6352
rect 170642 6296 170647 6352
rect 162761 6294 170647 6296
rect 162761 6291 162827 6294
rect 170581 6291 170647 6294
rect 177021 6354 177087 6357
rect 214557 6354 214623 6357
rect 177021 6352 214623 6354
rect 177021 6296 177026 6352
rect 177082 6296 214562 6352
rect 214618 6296 214623 6352
rect 177021 6294 214623 6296
rect 177021 6291 177087 6294
rect 214557 6291 214623 6294
rect 221365 6354 221431 6357
rect 252553 6354 252619 6357
rect 221365 6352 252619 6354
rect 221365 6296 221370 6352
rect 221426 6296 252558 6352
rect 252614 6296 252619 6352
rect 221365 6294 252619 6296
rect 221365 6291 221431 6294
rect 252553 6291 252619 6294
rect 182909 6218 182975 6221
rect 94497 6216 152842 6218
rect 94497 6160 94502 6216
rect 94558 6160 108670 6216
rect 108726 6160 148138 6216
rect 148194 6160 152842 6216
rect 94497 6158 152842 6160
rect 157290 6216 182975 6218
rect 157290 6160 182914 6216
rect 182970 6160 182975 6216
rect 157290 6158 182975 6160
rect 94497 6155 94563 6158
rect 108665 6155 108731 6158
rect 148133 6155 148199 6158
rect 150249 6082 150315 6085
rect 157290 6082 157350 6158
rect 182909 6155 182975 6158
rect 218973 6218 219039 6221
rect 221457 6218 221523 6221
rect 221733 6218 221799 6221
rect 222101 6218 222167 6221
rect 218973 6216 222167 6218
rect 218973 6160 218978 6216
rect 219034 6160 221462 6216
rect 221518 6160 221738 6216
rect 221794 6160 222106 6216
rect 222162 6160 222167 6216
rect 218973 6158 222167 6160
rect 218973 6155 219039 6158
rect 221457 6155 221523 6158
rect 221733 6155 221799 6158
rect 222101 6155 222167 6158
rect 223389 6218 223455 6221
rect 224125 6218 224191 6221
rect 223389 6216 224191 6218
rect 223389 6160 223394 6216
rect 223450 6160 224130 6216
rect 224186 6160 224191 6216
rect 223389 6158 224191 6160
rect 223389 6155 223455 6158
rect 224125 6155 224191 6158
rect 224861 6218 224927 6221
rect 225597 6218 225663 6221
rect 224861 6216 225663 6218
rect 224861 6160 224866 6216
rect 224922 6160 225602 6216
rect 225658 6160 225663 6216
rect 224861 6158 225663 6160
rect 224861 6155 224927 6158
rect 225597 6155 225663 6158
rect 226333 6218 226399 6221
rect 249609 6218 249675 6221
rect 226333 6216 249675 6218
rect 226333 6160 226338 6216
rect 226394 6160 249614 6216
rect 249670 6160 249675 6216
rect 226333 6158 249675 6160
rect 253890 6218 253950 6430
rect 258766 6354 258826 6566
rect 263409 6624 269087 6626
rect 263409 6568 263414 6624
rect 263470 6568 269026 6624
rect 269082 6568 269087 6624
rect 263409 6566 269087 6568
rect 263409 6563 263475 6566
rect 269021 6563 269087 6566
rect 271873 6626 271939 6629
rect 271873 6624 272504 6626
rect 271873 6568 271878 6624
rect 271934 6568 272504 6624
rect 271873 6566 272504 6568
rect 271873 6563 271939 6566
rect 271333 6560 271649 6561
rect 271333 6496 271339 6560
rect 271403 6496 271419 6560
rect 271483 6496 271499 6560
rect 271563 6496 271579 6560
rect 271643 6496 271649 6560
rect 271333 6495 271649 6496
rect 263409 6490 263475 6493
rect 268193 6490 268259 6493
rect 263409 6488 268259 6490
rect 263409 6432 263414 6488
rect 263470 6432 268198 6488
rect 268254 6432 268259 6488
rect 263409 6430 268259 6432
rect 263409 6427 263475 6430
rect 268193 6427 268259 6430
rect 268745 6490 268811 6493
rect 268745 6488 270970 6490
rect 268745 6432 268750 6488
rect 268806 6432 270970 6488
rect 268745 6430 270970 6432
rect 268745 6427 268811 6430
rect 268377 6354 268443 6357
rect 269113 6354 269179 6357
rect 258766 6352 269179 6354
rect 258766 6296 268382 6352
rect 268438 6296 269118 6352
rect 269174 6296 269179 6352
rect 258766 6294 269179 6296
rect 270910 6354 270970 6430
rect 271830 6430 272504 6490
rect 271830 6354 271890 6430
rect 270910 6294 271890 6354
rect 271965 6354 272031 6357
rect 271965 6352 272504 6354
rect 271965 6296 271970 6352
rect 272026 6296 272504 6352
rect 271965 6294 272504 6296
rect 268377 6291 268443 6294
rect 269113 6291 269179 6294
rect 271965 6291 272031 6294
rect 261477 6218 261543 6221
rect 262070 6218 262076 6220
rect 253890 6216 262076 6218
rect 253890 6160 261482 6216
rect 261538 6160 262076 6216
rect 253890 6158 262076 6160
rect 226333 6155 226399 6158
rect 249609 6155 249675 6158
rect 261477 6155 261543 6158
rect 262070 6156 262076 6158
rect 262140 6156 262146 6220
rect 267273 6218 267339 6221
rect 268142 6218 268148 6220
rect 267273 6216 268148 6218
rect 267273 6160 267278 6216
rect 267334 6160 268148 6216
rect 267273 6158 268148 6160
rect 267273 6155 267339 6158
rect 268142 6156 268148 6158
rect 268212 6156 268218 6220
rect 268929 6218 268995 6221
rect 268929 6216 272504 6218
rect 268929 6160 268934 6216
rect 268990 6160 272504 6216
rect 268929 6158 272504 6160
rect 268929 6155 268995 6158
rect 150249 6080 157350 6082
rect 150249 6024 150254 6080
rect 150310 6024 157350 6080
rect 150249 6022 157350 6024
rect 182081 6082 182147 6085
rect 228081 6082 228147 6085
rect 182081 6080 228147 6082
rect 182081 6024 182086 6080
rect 182142 6024 228086 6080
rect 228142 6024 228147 6080
rect 182081 6022 228147 6024
rect 150249 6019 150315 6022
rect 182081 6019 182147 6022
rect 228081 6019 228147 6022
rect 269021 6082 269087 6085
rect 271781 6082 271847 6085
rect 269021 6080 271522 6082
rect 269021 6024 269026 6080
rect 269082 6024 271522 6080
rect 269021 6022 271522 6024
rect 269021 6019 269087 6022
rect 34744 6016 35060 6017
rect 34744 5952 34750 6016
rect 34814 5952 34830 6016
rect 34894 5952 34910 6016
rect 34974 5952 34990 6016
rect 35054 5952 35060 6016
rect 34744 5951 35060 5952
rect 102341 6016 102657 6017
rect 102341 5952 102347 6016
rect 102411 5952 102427 6016
rect 102491 5952 102507 6016
rect 102571 5952 102587 6016
rect 102651 5952 102657 6016
rect 102341 5951 102657 5952
rect 169938 6016 170254 6017
rect 169938 5952 169944 6016
rect 170008 5952 170024 6016
rect 170088 5952 170104 6016
rect 170168 5952 170184 6016
rect 170248 5952 170254 6016
rect 169938 5951 170254 5952
rect 237535 6016 237851 6017
rect 237535 5952 237541 6016
rect 237605 5952 237621 6016
rect 237685 5952 237701 6016
rect 237765 5952 237781 6016
rect 237845 5952 237851 6016
rect 237535 5951 237851 5952
rect 130193 5946 130259 5949
rect 188429 5946 188495 5949
rect 130193 5944 157350 5946
rect 130193 5888 130198 5944
rect 130254 5888 157350 5944
rect 130193 5886 157350 5888
rect 130193 5883 130259 5886
rect 43161 5810 43227 5813
rect 43621 5810 43687 5813
rect 45369 5810 45435 5813
rect 43161 5808 45435 5810
rect 43161 5752 43166 5808
rect 43222 5752 43626 5808
rect 43682 5752 45374 5808
rect 45430 5752 45435 5808
rect 43161 5750 45435 5752
rect 43161 5747 43227 5750
rect 43621 5747 43687 5750
rect 45369 5747 45435 5750
rect 81985 5810 82051 5813
rect 100569 5810 100635 5813
rect 81985 5808 100635 5810
rect 81985 5752 81990 5808
rect 82046 5752 100574 5808
rect 100630 5752 100635 5808
rect 81985 5750 100635 5752
rect 81985 5747 82051 5750
rect 100569 5747 100635 5750
rect 108849 5810 108915 5813
rect 111517 5810 111583 5813
rect 108849 5808 111583 5810
rect 108849 5752 108854 5808
rect 108910 5752 111522 5808
rect 111578 5752 111583 5808
rect 108849 5750 111583 5752
rect 157290 5810 157350 5886
rect 170446 5944 188495 5946
rect 170446 5888 188434 5944
rect 188490 5888 188495 5944
rect 170446 5886 188495 5888
rect 170446 5810 170506 5886
rect 188429 5883 188495 5886
rect 211153 5946 211219 5949
rect 237005 5946 237071 5949
rect 211153 5944 237071 5946
rect 211153 5888 211158 5944
rect 211214 5888 237010 5944
rect 237066 5888 237071 5944
rect 211153 5886 237071 5888
rect 211153 5883 211219 5886
rect 237005 5883 237071 5886
rect 263041 5946 263107 5949
rect 268193 5946 268259 5949
rect 263041 5944 268259 5946
rect 263041 5888 263046 5944
rect 263102 5888 268198 5944
rect 268254 5888 268259 5944
rect 263041 5886 268259 5888
rect 263041 5883 263107 5886
rect 268193 5883 268259 5886
rect 268469 5946 268535 5949
rect 268469 5944 271338 5946
rect 268469 5888 268474 5944
rect 268530 5888 271338 5944
rect 268469 5886 271338 5888
rect 268469 5883 268535 5886
rect 157290 5750 170506 5810
rect 170581 5810 170647 5813
rect 231669 5810 231735 5813
rect 232313 5810 232379 5813
rect 251817 5810 251883 5813
rect 262305 5810 262371 5813
rect 170581 5808 232379 5810
rect 170581 5752 170586 5808
rect 170642 5752 231674 5808
rect 231730 5752 232318 5808
rect 232374 5752 232379 5808
rect 170581 5750 232379 5752
rect 108849 5747 108915 5750
rect 111517 5747 111583 5750
rect 170581 5747 170647 5750
rect 231669 5747 231735 5750
rect 232313 5747 232379 5750
rect 234570 5808 251883 5810
rect 234570 5752 251822 5808
rect 251878 5752 251883 5808
rect 234570 5750 251883 5752
rect 42701 5674 42767 5677
rect 43713 5674 43779 5677
rect 42701 5672 43779 5674
rect 42701 5616 42706 5672
rect 42762 5616 43718 5672
rect 43774 5616 43779 5672
rect 42701 5614 43779 5616
rect 42701 5611 42767 5614
rect 43713 5611 43779 5614
rect 44541 5674 44607 5677
rect 81893 5674 81959 5677
rect 44541 5672 81959 5674
rect 44541 5616 44546 5672
rect 44602 5616 81898 5672
rect 81954 5616 81959 5672
rect 44541 5614 81959 5616
rect 44541 5611 44607 5614
rect 81893 5611 81959 5614
rect 85573 5674 85639 5677
rect 119429 5674 119495 5677
rect 85573 5672 119495 5674
rect 85573 5616 85578 5672
rect 85634 5616 119434 5672
rect 119490 5616 119495 5672
rect 85573 5614 119495 5616
rect 85573 5611 85639 5614
rect 119429 5611 119495 5614
rect 143533 5674 143599 5677
rect 208393 5674 208459 5677
rect 143533 5672 208459 5674
rect 143533 5616 143538 5672
rect 143594 5616 208398 5672
rect 208454 5616 208459 5672
rect 143533 5614 208459 5616
rect 143533 5611 143599 5614
rect 208393 5611 208459 5614
rect 212533 5674 212599 5677
rect 214649 5674 214715 5677
rect 212533 5672 214715 5674
rect 212533 5616 212538 5672
rect 212594 5616 214654 5672
rect 214710 5616 214715 5672
rect 212533 5614 214715 5616
rect 212533 5611 212599 5614
rect 214649 5611 214715 5614
rect 216305 5674 216371 5677
rect 226333 5674 226399 5677
rect 216305 5672 226399 5674
rect 216305 5616 216310 5672
rect 216366 5616 226338 5672
rect 226394 5616 226399 5672
rect 216305 5614 226399 5616
rect 216305 5611 216371 5614
rect 226333 5611 226399 5614
rect 226609 5674 226675 5677
rect 234570 5674 234630 5750
rect 251817 5747 251883 5750
rect 253890 5808 262371 5810
rect 253890 5752 262310 5808
rect 262366 5752 262371 5808
rect 253890 5750 262371 5752
rect 226609 5672 234630 5674
rect 226609 5616 226614 5672
rect 226670 5616 234630 5672
rect 226609 5614 234630 5616
rect 235349 5674 235415 5677
rect 253890 5674 253950 5750
rect 262305 5747 262371 5750
rect 262949 5810 263015 5813
rect 267733 5810 267799 5813
rect 262949 5808 267799 5810
rect 262949 5752 262954 5808
rect 263010 5752 267738 5808
rect 267794 5752 267799 5808
rect 262949 5750 267799 5752
rect 262949 5747 263015 5750
rect 267733 5747 267799 5750
rect 268009 5810 268075 5813
rect 270309 5810 270375 5813
rect 268009 5808 270375 5810
rect 268009 5752 268014 5808
rect 268070 5752 270314 5808
rect 270370 5752 270375 5808
rect 268009 5750 270375 5752
rect 268009 5747 268075 5750
rect 270309 5747 270375 5750
rect 270585 5810 270651 5813
rect 271086 5810 271092 5812
rect 270585 5808 271092 5810
rect 270585 5752 270590 5808
rect 270646 5752 271092 5808
rect 270585 5750 271092 5752
rect 270585 5747 270651 5750
rect 271086 5748 271092 5750
rect 271156 5748 271162 5812
rect 263133 5674 263199 5677
rect 266905 5676 266971 5677
rect 235349 5672 253950 5674
rect 235349 5616 235354 5672
rect 235410 5616 253950 5672
rect 235349 5614 253950 5616
rect 262262 5672 263199 5674
rect 262262 5616 263138 5672
rect 263194 5616 263199 5672
rect 262262 5614 263199 5616
rect 226609 5611 226675 5614
rect 235349 5611 235415 5614
rect 104893 5538 104959 5541
rect 117405 5538 117471 5541
rect 104893 5536 117471 5538
rect 104893 5480 104898 5536
rect 104954 5480 117410 5536
rect 117466 5480 117471 5536
rect 104893 5478 117471 5480
rect 104893 5475 104959 5478
rect 117405 5475 117471 5478
rect 215109 5538 215175 5541
rect 230606 5538 230612 5540
rect 215109 5536 230612 5538
rect 215109 5480 215114 5536
rect 215170 5480 230612 5536
rect 215109 5478 230612 5480
rect 215109 5475 215175 5478
rect 230606 5476 230612 5478
rect 230676 5476 230682 5540
rect 262262 5538 262322 5614
rect 263133 5611 263199 5614
rect 266854 5612 266860 5676
rect 266924 5674 266971 5676
rect 267733 5676 267799 5677
rect 267733 5674 267780 5676
rect 266924 5672 267016 5674
rect 266966 5616 267016 5672
rect 266924 5614 267016 5616
rect 267688 5672 267780 5674
rect 267688 5616 267738 5672
rect 267688 5614 267780 5616
rect 266924 5612 266971 5614
rect 266905 5611 266971 5612
rect 267733 5612 267780 5614
rect 267844 5612 267850 5676
rect 267917 5674 267983 5677
rect 268326 5674 268332 5676
rect 267917 5672 268332 5674
rect 267917 5616 267922 5672
rect 267978 5616 268332 5672
rect 267917 5614 268332 5616
rect 267733 5611 267799 5612
rect 267917 5611 267983 5614
rect 268326 5612 268332 5614
rect 268396 5612 268402 5676
rect 269246 5612 269252 5676
rect 269316 5674 269322 5676
rect 269389 5674 269455 5677
rect 269316 5672 269455 5674
rect 269316 5616 269394 5672
rect 269450 5616 269455 5672
rect 269316 5614 269455 5616
rect 269316 5612 269322 5614
rect 269389 5611 269455 5614
rect 269573 5674 269639 5677
rect 270493 5676 270559 5677
rect 269798 5674 269804 5676
rect 269573 5672 269804 5674
rect 269573 5616 269578 5672
rect 269634 5616 269804 5672
rect 269573 5614 269804 5616
rect 269573 5611 269639 5614
rect 269798 5612 269804 5614
rect 269868 5612 269874 5676
rect 270493 5674 270540 5676
rect 270448 5672 270540 5674
rect 270448 5616 270498 5672
rect 270448 5614 270540 5616
rect 270493 5612 270540 5614
rect 270604 5612 270610 5676
rect 271278 5674 271338 5886
rect 271462 5810 271522 6022
rect 271781 6080 272504 6082
rect 271781 6024 271786 6080
rect 271842 6024 272504 6080
rect 271781 6022 272504 6024
rect 271781 6019 271847 6022
rect 271689 5946 271755 5949
rect 271689 5944 272504 5946
rect 271689 5888 271694 5944
rect 271750 5888 272504 5944
rect 271689 5886 272504 5888
rect 271689 5883 271755 5886
rect 271462 5750 272504 5810
rect 271278 5614 272504 5674
rect 270493 5611 270559 5612
rect 253890 5478 262322 5538
rect 267181 5538 267247 5541
rect 268929 5538 268995 5541
rect 267181 5536 268995 5538
rect 267181 5480 267186 5536
rect 267242 5480 268934 5536
rect 268990 5480 268995 5536
rect 267181 5478 268995 5480
rect 68542 5472 68858 5473
rect 68542 5408 68548 5472
rect 68612 5408 68628 5472
rect 68692 5408 68708 5472
rect 68772 5408 68788 5472
rect 68852 5408 68858 5472
rect 68542 5407 68858 5408
rect 136139 5472 136455 5473
rect 136139 5408 136145 5472
rect 136209 5408 136225 5472
rect 136289 5408 136305 5472
rect 136369 5408 136385 5472
rect 136449 5408 136455 5472
rect 136139 5407 136455 5408
rect 203736 5472 204052 5473
rect 203736 5408 203742 5472
rect 203806 5408 203822 5472
rect 203886 5408 203902 5472
rect 203966 5408 203982 5472
rect 204046 5408 204052 5472
rect 203736 5407 204052 5408
rect 42057 5402 42123 5405
rect 47945 5402 48011 5405
rect 42057 5400 48011 5402
rect 42057 5344 42062 5400
rect 42118 5344 47950 5400
rect 48006 5344 48011 5400
rect 42057 5342 48011 5344
rect 42057 5339 42123 5342
rect 47945 5339 48011 5342
rect 91461 5402 91527 5405
rect 109401 5402 109467 5405
rect 91461 5400 109467 5402
rect 91461 5344 91466 5400
rect 91522 5344 109406 5400
rect 109462 5344 109467 5400
rect 91461 5342 109467 5344
rect 91461 5339 91527 5342
rect 109401 5339 109467 5342
rect 146293 5402 146359 5405
rect 177573 5402 177639 5405
rect 146293 5400 177639 5402
rect 146293 5344 146298 5400
rect 146354 5344 177578 5400
rect 177634 5344 177639 5400
rect 146293 5342 177639 5344
rect 146293 5339 146359 5342
rect 177573 5339 177639 5342
rect 219249 5402 219315 5405
rect 230289 5402 230355 5405
rect 219249 5400 230355 5402
rect 219249 5344 219254 5400
rect 219310 5344 230294 5400
rect 230350 5344 230355 5400
rect 219249 5342 230355 5344
rect 219249 5339 219315 5342
rect 230289 5339 230355 5342
rect 230565 5402 230631 5405
rect 253890 5402 253950 5478
rect 267181 5475 267247 5478
rect 268929 5475 268995 5478
rect 271781 5538 271847 5541
rect 271781 5536 272504 5538
rect 271781 5480 271786 5536
rect 271842 5480 272504 5536
rect 271781 5478 272504 5480
rect 271781 5475 271847 5478
rect 271333 5472 271649 5473
rect 271333 5408 271339 5472
rect 271403 5408 271419 5472
rect 271483 5408 271499 5472
rect 271563 5408 271579 5472
rect 271643 5408 271649 5472
rect 271333 5407 271649 5408
rect 230565 5400 253950 5402
rect 230565 5344 230570 5400
rect 230626 5344 253950 5400
rect 230565 5342 253950 5344
rect 264053 5402 264119 5405
rect 267273 5402 267339 5405
rect 264053 5400 267339 5402
rect 264053 5344 264058 5400
rect 264114 5344 267278 5400
rect 267334 5344 267339 5400
rect 264053 5342 267339 5344
rect 230565 5339 230631 5342
rect 264053 5339 264119 5342
rect 267273 5339 267339 5342
rect 268837 5402 268903 5405
rect 271137 5402 271203 5405
rect 268837 5400 271203 5402
rect 268837 5344 268842 5400
rect 268898 5344 271142 5400
rect 271198 5344 271203 5400
rect 268837 5342 271203 5344
rect 268837 5339 268903 5342
rect 271137 5339 271203 5342
rect 271965 5402 272031 5405
rect 271965 5400 272504 5402
rect 271965 5344 271970 5400
rect 272026 5344 272504 5400
rect 271965 5342 272504 5344
rect 271965 5339 272031 5342
rect 67541 5266 67607 5269
rect 80329 5266 80395 5269
rect 67541 5264 80395 5266
rect 67541 5208 67546 5264
rect 67602 5208 80334 5264
rect 80390 5208 80395 5264
rect 67541 5206 80395 5208
rect 67541 5203 67607 5206
rect 80329 5203 80395 5206
rect 80881 5266 80947 5269
rect 108389 5266 108455 5269
rect 122189 5266 122255 5269
rect 80881 5264 122255 5266
rect 80881 5208 80886 5264
rect 80942 5208 108394 5264
rect 108450 5208 122194 5264
rect 122250 5208 122255 5264
rect 80881 5206 122255 5208
rect 80881 5203 80947 5206
rect 108389 5203 108455 5206
rect 122189 5203 122255 5206
rect 150525 5266 150591 5269
rect 151353 5266 151419 5269
rect 158621 5266 158687 5269
rect 150525 5264 158687 5266
rect 150525 5208 150530 5264
rect 150586 5208 151358 5264
rect 151414 5208 158626 5264
rect 158682 5208 158687 5264
rect 150525 5206 158687 5208
rect 150525 5203 150591 5206
rect 151353 5203 151419 5206
rect 158621 5203 158687 5206
rect 160553 5266 160619 5269
rect 222285 5266 222351 5269
rect 160553 5264 222351 5266
rect 160553 5208 160558 5264
rect 160614 5208 222290 5264
rect 222346 5208 222351 5264
rect 160553 5206 222351 5208
rect 160553 5203 160619 5206
rect 222285 5203 222351 5206
rect 228265 5266 228331 5269
rect 240317 5266 240383 5269
rect 228265 5264 240383 5266
rect 228265 5208 228270 5264
rect 228326 5208 240322 5264
rect 240378 5208 240383 5264
rect 228265 5206 240383 5208
rect 228265 5203 228331 5206
rect 240317 5203 240383 5206
rect 240501 5266 240567 5269
rect 260649 5266 260715 5269
rect 263225 5268 263291 5269
rect 240501 5264 260715 5266
rect 240501 5208 240506 5264
rect 240562 5208 260654 5264
rect 260710 5208 260715 5264
rect 240501 5206 260715 5208
rect 240501 5203 240567 5206
rect 260649 5203 260715 5206
rect 263174 5204 263180 5268
rect 263244 5266 263291 5268
rect 268929 5266 268995 5269
rect 263244 5264 263336 5266
rect 263286 5208 263336 5264
rect 263244 5206 263336 5208
rect 268929 5264 272504 5266
rect 268929 5208 268934 5264
rect 268990 5208 272504 5264
rect 268929 5206 272504 5208
rect 263244 5204 263291 5206
rect 263225 5203 263291 5204
rect 268929 5203 268995 5206
rect 20713 5130 20779 5133
rect 42425 5130 42491 5133
rect 44265 5130 44331 5133
rect 20713 5128 44331 5130
rect 20713 5072 20718 5128
rect 20774 5072 42430 5128
rect 42486 5072 44270 5128
rect 44326 5072 44331 5128
rect 20713 5070 44331 5072
rect 20713 5067 20779 5070
rect 42425 5067 42491 5070
rect 44265 5067 44331 5070
rect 44633 5130 44699 5133
rect 91737 5130 91803 5133
rect 44633 5128 91803 5130
rect 44633 5072 44638 5128
rect 44694 5072 91742 5128
rect 91798 5072 91803 5128
rect 44633 5070 91803 5072
rect 44633 5067 44699 5070
rect 91737 5067 91803 5070
rect 100569 5130 100635 5133
rect 162117 5130 162183 5133
rect 100569 5128 162183 5130
rect 100569 5072 100574 5128
rect 100630 5072 162122 5128
rect 162178 5072 162183 5128
rect 100569 5070 162183 5072
rect 100569 5067 100635 5070
rect 162117 5067 162183 5070
rect 163129 5130 163195 5133
rect 220537 5130 220603 5133
rect 163129 5128 220603 5130
rect 163129 5072 163134 5128
rect 163190 5072 220542 5128
rect 220598 5072 220603 5128
rect 163129 5070 220603 5072
rect 163129 5067 163195 5070
rect 220537 5067 220603 5070
rect 230606 5068 230612 5132
rect 230676 5130 230682 5132
rect 258165 5130 258231 5133
rect 230676 5128 258231 5130
rect 230676 5072 258170 5128
rect 258226 5072 258231 5128
rect 230676 5070 258231 5072
rect 230676 5068 230682 5070
rect 258165 5067 258231 5070
rect 268377 5130 268443 5133
rect 271781 5130 271847 5133
rect 268377 5128 271847 5130
rect 268377 5072 268382 5128
rect 268438 5072 271786 5128
rect 271842 5072 271847 5128
rect 268377 5070 271847 5072
rect 268377 5067 268443 5070
rect 271781 5067 271847 5070
rect 271965 5130 272031 5133
rect 271965 5128 272504 5130
rect 271965 5072 271970 5128
rect 272026 5072 272504 5128
rect 271965 5070 272504 5072
rect 271965 5067 272031 5070
rect 42517 4994 42583 4997
rect 43805 4994 43871 4997
rect 42517 4992 43871 4994
rect 42517 4936 42522 4992
rect 42578 4936 43810 4992
rect 43866 4936 43871 4992
rect 42517 4934 43871 4936
rect 42517 4931 42583 4934
rect 43805 4931 43871 4934
rect 204253 4994 204319 4997
rect 229737 4994 229803 4997
rect 204253 4992 229803 4994
rect 204253 4936 204258 4992
rect 204314 4936 229742 4992
rect 229798 4936 229803 4992
rect 204253 4934 229803 4936
rect 204253 4931 204319 4934
rect 229737 4931 229803 4934
rect 268101 4994 268167 4997
rect 268101 4992 272504 4994
rect 268101 4936 268106 4992
rect 268162 4936 272504 4992
rect 268101 4934 272504 4936
rect 268101 4931 268167 4934
rect 34744 4928 35060 4929
rect 34744 4864 34750 4928
rect 34814 4864 34830 4928
rect 34894 4864 34910 4928
rect 34974 4864 34990 4928
rect 35054 4864 35060 4928
rect 34744 4863 35060 4864
rect 102341 4928 102657 4929
rect 102341 4864 102347 4928
rect 102411 4864 102427 4928
rect 102491 4864 102507 4928
rect 102571 4864 102587 4928
rect 102651 4864 102657 4928
rect 102341 4863 102657 4864
rect 169938 4928 170254 4929
rect 169938 4864 169944 4928
rect 170008 4864 170024 4928
rect 170088 4864 170104 4928
rect 170168 4864 170184 4928
rect 170248 4864 170254 4928
rect 169938 4863 170254 4864
rect 237535 4928 237851 4929
rect 237535 4864 237541 4928
rect 237605 4864 237621 4928
rect 237685 4864 237701 4928
rect 237765 4864 237781 4928
rect 237845 4864 237851 4928
rect 237535 4863 237851 4864
rect 214557 4858 214623 4861
rect 219709 4858 219775 4861
rect 214557 4856 219775 4858
rect 214557 4800 214562 4856
rect 214618 4800 219714 4856
rect 219770 4800 219775 4856
rect 214557 4798 219775 4800
rect 214557 4795 214623 4798
rect 219709 4795 219775 4798
rect 224861 4858 224927 4861
rect 227713 4858 227779 4861
rect 224861 4856 227779 4858
rect 224861 4800 224866 4856
rect 224922 4800 227718 4856
rect 227774 4800 227779 4856
rect 224861 4798 227779 4800
rect 224861 4795 224927 4798
rect 227713 4795 227779 4798
rect 228173 4858 228239 4861
rect 237281 4858 237347 4861
rect 228173 4856 237347 4858
rect 228173 4800 228178 4856
rect 228234 4800 237286 4856
rect 237342 4800 237347 4856
rect 228173 4798 237347 4800
rect 228173 4795 228239 4798
rect 237281 4795 237347 4798
rect 268837 4858 268903 4861
rect 268837 4856 272504 4858
rect 268837 4800 268842 4856
rect 268898 4800 272504 4856
rect 268837 4798 272504 4800
rect 268837 4795 268903 4798
rect 81433 4722 81499 4725
rect 94405 4722 94471 4725
rect 182541 4722 182607 4725
rect 81433 4720 182607 4722
rect 81433 4664 81438 4720
rect 81494 4664 94410 4720
rect 94466 4664 182546 4720
rect 182602 4664 182607 4720
rect 81433 4662 182607 4664
rect 81433 4659 81499 4662
rect 94405 4659 94471 4662
rect 182541 4659 182607 4662
rect 216213 4722 216279 4725
rect 217409 4722 217475 4725
rect 216213 4720 217475 4722
rect 216213 4664 216218 4720
rect 216274 4664 217414 4720
rect 217470 4664 217475 4720
rect 216213 4662 217475 4664
rect 216213 4659 216279 4662
rect 217409 4659 217475 4662
rect 217685 4722 217751 4725
rect 250621 4722 250687 4725
rect 217685 4720 250687 4722
rect 217685 4664 217690 4720
rect 217746 4664 250626 4720
rect 250682 4664 250687 4720
rect 217685 4662 250687 4664
rect 217685 4659 217751 4662
rect 250621 4659 250687 4662
rect 267733 4722 267799 4725
rect 272149 4722 272215 4725
rect 267733 4720 272028 4722
rect 267733 4664 267738 4720
rect 267794 4664 272028 4720
rect 267733 4662 272028 4664
rect 267733 4659 267799 4662
rect 42241 4586 42307 4589
rect 94313 4586 94379 4589
rect 42241 4584 94379 4586
rect 42241 4528 42246 4584
rect 42302 4528 94318 4584
rect 94374 4528 94379 4584
rect 42241 4526 94379 4528
rect 42241 4523 42307 4526
rect 94313 4523 94379 4526
rect 116209 4586 116275 4589
rect 151997 4586 152063 4589
rect 116209 4584 152063 4586
rect 116209 4528 116214 4584
rect 116270 4528 152002 4584
rect 152058 4528 152063 4584
rect 116209 4526 152063 4528
rect 116209 4523 116275 4526
rect 151997 4523 152063 4526
rect 160829 4586 160895 4589
rect 223389 4586 223455 4589
rect 226241 4586 226307 4589
rect 228725 4586 228791 4589
rect 242249 4586 242315 4589
rect 160829 4584 223455 4586
rect 160829 4528 160834 4584
rect 160890 4528 223394 4584
rect 223450 4528 223455 4584
rect 160829 4526 223455 4528
rect 160829 4523 160895 4526
rect 223389 4523 223455 4526
rect 226198 4584 242315 4586
rect 226198 4528 226246 4584
rect 226302 4528 228730 4584
rect 228786 4528 242254 4584
rect 242310 4528 242315 4584
rect 226198 4526 242315 4528
rect 226198 4523 226307 4526
rect 228725 4523 228791 4526
rect 242249 4523 242315 4526
rect 264881 4586 264947 4589
rect 264881 4584 271890 4586
rect 264881 4528 264886 4584
rect 264942 4528 271890 4584
rect 264881 4526 271890 4528
rect 264881 4523 264947 4526
rect 19333 4450 19399 4453
rect 46933 4450 46999 4453
rect 48129 4450 48195 4453
rect 19333 4448 48195 4450
rect 19333 4392 19338 4448
rect 19394 4392 46938 4448
rect 46994 4392 48134 4448
rect 48190 4392 48195 4448
rect 19333 4390 48195 4392
rect 19333 4387 19399 4390
rect 46933 4387 46999 4390
rect 48129 4387 48195 4390
rect 92473 4450 92539 4453
rect 113357 4450 113423 4453
rect 92473 4448 113423 4450
rect 92473 4392 92478 4448
rect 92534 4392 113362 4448
rect 113418 4392 113423 4448
rect 92473 4390 113423 4392
rect 92473 4387 92539 4390
rect 113357 4387 113423 4390
rect 151629 4450 151695 4453
rect 173801 4450 173867 4453
rect 226198 4450 226258 4523
rect 151629 4448 173867 4450
rect 151629 4392 151634 4448
rect 151690 4392 173806 4448
rect 173862 4392 173867 4448
rect 151629 4390 173867 4392
rect 151629 4387 151695 4390
rect 173801 4387 173867 4390
rect 209730 4390 226258 4450
rect 267273 4450 267339 4453
rect 271137 4450 271203 4453
rect 267273 4448 271203 4450
rect 267273 4392 267278 4448
rect 267334 4392 271142 4448
rect 271198 4392 271203 4448
rect 267273 4390 271203 4392
rect 68542 4384 68858 4385
rect 68542 4320 68548 4384
rect 68612 4320 68628 4384
rect 68692 4320 68708 4384
rect 68772 4320 68788 4384
rect 68852 4320 68858 4384
rect 68542 4319 68858 4320
rect 136139 4384 136455 4385
rect 136139 4320 136145 4384
rect 136209 4320 136225 4384
rect 136289 4320 136305 4384
rect 136369 4320 136385 4384
rect 136449 4320 136455 4384
rect 136139 4319 136455 4320
rect 203736 4384 204052 4385
rect 203736 4320 203742 4384
rect 203806 4320 203822 4384
rect 203886 4320 203902 4384
rect 203966 4320 203982 4384
rect 204046 4320 204052 4384
rect 203736 4319 204052 4320
rect 40953 4314 41019 4317
rect 41413 4314 41479 4317
rect 40953 4312 41479 4314
rect 40953 4256 40958 4312
rect 41014 4256 41418 4312
rect 41474 4256 41479 4312
rect 40953 4254 41479 4256
rect 40953 4251 41019 4254
rect 41413 4251 41479 4254
rect 44265 4314 44331 4317
rect 60733 4314 60799 4317
rect 44265 4312 60799 4314
rect 44265 4256 44270 4312
rect 44326 4256 60738 4312
rect 60794 4256 60799 4312
rect 44265 4254 60799 4256
rect 44265 4251 44331 4254
rect 60733 4251 60799 4254
rect 98085 4314 98151 4317
rect 99465 4314 99531 4317
rect 100845 4314 100911 4317
rect 101397 4314 101463 4317
rect 98085 4312 101463 4314
rect 98085 4256 98090 4312
rect 98146 4256 99470 4312
rect 99526 4256 100850 4312
rect 100906 4256 101402 4312
rect 101458 4256 101463 4312
rect 98085 4254 101463 4256
rect 98085 4251 98151 4254
rect 99465 4251 99531 4254
rect 100845 4251 100911 4254
rect 101397 4251 101463 4254
rect 175917 4178 175983 4181
rect 209730 4178 209790 4390
rect 267273 4387 267339 4390
rect 271137 4387 271203 4390
rect 271333 4384 271649 4385
rect 271333 4320 271339 4384
rect 271403 4320 271419 4384
rect 271483 4320 271499 4384
rect 271563 4320 271579 4384
rect 271643 4320 271649 4384
rect 271333 4319 271649 4320
rect 224677 4314 224743 4317
rect 242893 4314 242959 4317
rect 224677 4312 242959 4314
rect 224677 4256 224682 4312
rect 224738 4256 242898 4312
rect 242954 4256 242959 4312
rect 224677 4254 242959 4256
rect 224677 4251 224743 4254
rect 242893 4251 242959 4254
rect 255037 4314 255103 4317
rect 260189 4314 260255 4317
rect 255037 4312 260255 4314
rect 255037 4256 255042 4312
rect 255098 4256 260194 4312
rect 260250 4256 260255 4312
rect 255037 4254 260255 4256
rect 255037 4251 255103 4254
rect 260189 4251 260255 4254
rect 266445 4314 266511 4317
rect 268561 4314 268627 4317
rect 266445 4312 268627 4314
rect 266445 4256 266450 4312
rect 266506 4256 268566 4312
rect 268622 4256 268627 4312
rect 266445 4254 268627 4256
rect 271830 4314 271890 4526
rect 271968 4450 272028 4662
rect 272149 4720 272504 4722
rect 272149 4664 272154 4720
rect 272210 4664 272504 4720
rect 272149 4662 272504 4664
rect 272149 4659 272215 4662
rect 272304 4526 272504 4586
rect 271968 4390 272504 4450
rect 271830 4254 272504 4314
rect 266445 4251 266511 4254
rect 268561 4251 268627 4254
rect 175917 4176 209790 4178
rect 175917 4120 175922 4176
rect 175978 4120 209790 4176
rect 175917 4118 209790 4120
rect 213637 4178 213703 4181
rect 214005 4178 214071 4181
rect 216029 4178 216095 4181
rect 213637 4176 216095 4178
rect 213637 4120 213642 4176
rect 213698 4120 214010 4176
rect 214066 4120 216034 4176
rect 216090 4120 216095 4176
rect 213637 4118 216095 4120
rect 175917 4115 175983 4118
rect 213637 4115 213703 4118
rect 214005 4115 214071 4118
rect 216029 4115 216095 4118
rect 223205 4178 223271 4181
rect 225873 4178 225939 4181
rect 223205 4176 225939 4178
rect 223205 4120 223210 4176
rect 223266 4120 225878 4176
rect 225934 4120 225939 4176
rect 223205 4118 225939 4120
rect 223205 4115 223271 4118
rect 225873 4115 225939 4118
rect 226701 4178 226767 4181
rect 230749 4178 230815 4181
rect 226701 4176 230815 4178
rect 226701 4120 226706 4176
rect 226762 4120 230754 4176
rect 230810 4120 230815 4176
rect 226701 4118 230815 4120
rect 226701 4115 226767 4118
rect 230749 4115 230815 4118
rect 244181 4178 244247 4181
rect 244181 4176 272504 4178
rect 244181 4120 244186 4176
rect 244242 4120 272504 4176
rect 244181 4118 272504 4120
rect 244181 4115 244247 4118
rect 49785 4042 49851 4045
rect 51625 4042 51691 4045
rect 49785 4040 51691 4042
rect 49785 3984 49790 4040
rect 49846 3984 51630 4040
rect 51686 3984 51691 4040
rect 49785 3982 51691 3984
rect 49785 3979 49851 3982
rect 51625 3979 51691 3982
rect 96153 4042 96219 4045
rect 110505 4042 110571 4045
rect 96153 4040 110571 4042
rect 96153 3984 96158 4040
rect 96214 3984 110510 4040
rect 110566 3984 110571 4040
rect 96153 3982 110571 3984
rect 96153 3979 96219 3982
rect 110505 3979 110571 3982
rect 149789 4042 149855 4045
rect 212349 4042 212415 4045
rect 149789 4040 212415 4042
rect 149789 3984 149794 4040
rect 149850 3984 212354 4040
rect 212410 3984 212415 4040
rect 149789 3982 212415 3984
rect 149789 3979 149855 3982
rect 212349 3979 212415 3982
rect 216489 4042 216555 4045
rect 238201 4042 238267 4045
rect 216489 4040 238267 4042
rect 216489 3984 216494 4040
rect 216550 3984 238206 4040
rect 238262 3984 238267 4040
rect 216489 3982 238267 3984
rect 216489 3979 216555 3982
rect 238201 3979 238267 3982
rect 240777 4042 240843 4045
rect 268009 4042 268075 4045
rect 240777 4040 268075 4042
rect 240777 3984 240782 4040
rect 240838 3984 268014 4040
rect 268070 3984 268075 4040
rect 240777 3982 268075 3984
rect 240777 3979 240843 3982
rect 268009 3979 268075 3982
rect 268469 4042 268535 4045
rect 271137 4042 271203 4045
rect 268469 4040 271203 4042
rect 268469 3984 268474 4040
rect 268530 3984 271142 4040
rect 271198 3984 271203 4040
rect 268469 3982 271203 3984
rect 268469 3979 268535 3982
rect 271137 3979 271203 3982
rect 271278 3982 272504 4042
rect 119981 3906 120047 3909
rect 159909 3906 159975 3909
rect 119981 3904 159975 3906
rect 119981 3848 119986 3904
rect 120042 3848 159914 3904
rect 159970 3848 159975 3904
rect 119981 3846 159975 3848
rect 119981 3843 120047 3846
rect 159909 3843 159975 3846
rect 216121 3906 216187 3909
rect 217501 3906 217567 3909
rect 216121 3904 217567 3906
rect 216121 3848 216126 3904
rect 216182 3848 217506 3904
rect 217562 3848 217567 3904
rect 216121 3846 217567 3848
rect 216121 3843 216187 3846
rect 217501 3843 217567 3846
rect 227437 3906 227503 3909
rect 229093 3906 229159 3909
rect 227437 3904 229159 3906
rect 227437 3848 227442 3904
rect 227498 3848 229098 3904
rect 229154 3848 229159 3904
rect 227437 3846 229159 3848
rect 227437 3843 227503 3846
rect 229093 3843 229159 3846
rect 242525 3906 242591 3909
rect 271278 3906 271338 3982
rect 242525 3904 271338 3906
rect 242525 3848 242530 3904
rect 242586 3848 271338 3904
rect 242525 3846 271338 3848
rect 271462 3846 272504 3906
rect 242525 3843 242591 3846
rect 34744 3840 35060 3841
rect 34744 3776 34750 3840
rect 34814 3776 34830 3840
rect 34894 3776 34910 3840
rect 34974 3776 34990 3840
rect 35054 3776 35060 3840
rect 34744 3775 35060 3776
rect 102341 3840 102657 3841
rect 102341 3776 102347 3840
rect 102411 3776 102427 3840
rect 102491 3776 102507 3840
rect 102571 3776 102587 3840
rect 102651 3776 102657 3840
rect 102341 3775 102657 3776
rect 169938 3840 170254 3841
rect 169938 3776 169944 3840
rect 170008 3776 170024 3840
rect 170088 3776 170104 3840
rect 170168 3776 170184 3840
rect 170248 3776 170254 3840
rect 169938 3775 170254 3776
rect 237535 3840 237851 3841
rect 237535 3776 237541 3840
rect 237605 3776 237621 3840
rect 237685 3776 237701 3840
rect 237765 3776 237781 3840
rect 237845 3776 237851 3840
rect 237535 3775 237851 3776
rect 207197 3770 207263 3773
rect 214465 3770 214531 3773
rect 207197 3768 214531 3770
rect 207197 3712 207202 3768
rect 207258 3712 214470 3768
rect 214526 3712 214531 3768
rect 207197 3710 214531 3712
rect 207197 3707 207263 3710
rect 214465 3707 214531 3710
rect 215334 3708 215340 3772
rect 215404 3770 215410 3772
rect 216581 3770 216647 3773
rect 215404 3768 216647 3770
rect 215404 3712 216586 3768
rect 216642 3712 216647 3768
rect 215404 3710 216647 3712
rect 215404 3708 215410 3710
rect 216581 3707 216647 3710
rect 218789 3770 218855 3773
rect 227897 3770 227963 3773
rect 218789 3768 227963 3770
rect 218789 3712 218794 3768
rect 218850 3712 227902 3768
rect 227958 3712 227963 3768
rect 218789 3710 227963 3712
rect 218789 3707 218855 3710
rect 227897 3707 227963 3710
rect 237925 3770 237991 3773
rect 243721 3770 243787 3773
rect 237925 3768 243787 3770
rect 237925 3712 237930 3768
rect 237986 3712 243726 3768
rect 243782 3712 243787 3768
rect 237925 3710 243787 3712
rect 237925 3707 237991 3710
rect 243721 3707 243787 3710
rect 267365 3770 267431 3773
rect 267590 3770 267596 3772
rect 267365 3768 267596 3770
rect 267365 3712 267370 3768
rect 267426 3712 267596 3768
rect 267365 3710 267596 3712
rect 267365 3707 267431 3710
rect 267590 3708 267596 3710
rect 267660 3708 267666 3772
rect 268009 3770 268075 3773
rect 271462 3770 271522 3846
rect 268009 3768 271522 3770
rect 268009 3712 268014 3768
rect 268070 3712 271522 3768
rect 268009 3710 271522 3712
rect 271597 3770 271663 3773
rect 271597 3768 272504 3770
rect 271597 3712 271602 3768
rect 271658 3712 272504 3768
rect 271597 3710 272504 3712
rect 268009 3707 268075 3710
rect 271597 3707 271663 3710
rect 85665 3634 85731 3637
rect 96613 3634 96679 3637
rect 85665 3632 96679 3634
rect 85665 3576 85670 3632
rect 85726 3576 96618 3632
rect 96674 3576 96679 3632
rect 85665 3574 96679 3576
rect 85665 3571 85731 3574
rect 96613 3571 96679 3574
rect 116117 3634 116183 3637
rect 120349 3634 120415 3637
rect 116117 3632 120415 3634
rect 116117 3576 116122 3632
rect 116178 3576 120354 3632
rect 120410 3576 120415 3632
rect 116117 3574 120415 3576
rect 116117 3571 116183 3574
rect 120349 3571 120415 3574
rect 144269 3634 144335 3637
rect 144729 3634 144795 3637
rect 144269 3632 144795 3634
rect 144269 3576 144274 3632
rect 144330 3576 144734 3632
rect 144790 3576 144795 3632
rect 144269 3574 144795 3576
rect 144269 3571 144335 3574
rect 144729 3571 144795 3574
rect 156689 3634 156755 3637
rect 161657 3634 161723 3637
rect 156689 3632 161723 3634
rect 156689 3576 156694 3632
rect 156750 3576 161662 3632
rect 161718 3576 161723 3632
rect 156689 3574 161723 3576
rect 156689 3571 156755 3574
rect 161657 3571 161723 3574
rect 208669 3634 208735 3637
rect 238109 3634 238175 3637
rect 208669 3632 238175 3634
rect 208669 3576 208674 3632
rect 208730 3576 238114 3632
rect 238170 3576 238175 3632
rect 208669 3574 238175 3576
rect 208669 3571 208735 3574
rect 238109 3571 238175 3574
rect 265433 3634 265499 3637
rect 267733 3634 267799 3637
rect 265433 3632 267799 3634
rect 265433 3576 265438 3632
rect 265494 3576 267738 3632
rect 267794 3576 267799 3632
rect 265433 3574 267799 3576
rect 265433 3571 265499 3574
rect 267733 3571 267799 3574
rect 267917 3634 267983 3637
rect 267917 3632 272504 3634
rect 267917 3576 267922 3632
rect 267978 3576 272504 3632
rect 267917 3574 272504 3576
rect 267917 3571 267983 3574
rect 39113 3498 39179 3501
rect 86585 3498 86651 3501
rect 39113 3496 86651 3498
rect 39113 3440 39118 3496
rect 39174 3440 86590 3496
rect 86646 3440 86651 3496
rect 39113 3438 86651 3440
rect 39113 3435 39179 3438
rect 86585 3435 86651 3438
rect 95877 3498 95943 3501
rect 109033 3498 109099 3501
rect 150065 3498 150131 3501
rect 214097 3498 214163 3501
rect 95877 3496 214163 3498
rect 95877 3440 95882 3496
rect 95938 3440 109038 3496
rect 109094 3440 150070 3496
rect 150126 3440 214102 3496
rect 214158 3440 214163 3496
rect 95877 3438 214163 3440
rect 95877 3435 95943 3438
rect 109033 3435 109099 3438
rect 150065 3435 150131 3438
rect 214097 3435 214163 3438
rect 228357 3498 228423 3501
rect 259269 3498 259335 3501
rect 228357 3496 259335 3498
rect 228357 3440 228362 3496
rect 228418 3440 259274 3496
rect 259330 3440 259335 3496
rect 228357 3438 259335 3440
rect 228357 3435 228423 3438
rect 259269 3435 259335 3438
rect 260833 3498 260899 3501
rect 271965 3498 272031 3501
rect 260833 3496 271890 3498
rect 260833 3440 260838 3496
rect 260894 3440 271890 3496
rect 260833 3438 271890 3440
rect 260833 3435 260899 3438
rect 24342 3300 24348 3364
rect 24412 3362 24418 3364
rect 24485 3362 24551 3365
rect 24412 3360 24551 3362
rect 24412 3304 24490 3360
rect 24546 3304 24551 3360
rect 24412 3302 24551 3304
rect 24412 3300 24418 3302
rect 24485 3299 24551 3302
rect 85665 3362 85731 3365
rect 120625 3362 120691 3365
rect 85665 3360 120691 3362
rect 85665 3304 85670 3360
rect 85726 3304 120630 3360
rect 120686 3304 120691 3360
rect 85665 3302 120691 3304
rect 85665 3299 85731 3302
rect 120625 3299 120691 3302
rect 155033 3362 155099 3365
rect 174169 3362 174235 3365
rect 155033 3360 174235 3362
rect 155033 3304 155038 3360
rect 155094 3304 174174 3360
rect 174230 3304 174235 3360
rect 155033 3302 174235 3304
rect 155033 3299 155099 3302
rect 174169 3299 174235 3302
rect 213545 3362 213611 3365
rect 237833 3362 237899 3365
rect 241513 3362 241579 3365
rect 213545 3360 237899 3362
rect 213545 3304 213550 3360
rect 213606 3304 237838 3360
rect 237894 3304 237899 3360
rect 213545 3302 237899 3304
rect 213545 3299 213611 3302
rect 237833 3299 237899 3302
rect 237974 3360 241579 3362
rect 237974 3304 241518 3360
rect 241574 3304 241579 3360
rect 237974 3302 241579 3304
rect 68542 3296 68858 3297
rect 68542 3232 68548 3296
rect 68612 3232 68628 3296
rect 68692 3232 68708 3296
rect 68772 3232 68788 3296
rect 68852 3232 68858 3296
rect 68542 3231 68858 3232
rect 136139 3296 136455 3297
rect 136139 3232 136145 3296
rect 136209 3232 136225 3296
rect 136289 3232 136305 3296
rect 136369 3232 136385 3296
rect 136449 3232 136455 3296
rect 136139 3231 136455 3232
rect 203736 3296 204052 3297
rect 203736 3232 203742 3296
rect 203806 3232 203822 3296
rect 203886 3232 203902 3296
rect 203966 3232 203982 3296
rect 204046 3232 204052 3296
rect 203736 3231 204052 3232
rect 82169 3226 82235 3229
rect 101673 3226 101739 3229
rect 82169 3224 101739 3226
rect 82169 3168 82174 3224
rect 82230 3168 101678 3224
rect 101734 3168 101739 3224
rect 82169 3166 101739 3168
rect 82169 3163 82235 3166
rect 101673 3163 101739 3166
rect 156045 3226 156111 3229
rect 156597 3226 156663 3229
rect 157057 3226 157123 3229
rect 156045 3224 157123 3226
rect 156045 3168 156050 3224
rect 156106 3168 156602 3224
rect 156658 3168 157062 3224
rect 157118 3168 157123 3224
rect 156045 3166 157123 3168
rect 156045 3163 156111 3166
rect 156597 3163 156663 3166
rect 157057 3163 157123 3166
rect 210969 3226 211035 3229
rect 237974 3226 238034 3302
rect 241513 3299 241579 3302
rect 267733 3362 267799 3365
rect 271137 3362 271203 3365
rect 267733 3360 271203 3362
rect 267733 3304 267738 3360
rect 267794 3304 271142 3360
rect 271198 3304 271203 3360
rect 267733 3302 271203 3304
rect 271830 3362 271890 3438
rect 271965 3496 272504 3498
rect 271965 3440 271970 3496
rect 272026 3440 272504 3496
rect 271965 3438 272504 3440
rect 271965 3435 272031 3438
rect 271830 3302 272504 3362
rect 267733 3299 267799 3302
rect 271137 3299 271203 3302
rect 271333 3296 271649 3297
rect 271333 3232 271339 3296
rect 271403 3232 271419 3296
rect 271483 3232 271499 3296
rect 271563 3232 271579 3296
rect 271643 3232 271649 3296
rect 271333 3231 271649 3232
rect 210969 3224 238034 3226
rect 210969 3168 210974 3224
rect 211030 3168 238034 3224
rect 210969 3166 238034 3168
rect 238661 3226 238727 3229
rect 240501 3226 240567 3229
rect 238661 3224 240567 3226
rect 238661 3168 238666 3224
rect 238722 3168 240506 3224
rect 240562 3168 240567 3224
rect 238661 3166 240567 3168
rect 210969 3163 211035 3166
rect 238661 3163 238727 3166
rect 240501 3163 240567 3166
rect 265893 3226 265959 3229
rect 267958 3226 267964 3228
rect 265893 3224 267964 3226
rect 265893 3168 265898 3224
rect 265954 3168 267964 3224
rect 265893 3166 267964 3168
rect 265893 3163 265959 3166
rect 267958 3164 267964 3166
rect 268028 3164 268034 3228
rect 268101 3226 268167 3229
rect 270769 3226 270835 3229
rect 268101 3224 270835 3226
rect 268101 3168 268106 3224
rect 268162 3168 270774 3224
rect 270830 3168 270835 3224
rect 268101 3166 270835 3168
rect 268101 3163 268167 3166
rect 270769 3163 270835 3166
rect 271781 3226 271847 3229
rect 271781 3224 272504 3226
rect 271781 3168 271786 3224
rect 271842 3168 272504 3224
rect 271781 3166 272504 3168
rect 271781 3163 271847 3166
rect 25221 3090 25287 3093
rect 54385 3090 54451 3093
rect 25221 3088 54451 3090
rect 25221 3032 25226 3088
rect 25282 3032 54390 3088
rect 54446 3032 54451 3088
rect 25221 3030 54451 3032
rect 25221 3027 25287 3030
rect 54385 3027 54451 3030
rect 82353 3090 82419 3093
rect 112529 3090 112595 3093
rect 82353 3088 112595 3090
rect 82353 3032 82358 3088
rect 82414 3032 112534 3088
rect 112590 3032 112595 3088
rect 82353 3030 112595 3032
rect 82353 3027 82419 3030
rect 112529 3027 112595 3030
rect 143717 3090 143783 3093
rect 160001 3090 160067 3093
rect 143717 3088 160067 3090
rect 143717 3032 143722 3088
rect 143778 3032 160006 3088
rect 160062 3032 160067 3088
rect 143717 3030 160067 3032
rect 143717 3027 143783 3030
rect 160001 3027 160067 3030
rect 216305 3090 216371 3093
rect 222193 3090 222259 3093
rect 216305 3088 222259 3090
rect 216305 3032 216310 3088
rect 216366 3032 222198 3088
rect 222254 3032 222259 3088
rect 216305 3030 222259 3032
rect 216305 3027 216371 3030
rect 222193 3027 222259 3030
rect 223205 3090 223271 3093
rect 262213 3090 262279 3093
rect 223205 3088 253950 3090
rect 223205 3032 223210 3088
rect 223266 3032 253950 3088
rect 223205 3030 253950 3032
rect 223205 3027 223271 3030
rect 19241 2956 19307 2957
rect 22921 2956 22987 2957
rect 19190 2954 19196 2956
rect 19150 2894 19196 2954
rect 19260 2952 19307 2956
rect 22870 2954 22876 2956
rect 19302 2896 19307 2952
rect 19190 2892 19196 2894
rect 19260 2892 19307 2896
rect 22830 2894 22876 2954
rect 22940 2952 22987 2956
rect 22982 2896 22987 2952
rect 22870 2892 22876 2894
rect 22940 2892 22987 2896
rect 19241 2891 19307 2892
rect 22921 2891 22987 2892
rect 41137 2954 41203 2957
rect 90081 2954 90147 2957
rect 41137 2952 90147 2954
rect 41137 2896 41142 2952
rect 41198 2896 90086 2952
rect 90142 2896 90147 2952
rect 41137 2894 90147 2896
rect 41137 2891 41203 2894
rect 90081 2891 90147 2894
rect 99373 2954 99439 2957
rect 115749 2954 115815 2957
rect 99373 2952 115815 2954
rect 99373 2896 99378 2952
rect 99434 2896 115754 2952
rect 115810 2896 115815 2952
rect 99373 2894 115815 2896
rect 99373 2891 99439 2894
rect 115749 2891 115815 2894
rect 140681 2954 140747 2957
rect 203793 2954 203859 2957
rect 204437 2954 204503 2957
rect 140681 2952 204503 2954
rect 140681 2896 140686 2952
rect 140742 2896 203798 2952
rect 203854 2896 204442 2952
rect 204498 2896 204503 2952
rect 140681 2894 204503 2896
rect 140681 2891 140747 2894
rect 203793 2891 203859 2894
rect 204437 2891 204503 2894
rect 213913 2954 213979 2957
rect 245009 2954 245075 2957
rect 213913 2952 245075 2954
rect 213913 2896 213918 2952
rect 213974 2896 245014 2952
rect 245070 2896 245075 2952
rect 213913 2894 245075 2896
rect 253890 2954 253950 3030
rect 262213 3088 272504 3090
rect 262213 3032 262218 3088
rect 262274 3032 272504 3088
rect 262213 3030 272504 3032
rect 262213 3027 262279 3030
rect 266813 2954 266879 2957
rect 253890 2952 266879 2954
rect 253890 2896 266818 2952
rect 266874 2896 266879 2952
rect 253890 2894 266879 2896
rect 213913 2891 213979 2894
rect 245009 2891 245075 2894
rect 266813 2891 266879 2894
rect 268009 2954 268075 2957
rect 271781 2954 271847 2957
rect 268009 2952 271847 2954
rect 268009 2896 268014 2952
rect 268070 2896 271786 2952
rect 271842 2896 271847 2952
rect 268009 2894 271847 2896
rect 268009 2891 268075 2894
rect 271781 2891 271847 2894
rect 271965 2954 272031 2957
rect 271965 2952 272504 2954
rect 271965 2896 271970 2952
rect 272026 2896 272504 2952
rect 271965 2894 272504 2896
rect 271965 2891 272031 2894
rect 19977 2820 20043 2821
rect 19926 2818 19932 2820
rect 19886 2758 19932 2818
rect 19996 2816 20043 2820
rect 20038 2760 20043 2816
rect 19926 2756 19932 2758
rect 19996 2756 20043 2760
rect 22134 2756 22140 2820
rect 22204 2818 22210 2820
rect 23381 2818 23447 2821
rect 22204 2816 23447 2818
rect 22204 2760 23386 2816
rect 23442 2760 23447 2816
rect 22204 2758 23447 2760
rect 22204 2756 22210 2758
rect 19977 2755 20043 2756
rect 23381 2755 23447 2758
rect 25078 2756 25084 2820
rect 25148 2818 25154 2820
rect 28073 2818 28139 2821
rect 25148 2816 28139 2818
rect 25148 2760 28078 2816
rect 28134 2760 28139 2816
rect 25148 2758 28139 2760
rect 25148 2756 25154 2758
rect 28073 2755 28139 2758
rect 60038 2756 60044 2820
rect 60108 2818 60114 2820
rect 60733 2818 60799 2821
rect 157241 2820 157307 2821
rect 157190 2818 157196 2820
rect 60108 2816 60799 2818
rect 60108 2760 60738 2816
rect 60794 2760 60799 2816
rect 60108 2758 60799 2760
rect 157150 2758 157196 2818
rect 157260 2816 157307 2820
rect 157302 2760 157307 2816
rect 60108 2756 60114 2758
rect 60733 2755 60799 2758
rect 157190 2756 157196 2758
rect 157260 2756 157307 2760
rect 159398 2756 159404 2820
rect 159468 2818 159474 2820
rect 160001 2818 160067 2821
rect 159468 2816 160067 2818
rect 159468 2760 160006 2816
rect 160062 2760 160067 2816
rect 159468 2758 160067 2760
rect 159468 2756 159474 2758
rect 157241 2755 157307 2756
rect 160001 2755 160067 2758
rect 189942 2756 189948 2820
rect 190012 2818 190018 2820
rect 190361 2818 190427 2821
rect 190012 2816 190427 2818
rect 190012 2760 190366 2816
rect 190422 2760 190427 2816
rect 190012 2758 190427 2760
rect 190012 2756 190018 2758
rect 190361 2755 190427 2758
rect 191414 2756 191420 2820
rect 191484 2818 191490 2820
rect 191741 2818 191807 2821
rect 191484 2816 191807 2818
rect 191484 2760 191746 2816
rect 191802 2760 191807 2816
rect 191484 2758 191807 2760
rect 191484 2756 191490 2758
rect 191741 2755 191807 2758
rect 202454 2756 202460 2820
rect 202524 2818 202530 2820
rect 202781 2818 202847 2821
rect 202524 2816 202847 2818
rect 202524 2760 202786 2816
rect 202842 2760 202847 2816
rect 202524 2758 202847 2760
rect 202524 2756 202530 2758
rect 202781 2755 202847 2758
rect 210877 2818 210943 2821
rect 217133 2818 217199 2821
rect 223297 2820 223363 2821
rect 223246 2818 223252 2820
rect 210877 2816 217199 2818
rect 210877 2760 210882 2816
rect 210938 2760 217138 2816
rect 217194 2760 217199 2816
rect 210877 2758 217199 2760
rect 223206 2758 223252 2818
rect 223316 2816 223363 2820
rect 223358 2760 223363 2816
rect 210877 2755 210943 2758
rect 217133 2755 217199 2758
rect 223246 2756 223252 2758
rect 223316 2756 223363 2760
rect 224718 2756 224724 2820
rect 224788 2818 224794 2820
rect 224861 2818 224927 2821
rect 226241 2820 226307 2821
rect 226190 2818 226196 2820
rect 224788 2816 224927 2818
rect 224788 2760 224866 2816
rect 224922 2760 224927 2816
rect 224788 2758 224927 2760
rect 226150 2758 226196 2818
rect 226260 2816 226307 2820
rect 226302 2760 226307 2816
rect 224788 2756 224794 2758
rect 223297 2755 223363 2756
rect 224861 2755 224927 2758
rect 226190 2756 226196 2758
rect 226260 2756 226307 2760
rect 226241 2755 226307 2756
rect 226517 2818 226583 2821
rect 231025 2818 231091 2821
rect 226517 2816 231091 2818
rect 226517 2760 226522 2816
rect 226578 2760 231030 2816
rect 231086 2760 231091 2816
rect 226517 2758 231091 2760
rect 226517 2755 226583 2758
rect 231025 2755 231091 2758
rect 235758 2756 235764 2820
rect 235828 2818 235834 2820
rect 235901 2818 235967 2821
rect 258073 2820 258139 2821
rect 258022 2818 258028 2820
rect 235828 2816 235967 2818
rect 235828 2760 235906 2816
rect 235962 2760 235967 2816
rect 235828 2758 235967 2760
rect 257982 2758 258028 2818
rect 258092 2816 258139 2820
rect 258134 2760 258139 2816
rect 235828 2756 235834 2758
rect 235901 2755 235967 2758
rect 258022 2756 258028 2758
rect 258092 2756 258139 2760
rect 258073 2755 258139 2756
rect 265249 2818 265315 2821
rect 268193 2818 268259 2821
rect 265249 2816 268259 2818
rect 265249 2760 265254 2816
rect 265310 2760 268198 2816
rect 268254 2760 268259 2816
rect 265249 2758 268259 2760
rect 265249 2755 265315 2758
rect 268193 2755 268259 2758
rect 270493 2820 270559 2821
rect 270493 2816 270540 2820
rect 270604 2818 270610 2820
rect 270769 2818 270835 2821
rect 270493 2760 270498 2816
rect 270493 2756 270540 2760
rect 270604 2758 270650 2818
rect 270769 2816 272504 2818
rect 270769 2760 270774 2816
rect 270830 2760 272504 2816
rect 270769 2758 272504 2760
rect 270604 2756 270610 2758
rect 270493 2755 270559 2756
rect 270769 2755 270835 2758
rect 34744 2752 35060 2753
rect 34744 2688 34750 2752
rect 34814 2688 34830 2752
rect 34894 2688 34910 2752
rect 34974 2688 34990 2752
rect 35054 2688 35060 2752
rect 34744 2687 35060 2688
rect 102341 2752 102657 2753
rect 102341 2688 102347 2752
rect 102411 2688 102427 2752
rect 102491 2688 102507 2752
rect 102571 2688 102587 2752
rect 102651 2688 102657 2752
rect 102341 2687 102657 2688
rect 169938 2752 170254 2753
rect 169938 2688 169944 2752
rect 170008 2688 170024 2752
rect 170088 2688 170104 2752
rect 170168 2688 170184 2752
rect 170248 2688 170254 2752
rect 169938 2687 170254 2688
rect 237535 2752 237851 2753
rect 237535 2688 237541 2752
rect 237605 2688 237621 2752
rect 237685 2688 237701 2752
rect 237765 2688 237781 2752
rect 237845 2688 237851 2752
rect 237535 2687 237851 2688
rect 97625 2682 97691 2685
rect 100753 2682 100819 2685
rect 97625 2680 100819 2682
rect 97625 2624 97630 2680
rect 97686 2624 100758 2680
rect 100814 2624 100819 2680
rect 97625 2622 100819 2624
rect 97625 2619 97691 2622
rect 100753 2619 100819 2622
rect 155125 2682 155191 2685
rect 158529 2682 158595 2685
rect 155125 2680 158595 2682
rect 155125 2624 155130 2680
rect 155186 2624 158534 2680
rect 158590 2624 158595 2680
rect 155125 2622 158595 2624
rect 155125 2619 155191 2622
rect 158529 2619 158595 2622
rect 213453 2682 213519 2685
rect 215661 2682 215727 2685
rect 213453 2680 215727 2682
rect 213453 2624 213458 2680
rect 213514 2624 215666 2680
rect 215722 2624 215727 2680
rect 213453 2622 215727 2624
rect 213453 2619 213519 2622
rect 215661 2619 215727 2622
rect 215845 2682 215911 2685
rect 223481 2682 223547 2685
rect 215845 2680 223547 2682
rect 215845 2624 215850 2680
rect 215906 2624 223486 2680
rect 223542 2624 223547 2680
rect 215845 2622 223547 2624
rect 215845 2619 215911 2622
rect 223481 2619 223547 2622
rect 223849 2682 223915 2685
rect 236085 2682 236151 2685
rect 223849 2680 236151 2682
rect 223849 2624 223854 2680
rect 223910 2624 236090 2680
rect 236146 2624 236151 2680
rect 223849 2622 236151 2624
rect 223849 2619 223915 2622
rect 236085 2619 236151 2622
rect 241513 2682 241579 2685
rect 252277 2682 252343 2685
rect 241513 2680 252343 2682
rect 241513 2624 241518 2680
rect 241574 2624 252282 2680
rect 252338 2624 252343 2680
rect 241513 2622 252343 2624
rect 241513 2619 241579 2622
rect 252277 2619 252343 2622
rect 266486 2620 266492 2684
rect 266556 2682 266562 2684
rect 266629 2682 266695 2685
rect 266556 2680 266695 2682
rect 266556 2624 266634 2680
rect 266690 2624 266695 2680
rect 266556 2622 266695 2624
rect 266556 2620 266562 2622
rect 266629 2619 266695 2622
rect 267181 2682 267247 2685
rect 267181 2680 272504 2682
rect 267181 2624 267186 2680
rect 267242 2624 272504 2680
rect 267181 2622 272504 2624
rect 267181 2619 267247 2622
rect 89897 2546 89963 2549
rect 103421 2546 103487 2549
rect 89897 2544 103487 2546
rect 89897 2488 89902 2544
rect 89958 2488 103426 2544
rect 103482 2488 103487 2544
rect 89897 2486 103487 2488
rect 89897 2483 89963 2486
rect 103421 2483 103487 2486
rect 149145 2546 149211 2549
rect 156413 2546 156479 2549
rect 149145 2544 156479 2546
rect 149145 2488 149150 2544
rect 149206 2488 156418 2544
rect 156474 2488 156479 2544
rect 149145 2486 156479 2488
rect 149145 2483 149211 2486
rect 156413 2483 156479 2486
rect 156781 2546 156847 2549
rect 163589 2546 163655 2549
rect 156781 2544 163655 2546
rect 156781 2488 156786 2544
rect 156842 2488 163594 2544
rect 163650 2488 163655 2544
rect 156781 2486 163655 2488
rect 156781 2483 156847 2486
rect 163589 2483 163655 2486
rect 186313 2546 186379 2549
rect 210417 2546 210483 2549
rect 186313 2544 210483 2546
rect 186313 2488 186318 2544
rect 186374 2488 210422 2544
rect 210478 2488 210483 2544
rect 186313 2486 210483 2488
rect 186313 2483 186379 2486
rect 210417 2483 210483 2486
rect 212349 2546 212415 2549
rect 216765 2546 216831 2549
rect 212349 2544 216831 2546
rect 212349 2488 212354 2544
rect 212410 2488 216770 2544
rect 216826 2488 216831 2544
rect 212349 2486 216831 2488
rect 212349 2483 212415 2486
rect 216765 2483 216831 2486
rect 217869 2546 217935 2549
rect 223614 2546 223620 2548
rect 217869 2544 223620 2546
rect 217869 2488 217874 2544
rect 217930 2488 223620 2544
rect 217869 2486 223620 2488
rect 217869 2483 217935 2486
rect 223614 2484 223620 2486
rect 223684 2484 223690 2548
rect 224677 2546 224743 2549
rect 243813 2546 243879 2549
rect 224677 2544 243879 2546
rect 224677 2488 224682 2544
rect 224738 2488 243818 2544
rect 243874 2488 243879 2544
rect 224677 2486 243879 2488
rect 224677 2483 224743 2486
rect 243813 2483 243879 2486
rect 267958 2484 267964 2548
rect 268028 2546 268034 2548
rect 268285 2546 268351 2549
rect 268028 2544 268351 2546
rect 268028 2488 268290 2544
rect 268346 2488 268351 2544
rect 268028 2486 268351 2488
rect 268028 2484 268034 2486
rect 268285 2483 268351 2486
rect 268469 2546 268535 2549
rect 268469 2544 272504 2546
rect 268469 2488 268474 2544
rect 268530 2488 272504 2544
rect 268469 2486 272504 2488
rect 268469 2483 268535 2486
rect 38193 2410 38259 2413
rect 84285 2410 84351 2413
rect 38193 2408 84351 2410
rect 38193 2352 38198 2408
rect 38254 2352 84290 2408
rect 84346 2352 84351 2408
rect 38193 2350 84351 2352
rect 38193 2347 38259 2350
rect 84285 2347 84351 2350
rect 99005 2410 99071 2413
rect 101213 2410 101279 2413
rect 138565 2410 138631 2413
rect 99005 2408 138631 2410
rect 99005 2352 99010 2408
rect 99066 2352 101218 2408
rect 101274 2352 138570 2408
rect 138626 2352 138631 2408
rect 99005 2350 138631 2352
rect 99005 2347 99071 2350
rect 101213 2347 101279 2350
rect 138565 2347 138631 2350
rect 139025 2410 139091 2413
rect 161933 2410 161999 2413
rect 139025 2408 161999 2410
rect 139025 2352 139030 2408
rect 139086 2352 161938 2408
rect 161994 2352 161999 2408
rect 139025 2350 161999 2352
rect 139025 2347 139091 2350
rect 161933 2347 161999 2350
rect 163405 2410 163471 2413
rect 173249 2410 173315 2413
rect 163405 2408 173315 2410
rect 163405 2352 163410 2408
rect 163466 2352 173254 2408
rect 173310 2352 173315 2408
rect 163405 2350 173315 2352
rect 163405 2347 163471 2350
rect 173249 2347 173315 2350
rect 190821 2410 190887 2413
rect 215753 2410 215819 2413
rect 216622 2410 216628 2412
rect 190821 2408 215819 2410
rect 190821 2352 190826 2408
rect 190882 2352 215758 2408
rect 215814 2352 215819 2408
rect 190821 2350 215819 2352
rect 190821 2347 190887 2350
rect 215753 2347 215819 2350
rect 215894 2350 216628 2410
rect 89805 2274 89871 2277
rect 103789 2274 103855 2277
rect 89805 2272 103855 2274
rect 89805 2216 89810 2272
rect 89866 2216 103794 2272
rect 103850 2216 103855 2272
rect 89805 2214 103855 2216
rect 89805 2211 89871 2214
rect 103789 2211 103855 2214
rect 155677 2274 155743 2277
rect 185025 2274 185091 2277
rect 155677 2272 185091 2274
rect 155677 2216 155682 2272
rect 155738 2216 185030 2272
rect 185086 2216 185091 2272
rect 155677 2214 185091 2216
rect 155677 2211 155743 2214
rect 185025 2211 185091 2214
rect 210417 2274 210483 2277
rect 215894 2274 215954 2350
rect 216622 2348 216628 2350
rect 216692 2348 216698 2412
rect 223389 2410 223455 2413
rect 225873 2410 225939 2413
rect 257613 2410 257679 2413
rect 271965 2410 272031 2413
rect 223389 2408 257679 2410
rect 223389 2352 223394 2408
rect 223450 2352 225878 2408
rect 225934 2352 257618 2408
rect 257674 2352 257679 2408
rect 223389 2350 257679 2352
rect 223389 2347 223455 2350
rect 225873 2347 225939 2350
rect 257613 2347 257679 2350
rect 267690 2350 271890 2410
rect 210417 2272 215954 2274
rect 210417 2216 210422 2272
rect 210478 2216 215954 2272
rect 210417 2214 215954 2216
rect 216673 2274 216739 2277
rect 223941 2274 224007 2277
rect 216673 2272 224007 2274
rect 216673 2216 216678 2272
rect 216734 2216 223946 2272
rect 224002 2216 224007 2272
rect 216673 2214 224007 2216
rect 210417 2211 210483 2214
rect 216673 2211 216739 2214
rect 223941 2211 224007 2214
rect 224166 2212 224172 2276
rect 224236 2274 224242 2276
rect 224677 2274 224743 2277
rect 224236 2272 224743 2274
rect 224236 2216 224682 2272
rect 224738 2216 224743 2272
rect 224236 2214 224743 2216
rect 224236 2212 224242 2214
rect 224677 2211 224743 2214
rect 225229 2274 225295 2277
rect 229829 2274 229895 2277
rect 225229 2272 229895 2274
rect 225229 2216 225234 2272
rect 225290 2216 229834 2272
rect 229890 2216 229895 2272
rect 225229 2214 229895 2216
rect 225229 2211 225295 2214
rect 229829 2211 229895 2214
rect 235993 2274 236059 2277
rect 267690 2274 267750 2350
rect 235993 2272 267750 2274
rect 235993 2216 235998 2272
rect 236054 2216 267750 2272
rect 235993 2214 267750 2216
rect 268745 2274 268811 2277
rect 271137 2274 271203 2277
rect 268745 2272 271203 2274
rect 268745 2216 268750 2272
rect 268806 2216 271142 2272
rect 271198 2216 271203 2272
rect 268745 2214 271203 2216
rect 271830 2274 271890 2350
rect 271965 2408 272504 2410
rect 271965 2352 271970 2408
rect 272026 2352 272504 2408
rect 271965 2350 272504 2352
rect 271965 2347 272031 2350
rect 271830 2214 272504 2274
rect 235993 2211 236059 2214
rect 268745 2211 268811 2214
rect 271137 2211 271203 2214
rect 68542 2208 68858 2209
rect 68542 2144 68548 2208
rect 68612 2144 68628 2208
rect 68692 2144 68708 2208
rect 68772 2144 68788 2208
rect 68852 2144 68858 2208
rect 68542 2143 68858 2144
rect 136139 2208 136455 2209
rect 136139 2144 136145 2208
rect 136209 2144 136225 2208
rect 136289 2144 136305 2208
rect 136369 2144 136385 2208
rect 136449 2144 136455 2208
rect 136139 2143 136455 2144
rect 203736 2208 204052 2209
rect 203736 2144 203742 2208
rect 203806 2144 203822 2208
rect 203886 2144 203902 2208
rect 203966 2144 203982 2208
rect 204046 2144 204052 2208
rect 203736 2143 204052 2144
rect 271333 2208 271649 2209
rect 271333 2144 271339 2208
rect 271403 2144 271419 2208
rect 271483 2144 271499 2208
rect 271563 2144 271579 2208
rect 271643 2144 271649 2208
rect 271333 2143 271649 2144
rect 86401 2138 86467 2141
rect 119337 2138 119403 2141
rect 86401 2136 119403 2138
rect 86401 2080 86406 2136
rect 86462 2080 119342 2136
rect 119398 2080 119403 2136
rect 86401 2078 119403 2080
rect 86401 2075 86467 2078
rect 119337 2075 119403 2078
rect 138841 2138 138907 2141
rect 141693 2138 141759 2141
rect 143993 2138 144059 2141
rect 138841 2136 144059 2138
rect 138841 2080 138846 2136
rect 138902 2080 141698 2136
rect 141754 2080 143998 2136
rect 144054 2080 144059 2136
rect 138841 2078 144059 2080
rect 138841 2075 138907 2078
rect 141693 2075 141759 2078
rect 143993 2075 144059 2078
rect 144637 2138 144703 2141
rect 176837 2138 176903 2141
rect 144637 2136 176903 2138
rect 144637 2080 144642 2136
rect 144698 2080 176842 2136
rect 176898 2080 176903 2136
rect 144637 2078 176903 2080
rect 144637 2075 144703 2078
rect 176837 2075 176903 2078
rect 215661 2138 215727 2141
rect 222101 2138 222167 2141
rect 215661 2136 222167 2138
rect 215661 2080 215666 2136
rect 215722 2080 222106 2136
rect 222162 2080 222167 2136
rect 215661 2078 222167 2080
rect 215661 2075 215727 2078
rect 222101 2075 222167 2078
rect 223205 2138 223271 2141
rect 268837 2138 268903 2141
rect 223205 2136 268903 2138
rect 223205 2080 223210 2136
rect 223266 2080 268842 2136
rect 268898 2080 268903 2136
rect 223205 2078 268903 2080
rect 223205 2075 223271 2078
rect 268837 2075 268903 2078
rect 269021 2138 269087 2141
rect 271781 2138 271847 2141
rect 269021 2136 271154 2138
rect 269021 2080 269026 2136
rect 269082 2080 271154 2136
rect 269021 2078 271154 2080
rect 269021 2075 269087 2078
rect 15837 2002 15903 2005
rect 49049 2002 49115 2005
rect 15837 2000 49115 2002
rect 15837 1944 15842 2000
rect 15898 1944 49054 2000
rect 49110 1944 49115 2000
rect 15837 1942 49115 1944
rect 15837 1939 15903 1942
rect 49049 1939 49115 1942
rect 54385 2002 54451 2005
rect 89069 2002 89135 2005
rect 89621 2002 89687 2005
rect 123293 2002 123359 2005
rect 54385 2000 123359 2002
rect 54385 1944 54390 2000
rect 54446 1944 89074 2000
rect 89130 1944 89626 2000
rect 89682 1944 123298 2000
rect 123354 1944 123359 2000
rect 54385 1942 123359 1944
rect 54385 1939 54451 1942
rect 89069 1939 89135 1942
rect 89621 1939 89687 1942
rect 123293 1939 123359 1942
rect 139209 2002 139275 2005
rect 163405 2002 163471 2005
rect 220077 2002 220143 2005
rect 271094 2002 271154 2078
rect 271781 2136 272504 2138
rect 271781 2080 271786 2136
rect 271842 2080 272504 2136
rect 271781 2078 272504 2080
rect 271781 2075 271847 2078
rect 271965 2002 272031 2005
rect 139209 2000 163471 2002
rect 139209 1944 139214 2000
rect 139270 1944 163410 2000
rect 163466 1944 163471 2000
rect 139209 1942 163471 1944
rect 139209 1939 139275 1942
rect 163405 1939 163471 1942
rect 166030 1942 171150 2002
rect 40309 1866 40375 1869
rect 88333 1866 88399 1869
rect 40309 1864 88399 1866
rect 40309 1808 40314 1864
rect 40370 1808 88338 1864
rect 88394 1808 88399 1864
rect 40309 1806 88399 1808
rect 40309 1803 40375 1806
rect 88333 1803 88399 1806
rect 99465 1866 99531 1869
rect 105445 1866 105511 1869
rect 99465 1864 105511 1866
rect 99465 1808 99470 1864
rect 99526 1808 105450 1864
rect 105506 1808 105511 1864
rect 99465 1806 105511 1808
rect 99465 1803 99531 1806
rect 105445 1803 105511 1806
rect 141417 1866 141483 1869
rect 143165 1866 143231 1869
rect 141417 1864 143231 1866
rect 141417 1808 141422 1864
rect 141478 1808 143170 1864
rect 143226 1808 143231 1864
rect 141417 1806 143231 1808
rect 141417 1803 141483 1806
rect 143165 1803 143231 1806
rect 150433 1866 150499 1869
rect 166030 1866 166090 1942
rect 171090 1866 171150 1942
rect 220077 2000 270234 2002
rect 220077 1944 220082 2000
rect 220138 1944 270234 2000
rect 220077 1942 270234 1944
rect 271094 2000 272031 2002
rect 271094 1944 271970 2000
rect 272026 1944 272031 2000
rect 271094 1942 272031 1944
rect 220077 1939 220143 1942
rect 181989 1866 182055 1869
rect 150433 1864 166090 1866
rect 150433 1808 150438 1864
rect 150494 1808 166090 1864
rect 150433 1806 166090 1808
rect 166214 1806 170506 1866
rect 171090 1864 182055 1866
rect 171090 1808 181994 1864
rect 182050 1808 182055 1864
rect 171090 1806 182055 1808
rect 150433 1803 150499 1806
rect 21398 1668 21404 1732
rect 21468 1730 21474 1732
rect 22185 1730 22251 1733
rect 21468 1728 22251 1730
rect 21468 1672 22190 1728
rect 22246 1672 22251 1728
rect 21468 1670 22251 1672
rect 21468 1668 21474 1670
rect 22185 1667 22251 1670
rect 36813 1730 36879 1733
rect 83825 1730 83891 1733
rect 36813 1728 83891 1730
rect 36813 1672 36818 1728
rect 36874 1672 83830 1728
rect 83886 1672 83891 1728
rect 36813 1670 83891 1672
rect 36813 1667 36879 1670
rect 83825 1667 83891 1670
rect 153101 1730 153167 1733
rect 166214 1730 166274 1806
rect 153101 1728 166274 1730
rect 153101 1672 153106 1728
rect 153162 1672 166274 1728
rect 153101 1670 166274 1672
rect 170446 1730 170506 1806
rect 181989 1803 182055 1806
rect 220997 1866 221063 1869
rect 270174 1866 270234 1942
rect 271965 1939 272031 1942
rect 272149 2002 272215 2005
rect 272149 2000 272504 2002
rect 272149 1944 272154 2000
rect 272210 1944 272504 2000
rect 272149 1942 272504 1944
rect 272149 1939 272215 1942
rect 220997 1864 270050 1866
rect 220997 1808 221002 1864
rect 221058 1808 270050 1864
rect 220997 1806 270050 1808
rect 270174 1806 272504 1866
rect 220997 1803 221063 1806
rect 215334 1730 215340 1732
rect 170446 1670 215340 1730
rect 153101 1667 153167 1670
rect 215334 1668 215340 1670
rect 215404 1668 215410 1732
rect 215753 1730 215819 1733
rect 224769 1730 224835 1733
rect 215753 1728 224835 1730
rect 215753 1672 215758 1728
rect 215814 1672 224774 1728
rect 224830 1672 224835 1728
rect 215753 1670 224835 1672
rect 215753 1667 215819 1670
rect 224769 1667 224835 1670
rect 267406 1668 267412 1732
rect 267476 1730 267482 1732
rect 267641 1730 267707 1733
rect 267476 1728 267707 1730
rect 267476 1672 267646 1728
rect 267702 1672 267707 1728
rect 267476 1670 267707 1672
rect 269990 1730 270050 1806
rect 269990 1670 272504 1730
rect 267476 1668 267482 1670
rect 267641 1667 267707 1670
rect 34744 1664 35060 1665
rect 34744 1600 34750 1664
rect 34814 1600 34830 1664
rect 34894 1600 34910 1664
rect 34974 1600 34990 1664
rect 35054 1600 35060 1664
rect 34744 1599 35060 1600
rect 102341 1664 102657 1665
rect 102341 1600 102347 1664
rect 102411 1600 102427 1664
rect 102491 1600 102507 1664
rect 102571 1600 102587 1664
rect 102651 1600 102657 1664
rect 102341 1599 102657 1600
rect 169938 1664 170254 1665
rect 169938 1600 169944 1664
rect 170008 1600 170024 1664
rect 170088 1600 170104 1664
rect 170168 1600 170184 1664
rect 170248 1600 170254 1664
rect 169938 1599 170254 1600
rect 237535 1664 237851 1665
rect 237535 1600 237541 1664
rect 237605 1600 237621 1664
rect 237685 1600 237701 1664
rect 237765 1600 237781 1664
rect 237845 1600 237851 1664
rect 237535 1599 237851 1600
rect 59353 1596 59419 1597
rect 59302 1594 59308 1596
rect 59262 1534 59308 1594
rect 59372 1592 59419 1596
rect 59414 1536 59419 1592
rect 59302 1532 59308 1534
rect 59372 1532 59419 1536
rect 59353 1531 59419 1532
rect 80053 1596 80119 1597
rect 80053 1592 80100 1596
rect 80164 1594 80170 1596
rect 81341 1594 81407 1597
rect 82997 1596 83063 1597
rect 83733 1596 83799 1597
rect 81566 1594 81572 1596
rect 80053 1536 80058 1592
rect 80053 1532 80100 1536
rect 80164 1534 80210 1594
rect 81341 1592 81572 1594
rect 81341 1536 81346 1592
rect 81402 1536 81572 1592
rect 81341 1534 81572 1536
rect 80164 1532 80170 1534
rect 80053 1531 80119 1532
rect 81341 1531 81407 1534
rect 81566 1532 81572 1534
rect 81636 1532 81642 1596
rect 82997 1592 83044 1596
rect 83108 1594 83114 1596
rect 82997 1536 83002 1592
rect 82997 1532 83044 1536
rect 83108 1534 83154 1594
rect 83733 1592 83780 1596
rect 83844 1594 83850 1596
rect 83733 1536 83738 1592
rect 83108 1532 83114 1534
rect 83733 1532 83780 1536
rect 83844 1534 83890 1594
rect 83844 1532 83850 1534
rect 99230 1532 99236 1596
rect 99300 1594 99306 1596
rect 100753 1594 100819 1597
rect 121637 1594 121703 1597
rect 99300 1592 100819 1594
rect 99300 1536 100758 1592
rect 100814 1536 100819 1592
rect 99300 1534 100819 1536
rect 99300 1532 99306 1534
rect 82997 1531 83063 1532
rect 83733 1531 83799 1532
rect 100753 1531 100819 1534
rect 108990 1592 121703 1594
rect 108990 1536 121642 1592
rect 121698 1536 121703 1592
rect 108990 1534 121703 1536
rect 841 1460 907 1461
rect 790 1458 796 1460
rect 750 1398 796 1458
rect 860 1456 907 1460
rect 902 1400 907 1456
rect 790 1396 796 1398
rect 860 1396 907 1400
rect 16246 1396 16252 1460
rect 16316 1458 16322 1460
rect 16573 1458 16639 1461
rect 16316 1456 16639 1458
rect 16316 1400 16578 1456
rect 16634 1400 16639 1456
rect 16316 1398 16639 1400
rect 16316 1396 16322 1398
rect 841 1395 907 1396
rect 16573 1395 16639 1398
rect 20662 1396 20668 1460
rect 20732 1458 20738 1460
rect 22093 1458 22159 1461
rect 20732 1456 22159 1458
rect 20732 1400 22098 1456
rect 22154 1400 22159 1456
rect 20732 1398 22159 1400
rect 20732 1396 20738 1398
rect 22093 1395 22159 1398
rect 32438 1396 32444 1460
rect 32508 1458 32514 1460
rect 33133 1458 33199 1461
rect 32508 1456 33199 1458
rect 32508 1400 33138 1456
rect 33194 1400 33199 1456
rect 32508 1398 33199 1400
rect 32508 1396 32514 1398
rect 33133 1395 33199 1398
rect 53925 1460 53991 1461
rect 53925 1456 53972 1460
rect 54036 1458 54042 1460
rect 54201 1458 54267 1461
rect 89069 1458 89135 1461
rect 108990 1458 109050 1534
rect 121637 1531 121703 1534
rect 155769 1594 155835 1597
rect 156873 1594 156939 1597
rect 155769 1592 156939 1594
rect 155769 1536 155774 1592
rect 155830 1536 156878 1592
rect 156934 1536 156939 1592
rect 155769 1534 156939 1536
rect 155769 1531 155835 1534
rect 156873 1531 156939 1534
rect 191097 1594 191163 1597
rect 191097 1592 200130 1594
rect 191097 1536 191102 1592
rect 191158 1536 200130 1592
rect 191097 1534 200130 1536
rect 191097 1531 191163 1534
rect 117313 1460 117379 1461
rect 128353 1460 128419 1461
rect 117262 1458 117268 1460
rect 53925 1400 53930 1456
rect 53925 1396 53972 1400
rect 54036 1398 54082 1458
rect 54201 1456 109050 1458
rect 54201 1400 54206 1456
rect 54262 1400 89074 1456
rect 89130 1400 109050 1456
rect 54201 1398 109050 1400
rect 117222 1398 117268 1458
rect 117332 1456 117379 1460
rect 128302 1458 128308 1460
rect 117374 1400 117379 1456
rect 54036 1396 54042 1398
rect 53925 1395 53991 1396
rect 54201 1395 54267 1398
rect 89069 1395 89135 1398
rect 117262 1396 117268 1398
rect 117332 1396 117379 1400
rect 128262 1398 128308 1458
rect 128372 1456 128419 1460
rect 128414 1400 128419 1456
rect 128302 1396 128308 1398
rect 128372 1396 128419 1400
rect 134926 1396 134932 1460
rect 134996 1458 135002 1460
rect 135253 1458 135319 1461
rect 134996 1456 135319 1458
rect 134996 1400 135258 1456
rect 135314 1400 135319 1456
rect 134996 1398 135319 1400
rect 134996 1396 135002 1398
rect 117313 1395 117379 1396
rect 128353 1395 128419 1396
rect 135253 1395 135319 1398
rect 137318 1396 137324 1460
rect 137388 1458 137394 1460
rect 138013 1458 138079 1461
rect 137388 1456 138079 1458
rect 137388 1400 138018 1456
rect 138074 1400 138079 1456
rect 137388 1398 138079 1400
rect 137388 1396 137394 1398
rect 138013 1395 138079 1398
rect 144678 1396 144684 1460
rect 144748 1458 144754 1460
rect 144913 1458 144979 1461
rect 144748 1456 144979 1458
rect 144748 1400 144918 1456
rect 144974 1400 144979 1456
rect 144748 1398 144979 1400
rect 144748 1396 144754 1398
rect 144913 1395 144979 1398
rect 155718 1396 155724 1460
rect 155788 1458 155794 1460
rect 155953 1458 156019 1461
rect 155788 1456 156019 1458
rect 155788 1400 155958 1456
rect 156014 1400 156019 1456
rect 155788 1398 156019 1400
rect 155788 1396 155794 1398
rect 155953 1395 156019 1398
rect 156454 1396 156460 1460
rect 156524 1458 156530 1460
rect 157425 1458 157491 1461
rect 156524 1456 157491 1458
rect 156524 1400 157430 1456
rect 157486 1400 157491 1456
rect 156524 1398 157491 1400
rect 156524 1396 156530 1398
rect 157425 1395 157491 1398
rect 157885 1460 157951 1461
rect 157885 1456 157932 1460
rect 157996 1458 158002 1460
rect 157885 1400 157890 1456
rect 157885 1396 157932 1400
rect 157996 1398 158042 1458
rect 157996 1396 158002 1398
rect 163814 1396 163820 1460
rect 163884 1458 163890 1460
rect 164233 1458 164299 1461
rect 163884 1456 164299 1458
rect 163884 1400 164238 1456
rect 164294 1400 164299 1456
rect 163884 1398 164299 1400
rect 163884 1396 163890 1398
rect 157885 1395 157951 1396
rect 164233 1395 164299 1398
rect 168230 1396 168236 1460
rect 168300 1458 168306 1460
rect 168373 1458 168439 1461
rect 186313 1460 186379 1461
rect 186262 1458 186268 1460
rect 168300 1456 168439 1458
rect 168300 1400 168378 1456
rect 168434 1400 168439 1456
rect 168300 1398 168439 1400
rect 186222 1398 186268 1458
rect 186332 1456 186379 1460
rect 186374 1400 186379 1456
rect 168300 1396 168306 1398
rect 168373 1395 168439 1398
rect 186262 1396 186268 1398
rect 186332 1396 186379 1400
rect 194358 1396 194364 1460
rect 194428 1458 194434 1460
rect 194685 1458 194751 1461
rect 194428 1456 194751 1458
rect 194428 1400 194690 1456
rect 194746 1400 194751 1456
rect 194428 1398 194751 1400
rect 194428 1396 194434 1398
rect 186313 1395 186379 1396
rect 194685 1395 194751 1398
rect 195830 1396 195836 1460
rect 195900 1458 195906 1460
rect 195973 1458 196039 1461
rect 195900 1456 196039 1458
rect 195900 1400 195978 1456
rect 196034 1400 196039 1456
rect 195900 1398 196039 1400
rect 200070 1458 200130 1534
rect 201718 1532 201724 1596
rect 201788 1594 201794 1596
rect 202873 1594 202939 1597
rect 223389 1594 223455 1597
rect 201788 1592 202939 1594
rect 201788 1536 202878 1592
rect 202934 1536 202939 1592
rect 201788 1534 202939 1536
rect 201788 1532 201794 1534
rect 202873 1531 202939 1534
rect 215250 1592 223455 1594
rect 215250 1536 223394 1592
rect 223450 1536 223455 1592
rect 215250 1534 223455 1536
rect 215250 1458 215310 1534
rect 223389 1531 223455 1534
rect 223573 1594 223639 1597
rect 235717 1594 235783 1597
rect 223573 1592 235783 1594
rect 223573 1536 223578 1592
rect 223634 1536 235722 1592
rect 235778 1536 235783 1592
rect 223573 1534 235783 1536
rect 223573 1531 223639 1534
rect 235717 1531 235783 1534
rect 269021 1594 269087 1597
rect 269021 1592 272504 1594
rect 269021 1536 269026 1592
rect 269082 1536 272504 1592
rect 269021 1534 272504 1536
rect 269021 1531 269087 1534
rect 216673 1460 216739 1461
rect 216622 1458 216628 1460
rect 200070 1398 215310 1458
rect 216582 1398 216628 1458
rect 216692 1456 216739 1460
rect 216734 1400 216739 1456
rect 195900 1396 195906 1398
rect 195973 1395 196039 1398
rect 216622 1396 216628 1398
rect 216692 1396 216739 1400
rect 220302 1396 220308 1460
rect 220372 1458 220378 1460
rect 220813 1458 220879 1461
rect 224033 1460 224099 1461
rect 223982 1458 223988 1460
rect 220372 1456 220879 1458
rect 220372 1400 220818 1456
rect 220874 1400 220879 1456
rect 220372 1398 220879 1400
rect 223942 1398 223988 1458
rect 224052 1456 224099 1460
rect 224094 1400 224099 1456
rect 220372 1396 220378 1398
rect 216673 1395 216739 1396
rect 220813 1395 220879 1398
rect 223982 1396 223988 1398
rect 224052 1396 224099 1400
rect 225454 1396 225460 1460
rect 225524 1458 225530 1460
rect 225597 1458 225663 1461
rect 237281 1460 237347 1461
rect 237230 1458 237236 1460
rect 225524 1456 225663 1458
rect 225524 1400 225602 1456
rect 225658 1400 225663 1456
rect 225524 1398 225663 1400
rect 237190 1398 237236 1458
rect 237300 1456 237347 1460
rect 237342 1400 237347 1456
rect 225524 1396 225530 1398
rect 224033 1395 224099 1396
rect 225597 1395 225663 1398
rect 237230 1396 237236 1398
rect 237300 1396 237347 1400
rect 242750 1396 242756 1460
rect 242820 1458 242826 1460
rect 242893 1458 242959 1461
rect 242820 1456 242959 1458
rect 242820 1400 242898 1456
rect 242954 1400 242959 1456
rect 242820 1398 242959 1400
rect 242820 1396 242826 1398
rect 237281 1395 237347 1396
rect 242893 1395 242959 1398
rect 244038 1396 244044 1460
rect 244108 1458 244114 1460
rect 244273 1458 244339 1461
rect 244108 1456 244339 1458
rect 244108 1400 244278 1456
rect 244334 1400 244339 1456
rect 244108 1398 244339 1400
rect 244108 1396 244114 1398
rect 244273 1395 244339 1398
rect 247902 1396 247908 1460
rect 247972 1458 247978 1460
rect 248413 1458 248479 1461
rect 247972 1456 248479 1458
rect 247972 1400 248418 1456
rect 248474 1400 248479 1456
rect 247972 1398 248479 1400
rect 247972 1396 247978 1398
rect 248413 1395 248479 1398
rect 249374 1396 249380 1460
rect 249444 1458 249450 1460
rect 249793 1458 249859 1461
rect 249444 1456 249859 1458
rect 249444 1400 249798 1456
rect 249854 1400 249859 1456
rect 249444 1398 249859 1400
rect 249444 1396 249450 1398
rect 249793 1395 249859 1398
rect 250846 1396 250852 1460
rect 250916 1458 250922 1460
rect 251173 1458 251239 1461
rect 250916 1456 251239 1458
rect 250916 1400 251178 1456
rect 251234 1400 251239 1456
rect 250916 1398 251239 1400
rect 250916 1396 250922 1398
rect 251173 1395 251239 1398
rect 264830 1396 264836 1460
rect 264900 1458 264906 1460
rect 264973 1458 265039 1461
rect 264900 1456 265039 1458
rect 264900 1400 264978 1456
rect 265034 1400 265039 1456
rect 264900 1398 265039 1400
rect 264900 1396 264906 1398
rect 264973 1395 265039 1398
rect 268837 1458 268903 1461
rect 268837 1456 272504 1458
rect 268837 1400 268842 1456
rect 268898 1400 272504 1456
rect 268837 1398 272504 1400
rect 268837 1395 268903 1398
rect 1577 1324 1643 1325
rect 1526 1322 1532 1324
rect 1486 1262 1532 1322
rect 1596 1320 1643 1324
rect 1638 1264 1643 1320
rect 1526 1260 1532 1262
rect 1596 1260 1643 1264
rect 25814 1260 25820 1324
rect 25884 1322 25890 1324
rect 25957 1322 26023 1325
rect 25884 1320 26023 1322
rect 25884 1264 25962 1320
rect 26018 1264 26023 1320
rect 25884 1262 26023 1264
rect 25884 1260 25890 1262
rect 1577 1259 1643 1260
rect 25957 1259 26023 1262
rect 26550 1260 26556 1324
rect 26620 1322 26626 1324
rect 26693 1322 26759 1325
rect 26620 1320 26759 1322
rect 26620 1264 26698 1320
rect 26754 1264 26759 1320
rect 26620 1262 26759 1264
rect 26620 1260 26626 1262
rect 26693 1259 26759 1262
rect 27286 1260 27292 1324
rect 27356 1322 27362 1324
rect 27429 1322 27495 1325
rect 71313 1324 71379 1325
rect 73521 1324 73587 1325
rect 76465 1324 76531 1325
rect 77937 1324 78003 1325
rect 79409 1324 79475 1325
rect 71262 1322 71268 1324
rect 27356 1320 27495 1322
rect 27356 1264 27434 1320
rect 27490 1264 27495 1320
rect 27356 1262 27495 1264
rect 71222 1262 71268 1322
rect 71332 1320 71379 1324
rect 73470 1322 73476 1324
rect 71374 1264 71379 1320
rect 27356 1260 27362 1262
rect 27429 1259 27495 1262
rect 71262 1260 71268 1262
rect 71332 1260 71379 1264
rect 73430 1262 73476 1322
rect 73540 1320 73587 1324
rect 76414 1322 76420 1324
rect 73582 1264 73587 1320
rect 73470 1260 73476 1262
rect 73540 1260 73587 1264
rect 76374 1262 76420 1322
rect 76484 1320 76531 1324
rect 77886 1322 77892 1324
rect 76526 1264 76531 1320
rect 76414 1260 76420 1262
rect 76484 1260 76531 1264
rect 77846 1262 77892 1322
rect 77956 1320 78003 1324
rect 79358 1322 79364 1324
rect 77998 1264 78003 1320
rect 77886 1260 77892 1262
rect 77956 1260 78003 1264
rect 79318 1262 79364 1322
rect 79428 1320 79475 1324
rect 79470 1264 79475 1320
rect 79358 1260 79364 1262
rect 79428 1260 79475 1264
rect 71313 1259 71379 1260
rect 73521 1259 73587 1260
rect 76465 1259 76531 1260
rect 77937 1259 78003 1260
rect 79409 1259 79475 1260
rect 82077 1322 82143 1325
rect 87505 1324 87571 1325
rect 82302 1322 82308 1324
rect 82077 1320 82308 1322
rect 82077 1264 82082 1320
rect 82138 1264 82308 1320
rect 82077 1262 82308 1264
rect 82077 1259 82143 1262
rect 82302 1260 82308 1262
rect 82372 1260 82378 1324
rect 87454 1322 87460 1324
rect 87414 1262 87460 1322
rect 87524 1320 87571 1324
rect 87566 1264 87571 1320
rect 87454 1260 87460 1262
rect 87524 1260 87571 1264
rect 88926 1260 88932 1324
rect 88996 1322 89002 1324
rect 89345 1322 89411 1325
rect 88996 1320 89411 1322
rect 88996 1264 89350 1320
rect 89406 1264 89411 1320
rect 88996 1262 89411 1264
rect 88996 1260 89002 1262
rect 87505 1259 87571 1260
rect 89345 1259 89411 1262
rect 97441 1322 97507 1325
rect 104617 1322 104683 1325
rect 97441 1320 104683 1322
rect 97441 1264 97446 1320
rect 97502 1264 104622 1320
rect 104678 1264 104683 1320
rect 97441 1262 104683 1264
rect 97441 1259 97507 1262
rect 104617 1259 104683 1262
rect 140262 1260 140268 1324
rect 140332 1322 140338 1324
rect 140773 1322 140839 1325
rect 140332 1320 140839 1322
rect 140332 1264 140778 1320
rect 140834 1264 140839 1320
rect 140332 1262 140839 1264
rect 140332 1260 140338 1262
rect 140773 1259 140839 1262
rect 154982 1260 154988 1324
rect 155052 1322 155058 1324
rect 155217 1322 155283 1325
rect 155052 1320 155283 1322
rect 155052 1264 155222 1320
rect 155278 1264 155283 1320
rect 155052 1262 155283 1264
rect 155052 1260 155058 1262
rect 155217 1259 155283 1262
rect 156597 1322 156663 1325
rect 169293 1322 169359 1325
rect 156597 1320 169359 1322
rect 156597 1264 156602 1320
rect 156658 1264 169298 1320
rect 169354 1264 169359 1320
rect 156597 1262 169359 1264
rect 156597 1259 156663 1262
rect 169293 1259 169359 1262
rect 176653 1324 176719 1325
rect 179597 1324 179663 1325
rect 181897 1324 181963 1325
rect 176653 1320 176700 1324
rect 176764 1322 176770 1324
rect 176653 1264 176658 1320
rect 176653 1260 176700 1264
rect 176764 1262 176810 1322
rect 179597 1320 179644 1324
rect 179708 1322 179714 1324
rect 181846 1322 181852 1324
rect 179597 1264 179602 1320
rect 176764 1260 176770 1262
rect 179597 1260 179644 1264
rect 179708 1262 179754 1322
rect 181806 1262 181852 1322
rect 181916 1320 181963 1324
rect 181958 1264 181963 1320
rect 179708 1260 179714 1262
rect 181846 1260 181852 1262
rect 181916 1260 181963 1264
rect 176653 1259 176719 1260
rect 179597 1259 179663 1260
rect 181897 1259 181963 1260
rect 186957 1324 187023 1325
rect 186957 1320 187004 1324
rect 187068 1322 187074 1324
rect 186957 1264 186962 1320
rect 186957 1260 187004 1264
rect 187068 1262 187114 1322
rect 187068 1260 187074 1262
rect 199510 1260 199516 1324
rect 199580 1322 199586 1324
rect 199929 1322 199995 1325
rect 199580 1320 199995 1322
rect 199580 1264 199934 1320
rect 199990 1264 199995 1320
rect 199580 1262 199995 1264
rect 199580 1260 199586 1262
rect 186957 1259 187023 1260
rect 199929 1259 199995 1262
rect 210734 1260 210740 1324
rect 210804 1322 210810 1324
rect 211521 1322 211587 1325
rect 210804 1320 211587 1322
rect 210804 1264 211526 1320
rect 211582 1264 211587 1320
rect 210804 1262 211587 1264
rect 210804 1260 210810 1262
rect 211521 1259 211587 1262
rect 222510 1260 222516 1324
rect 222580 1322 222586 1324
rect 222745 1322 222811 1325
rect 222580 1320 222811 1322
rect 222580 1264 222750 1320
rect 222806 1264 222811 1320
rect 222580 1262 222811 1264
rect 222580 1260 222586 1262
rect 222745 1259 222811 1262
rect 226926 1260 226932 1324
rect 226996 1322 227002 1324
rect 227253 1322 227319 1325
rect 226996 1320 227319 1322
rect 226996 1264 227258 1320
rect 227314 1264 227319 1320
rect 226996 1262 227319 1264
rect 226996 1260 227002 1262
rect 227253 1259 227319 1262
rect 227662 1260 227668 1324
rect 227732 1322 227738 1324
rect 228265 1322 228331 1325
rect 227732 1320 228331 1322
rect 227732 1264 228270 1320
rect 228326 1264 228331 1320
rect 227732 1262 228331 1264
rect 227732 1260 227738 1262
rect 228265 1259 228331 1262
rect 234613 1322 234679 1325
rect 241513 1322 241579 1325
rect 234613 1320 241579 1322
rect 234613 1264 234618 1320
rect 234674 1264 241518 1320
rect 241574 1264 241579 1320
rect 234613 1262 241579 1264
rect 234613 1259 234679 1262
rect 241513 1259 241579 1262
rect 268886 1262 272504 1322
rect 10409 1186 10475 1189
rect 85297 1186 85363 1189
rect 87597 1186 87663 1189
rect 88190 1186 88196 1188
rect 10409 1184 16590 1186
rect 10409 1128 10414 1184
rect 10470 1128 16590 1184
rect 10409 1126 16590 1128
rect 10409 1123 10475 1126
rect 2313 1052 2379 1053
rect 4521 1052 4587 1053
rect 2262 1050 2268 1052
rect 2222 990 2268 1050
rect 2332 1048 2379 1052
rect 4470 1050 4476 1052
rect 2374 992 2379 1048
rect 2262 988 2268 990
rect 2332 988 2379 992
rect 4430 990 4476 1050
rect 4540 1048 4587 1052
rect 4582 992 4587 1048
rect 4470 988 4476 990
rect 4540 988 4587 992
rect 6678 988 6684 1052
rect 6748 1050 6754 1052
rect 6821 1050 6887 1053
rect 14089 1052 14155 1053
rect 14038 1050 14044 1052
rect 6748 1048 6887 1050
rect 6748 992 6826 1048
rect 6882 992 6887 1048
rect 6748 990 6887 992
rect 13998 990 14044 1050
rect 14108 1048 14155 1052
rect 14150 992 14155 1048
rect 6748 988 6754 990
rect 2313 987 2379 988
rect 4521 987 4587 988
rect 6821 987 6887 990
rect 14038 988 14044 990
rect 14108 988 14155 992
rect 16530 1050 16590 1126
rect 85297 1184 87522 1186
rect 85297 1128 85302 1184
rect 85358 1128 87522 1184
rect 85297 1126 87522 1128
rect 85297 1123 85363 1126
rect 68542 1120 68858 1121
rect 68542 1056 68548 1120
rect 68612 1056 68628 1120
rect 68692 1056 68708 1120
rect 68772 1056 68788 1120
rect 68852 1056 68858 1120
rect 68542 1055 68858 1056
rect 44357 1050 44423 1053
rect 70577 1052 70643 1053
rect 72049 1052 72115 1053
rect 74257 1052 74323 1053
rect 75729 1052 75795 1053
rect 77201 1052 77267 1053
rect 70526 1050 70532 1052
rect 16530 1048 44423 1050
rect 16530 992 44362 1048
rect 44418 992 44423 1048
rect 16530 990 44423 992
rect 70486 990 70532 1050
rect 70596 1048 70643 1052
rect 71998 1050 72004 1052
rect 70638 992 70643 1048
rect 14089 987 14155 988
rect 44357 987 44423 990
rect 70526 988 70532 990
rect 70596 988 70643 992
rect 71958 990 72004 1050
rect 72068 1048 72115 1052
rect 74206 1050 74212 1052
rect 72110 992 72115 1048
rect 71998 988 72004 990
rect 72068 988 72115 992
rect 74166 990 74212 1050
rect 74276 1048 74323 1052
rect 75678 1050 75684 1052
rect 74318 992 74323 1048
rect 74206 988 74212 990
rect 74276 988 74323 992
rect 75638 990 75684 1050
rect 75748 1048 75795 1052
rect 77150 1050 77156 1052
rect 75790 992 75795 1048
rect 75678 988 75684 990
rect 75748 988 75795 992
rect 77110 990 77156 1050
rect 77220 1048 77267 1052
rect 77262 992 77267 1048
rect 77150 988 77156 990
rect 77220 988 77267 992
rect 85982 988 85988 1052
rect 86052 1050 86058 1052
rect 86125 1050 86191 1053
rect 86052 1048 86191 1050
rect 86052 992 86130 1048
rect 86186 992 86191 1048
rect 86052 990 86191 992
rect 87462 1050 87522 1126
rect 87597 1184 88196 1186
rect 87597 1128 87602 1184
rect 87658 1128 88196 1184
rect 87597 1126 88196 1128
rect 87597 1123 87663 1126
rect 88190 1124 88196 1126
rect 88260 1124 88266 1188
rect 93853 1186 93919 1189
rect 94078 1186 94084 1188
rect 93853 1184 94084 1186
rect 93853 1128 93858 1184
rect 93914 1128 94084 1184
rect 93853 1126 94084 1128
rect 93853 1123 93919 1126
rect 94078 1124 94084 1126
rect 94148 1124 94154 1188
rect 94589 1186 94655 1189
rect 94814 1186 94820 1188
rect 94589 1184 94820 1186
rect 94589 1128 94594 1184
rect 94650 1128 94820 1184
rect 94589 1126 94820 1128
rect 94589 1123 94655 1126
rect 94814 1124 94820 1126
rect 94884 1124 94890 1188
rect 95325 1186 95391 1189
rect 95550 1186 95556 1188
rect 95325 1184 95556 1186
rect 95325 1128 95330 1184
rect 95386 1128 95556 1184
rect 95325 1126 95556 1128
rect 95325 1123 95391 1126
rect 95550 1124 95556 1126
rect 95620 1124 95626 1188
rect 96061 1186 96127 1189
rect 96286 1186 96292 1188
rect 96061 1184 96292 1186
rect 96061 1128 96066 1184
rect 96122 1128 96292 1184
rect 96061 1126 96292 1128
rect 96061 1123 96127 1126
rect 96286 1124 96292 1126
rect 96356 1124 96362 1188
rect 100569 1186 100635 1189
rect 106825 1186 106891 1189
rect 100569 1184 106891 1186
rect 100569 1128 100574 1184
rect 100630 1128 106830 1184
rect 106886 1128 106891 1184
rect 100569 1126 106891 1128
rect 100569 1123 100635 1126
rect 106825 1123 106891 1126
rect 160134 1124 160140 1188
rect 160204 1186 160210 1188
rect 160921 1186 160987 1189
rect 160204 1184 160987 1186
rect 160204 1128 160926 1184
rect 160982 1128 160987 1184
rect 160204 1126 160987 1128
rect 160204 1124 160210 1126
rect 160921 1123 160987 1126
rect 161606 1124 161612 1188
rect 161676 1186 161682 1188
rect 161749 1186 161815 1189
rect 161676 1184 161815 1186
rect 161676 1128 161754 1184
rect 161810 1128 161815 1184
rect 161676 1126 161815 1128
rect 161676 1124 161682 1126
rect 161749 1123 161815 1126
rect 163078 1124 163084 1188
rect 163148 1186 163154 1188
rect 163865 1186 163931 1189
rect 165337 1188 165403 1189
rect 166073 1188 166139 1189
rect 166809 1188 166875 1189
rect 165286 1186 165292 1188
rect 163148 1184 163931 1186
rect 163148 1128 163870 1184
rect 163926 1128 163931 1184
rect 163148 1126 163931 1128
rect 165246 1126 165292 1186
rect 165356 1184 165403 1188
rect 166022 1186 166028 1188
rect 165398 1128 165403 1184
rect 163148 1124 163154 1126
rect 163865 1123 163931 1126
rect 165286 1124 165292 1126
rect 165356 1124 165403 1128
rect 165982 1126 166028 1186
rect 166092 1184 166139 1188
rect 166758 1186 166764 1188
rect 166134 1128 166139 1184
rect 166022 1124 166028 1126
rect 166092 1124 166139 1128
rect 166718 1126 166764 1186
rect 166828 1184 166875 1188
rect 166870 1128 166875 1184
rect 166758 1124 166764 1126
rect 166828 1124 166875 1128
rect 165337 1123 165403 1124
rect 166073 1123 166139 1124
rect 166809 1123 166875 1124
rect 171409 1186 171475 1189
rect 181897 1186 181963 1189
rect 184565 1186 184631 1189
rect 171409 1184 181963 1186
rect 171409 1128 171414 1184
rect 171470 1128 181902 1184
rect 181958 1128 181963 1184
rect 171409 1126 181963 1128
rect 171409 1123 171475 1126
rect 181897 1123 181963 1126
rect 182590 1184 184631 1186
rect 182590 1128 184570 1184
rect 184626 1128 184631 1184
rect 182590 1126 184631 1128
rect 136139 1120 136455 1121
rect 136139 1056 136145 1120
rect 136209 1056 136225 1120
rect 136289 1056 136305 1120
rect 136369 1056 136385 1120
rect 136449 1056 136455 1120
rect 136139 1055 136455 1056
rect 118417 1050 118483 1053
rect 87462 1048 118483 1050
rect 87462 992 118422 1048
rect 118478 992 118483 1048
rect 87462 990 118483 992
rect 86052 988 86058 990
rect 70577 987 70643 988
rect 72049 987 72115 988
rect 74257 987 74323 988
rect 75729 987 75795 988
rect 77201 987 77267 988
rect 86125 987 86191 990
rect 118417 987 118483 990
rect 142470 988 142476 1052
rect 142540 1050 142546 1052
rect 142981 1050 143047 1053
rect 142540 1048 143047 1050
rect 142540 992 142986 1048
rect 143042 992 143047 1048
rect 142540 990 143047 992
rect 142540 988 142546 990
rect 142981 987 143047 990
rect 149830 988 149836 1052
rect 149900 1050 149906 1052
rect 150065 1050 150131 1053
rect 149900 1048 150131 1050
rect 149900 992 150070 1048
rect 150126 992 150131 1048
rect 149900 990 150131 992
rect 149900 988 149906 990
rect 150065 987 150131 990
rect 151721 1050 151787 1053
rect 182590 1050 182650 1126
rect 184565 1123 184631 1126
rect 190678 1124 190684 1188
rect 190748 1186 190754 1188
rect 191281 1186 191347 1189
rect 190748 1184 191347 1186
rect 190748 1128 191286 1184
rect 191342 1128 191347 1184
rect 190748 1126 191347 1128
rect 190748 1124 190754 1126
rect 191281 1123 191347 1126
rect 198038 1124 198044 1188
rect 198108 1186 198114 1188
rect 198549 1186 198615 1189
rect 198108 1184 198615 1186
rect 198108 1128 198554 1184
rect 198610 1128 198615 1184
rect 198108 1126 198615 1128
rect 198108 1124 198114 1126
rect 198549 1123 198615 1126
rect 200982 1124 200988 1188
rect 201052 1186 201058 1188
rect 201401 1186 201467 1189
rect 201052 1184 201467 1186
rect 201052 1128 201406 1184
rect 201462 1128 201467 1184
rect 201052 1126 201467 1128
rect 201052 1124 201058 1126
rect 201401 1123 201467 1126
rect 218513 1186 218579 1189
rect 222377 1186 222443 1189
rect 228449 1188 228515 1189
rect 228398 1186 228404 1188
rect 218513 1184 222443 1186
rect 218513 1128 218518 1184
rect 218574 1128 222382 1184
rect 222438 1128 222443 1184
rect 218513 1126 222443 1128
rect 228358 1126 228404 1186
rect 228468 1184 228515 1188
rect 228510 1128 228515 1184
rect 218513 1123 218579 1126
rect 222377 1123 222443 1126
rect 228398 1124 228404 1126
rect 228468 1124 228515 1128
rect 228449 1123 228515 1124
rect 231301 1188 231367 1189
rect 232037 1188 232103 1189
rect 232773 1188 232839 1189
rect 231301 1184 231348 1188
rect 231412 1186 231418 1188
rect 231301 1128 231306 1184
rect 231301 1124 231348 1128
rect 231412 1126 231458 1186
rect 232037 1184 232084 1188
rect 232148 1186 232154 1188
rect 232037 1128 232042 1184
rect 231412 1124 231418 1126
rect 232037 1124 232084 1128
rect 232148 1126 232194 1186
rect 232773 1184 232820 1188
rect 232884 1186 232890 1188
rect 232773 1128 232778 1184
rect 232148 1124 232154 1126
rect 232773 1124 232820 1128
rect 232884 1126 232930 1186
rect 232884 1124 232890 1126
rect 236494 1124 236500 1188
rect 236564 1186 236570 1188
rect 236729 1186 236795 1189
rect 236564 1184 236795 1186
rect 236564 1128 236734 1184
rect 236790 1128 236795 1184
rect 236564 1126 236795 1128
rect 236564 1124 236570 1126
rect 231301 1123 231367 1124
rect 232037 1123 232103 1124
rect 232773 1123 232839 1124
rect 236729 1123 236795 1126
rect 247166 1124 247172 1188
rect 247236 1186 247242 1188
rect 248505 1186 248571 1189
rect 247236 1184 248571 1186
rect 247236 1128 248510 1184
rect 248566 1128 248571 1184
rect 247236 1126 248571 1128
rect 247236 1124 247242 1126
rect 248505 1123 248571 1126
rect 203736 1120 204052 1121
rect 203736 1056 203742 1120
rect 203806 1056 203822 1120
rect 203886 1056 203902 1120
rect 203966 1056 203982 1120
rect 204046 1056 204052 1120
rect 203736 1055 204052 1056
rect 151721 1048 182650 1050
rect 151721 992 151726 1048
rect 151782 992 182650 1048
rect 151721 990 182650 992
rect 183277 1052 183343 1053
rect 184749 1052 184815 1053
rect 183277 1048 183324 1052
rect 183388 1050 183394 1052
rect 183277 992 183282 1048
rect 151721 987 151787 990
rect 183277 988 183324 992
rect 183388 990 183434 1050
rect 184749 1048 184796 1052
rect 184860 1050 184866 1052
rect 184749 992 184754 1048
rect 183388 988 183394 990
rect 184749 988 184796 992
rect 184860 990 184906 1050
rect 184860 988 184866 990
rect 187734 988 187740 1052
rect 187804 1050 187810 1052
rect 188153 1050 188219 1053
rect 187804 1048 188219 1050
rect 187804 992 188158 1048
rect 188214 992 188219 1048
rect 187804 990 188219 992
rect 187804 988 187810 990
rect 183277 987 183343 988
rect 184749 987 184815 988
rect 188153 987 188219 990
rect 189206 988 189212 1052
rect 189276 1050 189282 1052
rect 189441 1050 189507 1053
rect 189276 1048 189507 1050
rect 189276 992 189446 1048
rect 189502 992 189507 1048
rect 189276 990 189507 992
rect 189276 988 189282 990
rect 189441 987 189507 990
rect 209998 988 210004 1052
rect 210068 1050 210074 1052
rect 210877 1050 210943 1053
rect 210068 1048 210943 1050
rect 210068 992 210882 1048
rect 210938 992 210943 1048
rect 210068 990 210943 992
rect 210068 988 210074 990
rect 210877 987 210943 990
rect 211470 988 211476 1052
rect 211540 1050 211546 1052
rect 211705 1050 211771 1053
rect 211540 1048 211771 1050
rect 211540 992 211710 1048
rect 211766 992 211771 1048
rect 211540 990 211771 992
rect 211540 988 211546 990
rect 211705 987 211771 990
rect 218973 1050 219039 1053
rect 268745 1050 268811 1053
rect 218973 1048 268811 1050
rect 218973 992 218978 1048
rect 219034 992 268750 1048
rect 268806 992 268811 1048
rect 218973 990 268811 992
rect 218973 987 219039 990
rect 268745 987 268811 990
rect 77569 914 77635 917
rect 100569 914 100635 917
rect 77569 912 100635 914
rect 77569 856 77574 912
rect 77630 856 100574 912
rect 100630 856 100635 912
rect 77569 854 100635 856
rect 77569 851 77635 854
rect 100569 851 100635 854
rect 100702 852 100708 916
rect 100772 914 100778 916
rect 101305 914 101371 917
rect 120901 914 120967 917
rect 100772 912 101371 914
rect 100772 856 101310 912
rect 101366 856 101371 912
rect 100772 854 101371 856
rect 100772 852 100778 854
rect 101305 851 101371 854
rect 113130 912 120967 914
rect 113130 856 120906 912
rect 120962 856 120967 912
rect 113130 854 120967 856
rect 2957 780 3023 781
rect 5165 780 5231 781
rect 2957 776 3004 780
rect 3068 778 3074 780
rect 2957 720 2962 776
rect 2957 716 3004 720
rect 3068 718 3114 778
rect 5165 776 5212 780
rect 5276 778 5282 780
rect 5165 720 5170 776
rect 3068 716 3074 718
rect 5165 716 5212 720
rect 5276 718 5322 778
rect 5276 716 5282 718
rect 5942 716 5948 780
rect 6012 778 6018 780
rect 6545 778 6611 781
rect 6012 776 6611 778
rect 6012 720 6550 776
rect 6606 720 6611 776
rect 6012 718 6611 720
rect 6012 716 6018 718
rect 2957 715 3023 716
rect 5165 715 5231 716
rect 6545 715 6611 718
rect 7414 716 7420 780
rect 7484 778 7490 780
rect 7557 778 7623 781
rect 7484 776 7623 778
rect 7484 720 7562 776
rect 7618 720 7623 776
rect 7484 718 7623 720
rect 7484 716 7490 718
rect 7557 715 7623 718
rect 8886 716 8892 780
rect 8956 778 8962 780
rect 9029 778 9095 781
rect 14825 780 14891 781
rect 14774 778 14780 780
rect 8956 776 9095 778
rect 8956 720 9034 776
rect 9090 720 9095 776
rect 8956 718 9095 720
rect 14734 718 14780 778
rect 14844 776 14891 780
rect 14886 720 14891 776
rect 8956 716 8962 718
rect 9029 715 9095 718
rect 14774 716 14780 718
rect 14844 716 14891 720
rect 15510 716 15516 780
rect 15580 778 15586 780
rect 15653 778 15719 781
rect 69105 780 69171 781
rect 69054 778 69060 780
rect 15580 776 15719 778
rect 15580 720 15658 776
rect 15714 720 15719 776
rect 15580 718 15719 720
rect 69014 718 69060 778
rect 69124 776 69171 780
rect 69166 720 69171 776
rect 15580 716 15586 718
rect 14825 715 14891 716
rect 15653 715 15719 718
rect 69054 716 69060 718
rect 69124 716 69171 720
rect 69105 715 69171 716
rect 69565 778 69631 781
rect 78581 780 78647 781
rect 69790 778 69796 780
rect 69565 776 69796 778
rect 69565 720 69570 776
rect 69626 720 69796 776
rect 69565 718 69796 720
rect 69565 715 69631 718
rect 69790 716 69796 718
rect 69860 716 69866 780
rect 78581 776 78628 780
rect 78692 778 78698 780
rect 79961 778 80027 781
rect 84469 780 84535 781
rect 80830 778 80836 780
rect 78581 720 78586 776
rect 78581 716 78628 720
rect 78692 718 78738 778
rect 79961 776 80836 778
rect 79961 720 79966 776
rect 80022 720 80836 776
rect 79961 718 80836 720
rect 78692 716 78698 718
rect 78581 715 78647 716
rect 79961 715 80027 718
rect 80830 716 80836 718
rect 80900 716 80906 780
rect 84469 776 84516 780
rect 84580 778 84586 780
rect 85021 778 85087 781
rect 86769 780 86835 781
rect 85246 778 85252 780
rect 84469 720 84474 776
rect 84469 716 84516 720
rect 84580 718 84626 778
rect 85021 776 85252 778
rect 85021 720 85026 776
rect 85082 720 85252 776
rect 85021 718 85252 720
rect 84580 716 84586 718
rect 84469 715 84535 716
rect 85021 715 85087 718
rect 85246 716 85252 718
rect 85316 716 85322 780
rect 86718 778 86724 780
rect 86678 718 86724 778
rect 86788 776 86835 780
rect 86830 720 86835 776
rect 86718 716 86724 718
rect 86788 716 86835 720
rect 90398 716 90404 780
rect 90468 778 90474 780
rect 90633 778 90699 781
rect 90468 776 90699 778
rect 90468 720 90638 776
rect 90694 720 90699 776
rect 90468 718 90699 720
rect 90468 716 90474 718
rect 86769 715 86835 716
rect 90633 715 90699 718
rect 91870 716 91876 780
rect 91940 778 91946 780
rect 92197 778 92263 781
rect 91940 776 92263 778
rect 91940 720 92202 776
rect 92258 720 92263 776
rect 91940 718 92263 720
rect 91940 716 91946 718
rect 92197 715 92263 718
rect 93342 716 93348 780
rect 93412 778 93418 780
rect 93485 778 93551 781
rect 93412 776 93551 778
rect 93412 720 93490 776
rect 93546 720 93551 776
rect 93412 718 93551 720
rect 93412 716 93418 718
rect 93485 715 93551 718
rect 97073 778 97139 781
rect 98453 780 98519 781
rect 97758 778 97764 780
rect 97073 776 97764 778
rect 97073 720 97078 776
rect 97134 720 97764 776
rect 97073 718 97764 720
rect 97073 715 97139 718
rect 97758 716 97764 718
rect 97828 716 97834 780
rect 98453 776 98500 780
rect 98564 778 98570 780
rect 98729 778 98795 781
rect 113130 778 113190 854
rect 120901 851 120967 854
rect 147029 914 147095 917
rect 171409 914 171475 917
rect 147029 912 171475 914
rect 147029 856 147034 912
rect 147090 856 171414 912
rect 171470 856 171475 912
rect 147029 854 171475 856
rect 147029 851 147095 854
rect 171409 851 171475 854
rect 171542 852 171548 916
rect 171612 914 171618 916
rect 171685 914 171751 917
rect 171612 912 171751 914
rect 171612 856 171690 912
rect 171746 856 171751 912
rect 171612 854 171751 856
rect 171612 852 171618 854
rect 171685 851 171751 854
rect 172237 916 172303 917
rect 172973 916 173039 917
rect 173801 916 173867 917
rect 172237 912 172284 916
rect 172348 914 172354 916
rect 172237 856 172242 912
rect 172237 852 172284 856
rect 172348 854 172394 914
rect 172973 912 173020 916
rect 173084 914 173090 916
rect 173750 914 173756 916
rect 172973 856 172978 912
rect 172348 852 172354 854
rect 172973 852 173020 856
rect 173084 854 173130 914
rect 173710 854 173756 914
rect 173820 912 173867 916
rect 173862 856 173867 912
rect 173084 852 173090 854
rect 173750 852 173756 854
rect 173820 852 173867 856
rect 172237 851 172303 852
rect 172973 851 173039 852
rect 173801 851 173867 852
rect 174445 916 174511 917
rect 175181 916 175247 917
rect 174445 912 174492 916
rect 174556 914 174562 916
rect 174445 856 174450 912
rect 174445 852 174492 856
rect 174556 854 174602 914
rect 175181 912 175228 916
rect 175292 914 175298 916
rect 175181 856 175186 912
rect 174556 852 174562 854
rect 175181 852 175228 856
rect 175292 854 175338 914
rect 175292 852 175298 854
rect 175958 852 175964 916
rect 176028 914 176034 916
rect 176561 914 176627 917
rect 176028 912 176627 914
rect 176028 856 176566 912
rect 176622 856 176627 912
rect 176028 854 176627 856
rect 176028 852 176034 854
rect 174445 851 174511 852
rect 175181 851 175247 852
rect 176561 851 176627 854
rect 177430 852 177436 916
rect 177500 914 177506 916
rect 177849 914 177915 917
rect 177500 912 177915 914
rect 177500 856 177854 912
rect 177910 856 177915 912
rect 177500 854 177915 856
rect 177500 852 177506 854
rect 177849 851 177915 854
rect 178166 852 178172 916
rect 178236 914 178242 916
rect 178401 914 178467 917
rect 178236 912 178467 914
rect 178236 856 178406 912
rect 178462 856 178467 912
rect 178236 854 178467 856
rect 178236 852 178242 854
rect 178401 851 178467 854
rect 178902 852 178908 916
rect 178972 914 178978 916
rect 179137 914 179203 917
rect 178972 912 179203 914
rect 178972 856 179142 912
rect 179198 856 179203 912
rect 178972 854 179203 856
rect 178972 852 178978 854
rect 179137 851 179203 854
rect 180374 852 180380 916
rect 180444 914 180450 916
rect 180517 914 180583 917
rect 180444 912 180583 914
rect 180444 856 180522 912
rect 180578 856 180583 912
rect 180444 854 180583 856
rect 180444 852 180450 854
rect 180517 851 180583 854
rect 181110 852 181116 916
rect 181180 914 181186 916
rect 181805 914 181871 917
rect 181180 912 181871 914
rect 181180 856 181810 912
rect 181866 856 181871 912
rect 181180 854 181871 856
rect 181180 852 181186 854
rect 181805 851 181871 854
rect 182541 916 182607 917
rect 182541 912 182588 916
rect 182652 914 182658 916
rect 182541 856 182546 912
rect 182541 852 182588 856
rect 182652 854 182698 914
rect 182652 852 182658 854
rect 184054 852 184060 916
rect 184124 914 184130 916
rect 184289 914 184355 917
rect 185577 916 185643 917
rect 188521 916 188587 917
rect 185526 914 185532 916
rect 184124 912 184355 914
rect 184124 856 184294 912
rect 184350 856 184355 912
rect 184124 854 184355 856
rect 185486 854 185532 914
rect 185596 912 185643 916
rect 188470 914 188476 916
rect 185638 856 185643 912
rect 184124 852 184130 854
rect 182541 851 182607 852
rect 184289 851 184355 854
rect 185526 852 185532 854
rect 185596 852 185643 856
rect 188430 854 188476 914
rect 188540 912 188587 916
rect 188582 856 188587 912
rect 188470 852 188476 854
rect 188540 852 188587 856
rect 192150 852 192156 916
rect 192220 914 192226 916
rect 192661 914 192727 917
rect 192937 916 193003 917
rect 193673 916 193739 917
rect 192886 914 192892 916
rect 192220 912 192727 914
rect 192220 856 192666 912
rect 192722 856 192727 912
rect 192220 854 192727 856
rect 192846 854 192892 914
rect 192956 912 193003 916
rect 193622 914 193628 916
rect 192998 856 193003 912
rect 192220 852 192226 854
rect 185577 851 185643 852
rect 188521 851 188587 852
rect 192661 851 192727 854
rect 192886 852 192892 854
rect 192956 852 193003 856
rect 193582 854 193628 914
rect 193692 912 193739 916
rect 193734 856 193739 912
rect 193622 852 193628 854
rect 193692 852 193739 856
rect 195094 852 195100 916
rect 195164 914 195170 916
rect 195789 914 195855 917
rect 196617 916 196683 917
rect 196566 914 196572 916
rect 195164 912 195855 914
rect 195164 856 195794 912
rect 195850 856 195855 912
rect 195164 854 195855 856
rect 196526 854 196572 914
rect 196636 912 196683 916
rect 196678 856 196683 912
rect 195164 852 195170 854
rect 192937 851 193003 852
rect 193673 851 193739 852
rect 195789 851 195855 854
rect 196566 852 196572 854
rect 196636 852 196683 856
rect 196617 851 196683 852
rect 197261 916 197327 917
rect 197261 912 197308 916
rect 197372 914 197378 916
rect 197261 856 197266 912
rect 197261 852 197308 856
rect 197372 854 197418 914
rect 197372 852 197378 854
rect 198774 852 198780 916
rect 198844 914 198850 916
rect 199929 914 199995 917
rect 198844 912 199995 914
rect 198844 856 199934 912
rect 199990 856 199995 912
rect 198844 854 199995 856
rect 198844 852 198850 854
rect 197261 851 197327 852
rect 199929 851 199995 854
rect 200246 852 200252 916
rect 200316 914 200322 916
rect 200665 914 200731 917
rect 200316 912 200731 914
rect 200316 856 200670 912
rect 200726 856 200731 912
rect 200316 854 200731 856
rect 200316 852 200322 854
rect 200665 851 200731 854
rect 203190 852 203196 916
rect 203260 914 203266 916
rect 203333 914 203399 917
rect 205817 916 205883 917
rect 205766 914 205772 916
rect 203260 912 203399 914
rect 203260 856 203338 912
rect 203394 856 203399 912
rect 203260 854 203399 856
rect 205726 854 205772 914
rect 205836 912 205883 916
rect 205878 856 205883 912
rect 203260 852 203266 854
rect 203333 851 203399 854
rect 205766 852 205772 854
rect 205836 852 205883 856
rect 206318 852 206324 916
rect 206388 914 206394 916
rect 206553 914 206619 917
rect 206388 912 206619 914
rect 206388 856 206558 912
rect 206614 856 206619 912
rect 206388 854 206619 856
rect 206388 852 206394 854
rect 205817 851 205883 852
rect 206553 851 206619 854
rect 207054 852 207060 916
rect 207124 914 207130 916
rect 207657 914 207723 917
rect 207124 912 207723 914
rect 207124 856 207662 912
rect 207718 856 207723 912
rect 207124 854 207723 856
rect 207124 852 207130 854
rect 207657 851 207723 854
rect 207790 852 207796 916
rect 207860 914 207866 916
rect 208301 914 208367 917
rect 207860 912 208367 914
rect 207860 856 208306 912
rect 208362 856 208367 912
rect 207860 854 208367 856
rect 207860 852 207866 854
rect 208301 851 208367 854
rect 208526 852 208532 916
rect 208596 914 208602 916
rect 208945 914 209011 917
rect 208596 912 209011 914
rect 208596 856 208950 912
rect 209006 856 209011 912
rect 208596 854 209011 856
rect 208596 852 208602 854
rect 208945 851 209011 854
rect 209262 852 209268 916
rect 209332 914 209338 916
rect 209773 914 209839 917
rect 212257 916 212323 917
rect 212206 914 212212 916
rect 209332 912 209839 914
rect 209332 856 209778 912
rect 209834 856 209839 912
rect 209332 854 209839 856
rect 212166 854 212212 914
rect 212276 912 212323 916
rect 212318 856 212323 912
rect 209332 852 209338 854
rect 209773 851 209839 854
rect 212206 852 212212 854
rect 212276 852 212323 856
rect 212942 852 212948 916
rect 213012 914 213018 916
rect 213453 914 213519 917
rect 213729 916 213795 917
rect 214465 916 214531 917
rect 213678 914 213684 916
rect 213012 912 213519 914
rect 213012 856 213458 912
rect 213514 856 213519 912
rect 213012 854 213519 856
rect 213638 854 213684 914
rect 213748 912 213795 916
rect 214414 914 214420 916
rect 213790 856 213795 912
rect 213012 852 213018 854
rect 212257 851 212323 852
rect 213453 851 213519 854
rect 213678 852 213684 854
rect 213748 852 213795 856
rect 214374 854 214420 914
rect 214484 912 214531 916
rect 214526 856 214531 912
rect 214414 852 214420 854
rect 214484 852 214531 856
rect 213729 851 213795 852
rect 214465 851 214531 852
rect 215109 916 215175 917
rect 215109 912 215156 916
rect 215220 914 215226 916
rect 215109 856 215114 912
rect 215109 852 215156 856
rect 215220 854 215266 914
rect 215220 852 215226 854
rect 215886 852 215892 916
rect 215956 914 215962 916
rect 216673 914 216739 917
rect 217409 916 217475 917
rect 217358 914 217364 916
rect 215956 912 216739 914
rect 215956 856 216678 912
rect 216734 856 216739 912
rect 215956 854 216739 856
rect 217318 854 217364 914
rect 217428 912 217475 916
rect 217470 856 217475 912
rect 215956 852 215962 854
rect 215109 851 215175 852
rect 216673 851 216739 854
rect 217358 852 217364 854
rect 217428 852 217475 856
rect 218094 852 218100 916
rect 218164 914 218170 916
rect 219433 914 219499 917
rect 218164 912 219499 914
rect 218164 856 219438 912
rect 219494 856 219499 912
rect 218164 854 219499 856
rect 218164 852 218170 854
rect 217409 851 217475 852
rect 219433 851 219499 854
rect 221038 852 221044 916
rect 221108 914 221114 916
rect 222193 914 222259 917
rect 221108 912 222259 914
rect 221108 856 222198 912
rect 222254 856 222259 912
rect 221108 854 222259 856
rect 221108 852 221114 854
rect 222193 851 222259 854
rect 222377 914 222443 917
rect 248045 914 248111 917
rect 258073 914 258139 917
rect 222377 912 248111 914
rect 222377 856 222382 912
rect 222438 856 248050 912
rect 248106 856 248111 912
rect 222377 854 248111 856
rect 222377 851 222443 854
rect 248045 851 248111 854
rect 248370 912 258139 914
rect 248370 856 258078 912
rect 258134 856 258139 912
rect 248370 854 258139 856
rect 117589 778 117655 781
rect 138841 780 138907 781
rect 138790 778 138796 780
rect 98453 720 98458 776
rect 98453 716 98500 720
rect 98564 718 98610 778
rect 98729 776 113190 778
rect 98729 720 98734 776
rect 98790 720 113190 776
rect 98729 718 113190 720
rect 113406 776 117655 778
rect 113406 720 117594 776
rect 117650 720 117655 776
rect 113406 718 117655 720
rect 138750 718 138796 778
rect 138860 776 138907 780
rect 138902 720 138907 776
rect 98564 716 98570 718
rect 98453 715 98519 716
rect 98729 715 98795 718
rect 3734 580 3740 644
rect 3804 642 3810 644
rect 4061 642 4127 645
rect 8201 644 8267 645
rect 8150 642 8156 644
rect 3804 640 4127 642
rect 3804 584 4066 640
rect 4122 584 4127 640
rect 3804 582 4127 584
rect 8110 582 8156 642
rect 8220 640 8267 644
rect 8262 584 8267 640
rect 3804 580 3810 582
rect 4061 579 4127 582
rect 8150 580 8156 582
rect 8220 580 8267 584
rect 8201 579 8267 580
rect 9581 644 9647 645
rect 9581 640 9628 644
rect 9692 642 9698 644
rect 10225 642 10291 645
rect 10358 642 10364 644
rect 9581 584 9586 640
rect 9581 580 9628 584
rect 9692 582 9738 642
rect 10225 640 10364 642
rect 10225 584 10230 640
rect 10286 584 10364 640
rect 10225 582 10364 584
rect 9692 580 9698 582
rect 9581 579 9647 580
rect 10225 579 10291 582
rect 10358 580 10364 582
rect 10428 580 10434 644
rect 10961 642 11027 645
rect 11094 642 11100 644
rect 10961 640 11100 642
rect 10961 584 10966 640
rect 11022 584 11100 640
rect 10961 582 11100 584
rect 10961 579 11027 582
rect 11094 580 11100 582
rect 11164 580 11170 644
rect 11830 580 11836 644
rect 11900 642 11906 644
rect 11973 642 12039 645
rect 11900 640 12039 642
rect 11900 584 11978 640
rect 12034 584 12039 640
rect 11900 582 12039 584
rect 11900 580 11906 582
rect 11973 579 12039 582
rect 12566 580 12572 644
rect 12636 642 12642 644
rect 12709 642 12775 645
rect 12636 640 12775 642
rect 12636 584 12714 640
rect 12770 584 12775 640
rect 12636 582 12775 584
rect 12636 580 12642 582
rect 12709 579 12775 582
rect 13302 580 13308 644
rect 13372 642 13378 644
rect 13445 642 13511 645
rect 13372 640 13511 642
rect 13372 584 13450 640
rect 13506 584 13511 640
rect 13372 582 13511 584
rect 13372 580 13378 582
rect 13445 579 13511 582
rect 16982 580 16988 644
rect 17052 642 17058 644
rect 17125 642 17191 645
rect 17052 640 17191 642
rect 17052 584 17130 640
rect 17186 584 17191 640
rect 17052 582 17191 584
rect 17052 580 17058 582
rect 17125 579 17191 582
rect 17718 580 17724 644
rect 17788 642 17794 644
rect 17861 642 17927 645
rect 17788 640 17927 642
rect 17788 584 17866 640
rect 17922 584 17927 640
rect 17788 582 17927 584
rect 17788 580 17794 582
rect 17861 579 17927 582
rect 18454 580 18460 644
rect 18524 642 18530 644
rect 18597 642 18663 645
rect 18524 640 18663 642
rect 18524 584 18602 640
rect 18658 584 18663 640
rect 18524 582 18663 584
rect 18524 580 18530 582
rect 18597 579 18663 582
rect 23606 580 23612 644
rect 23676 642 23682 644
rect 23933 642 23999 645
rect 23676 640 23999 642
rect 23676 584 23938 640
rect 23994 584 23999 640
rect 23676 582 23999 584
rect 23676 580 23682 582
rect 23933 579 23999 582
rect 28758 580 28764 644
rect 28828 642 28834 644
rect 28993 642 29059 645
rect 28828 640 29059 642
rect 28828 584 28998 640
rect 29054 584 29059 640
rect 28828 582 29059 584
rect 28828 580 28834 582
rect 28993 579 29059 582
rect 30230 580 30236 644
rect 30300 642 30306 644
rect 30373 642 30439 645
rect 30300 640 30439 642
rect 30300 584 30378 640
rect 30434 584 30439 640
rect 30300 582 30439 584
rect 30300 580 30306 582
rect 30373 579 30439 582
rect 35617 644 35683 645
rect 35617 640 35664 644
rect 35728 642 35734 644
rect 36261 642 36327 645
rect 36394 642 36400 644
rect 35617 584 35622 640
rect 35617 580 35664 584
rect 35728 582 35774 642
rect 36261 640 36400 642
rect 36261 584 36266 640
rect 36322 584 36400 640
rect 36261 582 36400 584
rect 35728 580 35734 582
rect 35617 579 35683 580
rect 36261 579 36327 582
rect 36394 580 36400 582
rect 36464 580 36470 644
rect 36905 642 36971 645
rect 37130 642 37136 644
rect 36905 640 37136 642
rect 36905 584 36910 640
rect 36966 584 37136 640
rect 36905 582 37136 584
rect 36905 579 36971 582
rect 37130 580 37136 582
rect 37200 580 37206 644
rect 37866 580 37872 644
rect 37936 642 37942 644
rect 38101 642 38167 645
rect 37936 640 38167 642
rect 37936 584 38106 640
rect 38162 584 38167 640
rect 37936 582 38167 584
rect 37936 580 37942 582
rect 38101 579 38167 582
rect 38561 644 38627 645
rect 38561 640 38608 644
rect 38672 642 38678 644
rect 39941 642 40007 645
rect 40769 644 40835 645
rect 40074 642 40080 644
rect 38561 584 38566 640
rect 38561 580 38608 584
rect 38672 582 38718 642
rect 39941 640 40080 642
rect 39941 584 39946 640
rect 40002 584 40080 640
rect 39941 582 40080 584
rect 38672 580 38678 582
rect 38561 579 38627 580
rect 39941 579 40007 582
rect 40074 580 40080 582
rect 40144 580 40150 644
rect 40769 640 40816 644
rect 40880 642 40886 644
rect 41413 642 41479 645
rect 41546 642 41552 644
rect 40769 584 40774 640
rect 40769 580 40816 584
rect 40880 582 40926 642
rect 41413 640 41552 642
rect 41413 584 41418 640
rect 41474 584 41552 640
rect 41413 582 41552 584
rect 40880 580 40886 582
rect 40769 579 40835 580
rect 41413 579 41479 582
rect 41546 580 41552 582
rect 41616 580 41622 644
rect 42057 642 42123 645
rect 42282 642 42288 644
rect 42057 640 42288 642
rect 42057 584 42062 640
rect 42118 584 42288 640
rect 42057 582 42288 584
rect 42057 579 42123 582
rect 42282 580 42288 582
rect 42352 580 42358 644
rect 43018 580 43024 644
rect 43088 642 43094 644
rect 43253 642 43319 645
rect 43088 640 43319 642
rect 43088 584 43258 640
rect 43314 584 43319 640
rect 43088 582 43319 584
rect 43088 580 43094 582
rect 43253 579 43319 582
rect 43754 580 43760 644
rect 43824 642 43830 644
rect 43989 642 44055 645
rect 43824 640 44055 642
rect 43824 584 43994 640
rect 44050 584 44055 640
rect 43824 582 44055 584
rect 43824 580 43830 582
rect 43989 579 44055 582
rect 44490 580 44496 644
rect 44560 642 44566 644
rect 44633 642 44699 645
rect 44560 640 44699 642
rect 44560 584 44638 640
rect 44694 584 44699 640
rect 44560 582 44699 584
rect 44560 580 44566 582
rect 44633 579 44699 582
rect 45226 580 45232 644
rect 45296 642 45302 644
rect 45461 642 45527 645
rect 45296 640 45527 642
rect 45296 584 45466 640
rect 45522 584 45527 640
rect 45296 582 45527 584
rect 45296 580 45302 582
rect 45461 579 45527 582
rect 45921 644 45987 645
rect 45921 640 45968 644
rect 46032 642 46038 644
rect 46565 642 46631 645
rect 46698 642 46704 644
rect 45921 584 45926 640
rect 45921 580 45968 584
rect 46032 582 46078 642
rect 46565 640 46704 642
rect 46565 584 46570 640
rect 46626 584 46704 640
rect 46565 582 46704 584
rect 46032 580 46038 582
rect 45921 579 45987 580
rect 46565 579 46631 582
rect 46698 580 46704 582
rect 46768 580 46774 644
rect 47209 642 47275 645
rect 47434 642 47440 644
rect 47209 640 47440 642
rect 47209 584 47214 640
rect 47270 584 47440 640
rect 47209 582 47440 584
rect 47209 579 47275 582
rect 47434 580 47440 582
rect 47504 580 47510 644
rect 48170 580 48176 644
rect 48240 642 48246 644
rect 48313 642 48379 645
rect 48240 640 48379 642
rect 48240 584 48318 640
rect 48374 584 48379 640
rect 48240 582 48379 584
rect 48240 580 48246 582
rect 48313 579 48379 582
rect 48906 580 48912 644
rect 48976 642 48982 644
rect 49141 642 49207 645
rect 48976 640 49207 642
rect 48976 584 49146 640
rect 49202 584 49207 640
rect 48976 582 49207 584
rect 48976 580 48982 582
rect 49141 579 49207 582
rect 49642 580 49648 644
rect 49712 642 49718 644
rect 49785 642 49851 645
rect 49712 640 49851 642
rect 49712 584 49790 640
rect 49846 584 49851 640
rect 49712 582 49851 584
rect 49712 580 49718 582
rect 49785 579 49851 582
rect 50378 580 50384 644
rect 50448 642 50454 644
rect 50613 642 50679 645
rect 50448 640 50679 642
rect 50448 584 50618 640
rect 50674 584 50679 640
rect 50448 582 50679 584
rect 50448 580 50454 582
rect 50613 579 50679 582
rect 51073 644 51139 645
rect 51073 640 51120 644
rect 51184 642 51190 644
rect 51717 642 51783 645
rect 51850 642 51856 644
rect 51073 584 51078 640
rect 51073 580 51120 584
rect 51184 582 51230 642
rect 51717 640 51856 642
rect 51717 584 51722 640
rect 51778 584 51856 640
rect 51717 582 51856 584
rect 51184 580 51190 582
rect 51073 579 51139 580
rect 51717 579 51783 582
rect 51850 580 51856 582
rect 51920 580 51926 644
rect 52361 642 52427 645
rect 53373 644 53439 645
rect 54845 644 54911 645
rect 52586 642 52592 644
rect 52361 640 52592 642
rect 52361 584 52366 640
rect 52422 584 52592 640
rect 52361 582 52592 584
rect 52361 579 52427 582
rect 52586 580 52592 582
rect 52656 580 52662 644
rect 53322 642 53328 644
rect 53282 582 53328 642
rect 53392 640 53439 644
rect 54794 642 54800 644
rect 53434 584 53439 640
rect 53322 580 53328 582
rect 53392 580 53439 584
rect 54754 582 54800 642
rect 54864 640 54911 644
rect 54906 584 54911 640
rect 54794 580 54800 582
rect 54864 580 54911 584
rect 55530 580 55536 644
rect 55600 642 55606 644
rect 55673 642 55739 645
rect 55600 640 55739 642
rect 55600 584 55678 640
rect 55734 584 55739 640
rect 55600 582 55739 584
rect 55600 580 55606 582
rect 53373 579 53439 580
rect 54845 579 54911 580
rect 55673 579 55739 582
rect 56225 644 56291 645
rect 57053 644 57119 645
rect 57789 644 57855 645
rect 56225 640 56272 644
rect 56336 642 56342 644
rect 57002 642 57008 644
rect 56225 584 56230 640
rect 56225 580 56272 584
rect 56336 582 56382 642
rect 56962 582 57008 642
rect 57072 640 57119 644
rect 57738 642 57744 644
rect 57114 584 57119 640
rect 56336 580 56342 582
rect 57002 580 57008 582
rect 57072 580 57119 584
rect 57698 582 57744 642
rect 57808 640 57855 644
rect 57850 584 57855 640
rect 57738 580 57744 582
rect 57808 580 57855 584
rect 58474 580 58480 644
rect 58544 642 58550 644
rect 58617 642 58683 645
rect 58544 640 58683 642
rect 58544 584 58622 640
rect 58678 584 58683 640
rect 58544 582 58683 584
rect 58544 580 58550 582
rect 56225 579 56291 580
rect 57053 579 57119 580
rect 57789 579 57855 580
rect 58617 579 58683 582
rect 60682 580 60688 644
rect 60752 642 60758 644
rect 60825 642 60891 645
rect 60752 640 60891 642
rect 60752 584 60830 640
rect 60886 584 60891 640
rect 60752 582 60891 584
rect 60752 580 60758 582
rect 60825 579 60891 582
rect 61418 580 61424 644
rect 61488 642 61494 644
rect 61561 642 61627 645
rect 61488 640 61627 642
rect 61488 584 61566 640
rect 61622 584 61627 640
rect 61488 582 61627 584
rect 61488 580 61494 582
rect 61561 579 61627 582
rect 62154 580 62160 644
rect 62224 642 62230 644
rect 62297 642 62363 645
rect 62941 644 63007 645
rect 62890 642 62896 644
rect 62224 640 62363 642
rect 62224 584 62302 640
rect 62358 584 62363 640
rect 62224 582 62363 584
rect 62850 582 62896 642
rect 62960 640 63007 644
rect 63002 584 63007 640
rect 62224 580 62230 582
rect 62297 579 62363 582
rect 62890 580 62896 582
rect 62960 580 63007 584
rect 63626 580 63632 644
rect 63696 642 63702 644
rect 63769 642 63835 645
rect 63696 640 63835 642
rect 63696 584 63774 640
rect 63830 584 63835 640
rect 63696 582 63835 584
rect 63696 580 63702 582
rect 62941 579 63007 580
rect 63769 579 63835 582
rect 64362 580 64368 644
rect 64432 642 64438 644
rect 64505 642 64571 645
rect 64432 640 64571 642
rect 64432 584 64510 640
rect 64566 584 64571 640
rect 64432 582 64571 584
rect 64432 580 64438 582
rect 64505 579 64571 582
rect 65098 580 65104 644
rect 65168 642 65174 644
rect 65609 642 65675 645
rect 65168 640 65675 642
rect 65168 584 65614 640
rect 65670 584 65675 640
rect 65168 582 65675 584
rect 65168 580 65174 582
rect 65609 579 65675 582
rect 72141 642 72207 645
rect 72734 642 72740 644
rect 72141 640 72740 642
rect 72141 584 72146 640
rect 72202 584 72740 640
rect 72141 582 72740 584
rect 72141 579 72207 582
rect 72734 580 72740 582
rect 72804 580 72810 644
rect 74717 642 74783 645
rect 74942 642 74948 644
rect 74717 640 74948 642
rect 74717 584 74722 640
rect 74778 584 74948 640
rect 74717 582 74948 584
rect 74717 579 74783 582
rect 74942 580 74948 582
rect 75012 580 75018 644
rect 82721 642 82787 645
rect 113406 642 113466 718
rect 117589 715 117655 718
rect 138790 716 138796 718
rect 138860 716 138907 720
rect 140998 716 141004 780
rect 141068 778 141074 780
rect 141969 778 142035 781
rect 141068 776 142035 778
rect 141068 720 141974 776
rect 142030 720 142035 776
rect 141068 718 142035 720
rect 141068 716 141074 718
rect 138841 715 138907 716
rect 141969 715 142035 718
rect 143206 716 143212 780
rect 143276 778 143282 780
rect 143533 778 143599 781
rect 143276 776 143599 778
rect 143276 720 143538 776
rect 143594 720 143599 776
rect 143276 718 143599 720
rect 143276 716 143282 718
rect 143533 715 143599 718
rect 143942 716 143948 780
rect 144012 778 144018 780
rect 144545 778 144611 781
rect 144012 776 144611 778
rect 144012 720 144550 776
rect 144606 720 144611 776
rect 144012 718 144611 720
rect 144012 716 144018 718
rect 144545 715 144611 718
rect 145414 716 145420 780
rect 145484 778 145490 780
rect 145833 778 145899 781
rect 146201 780 146267 781
rect 146150 778 146156 780
rect 145484 776 145899 778
rect 145484 720 145838 776
rect 145894 720 145899 776
rect 145484 718 145899 720
rect 146110 718 146156 778
rect 146220 776 146267 780
rect 146262 720 146267 776
rect 145484 716 145490 718
rect 145833 715 145899 718
rect 146150 716 146156 718
rect 146220 716 146267 720
rect 146886 716 146892 780
rect 146956 778 146962 780
rect 147121 778 147187 781
rect 146956 776 147187 778
rect 146956 720 147126 776
rect 147182 720 147187 776
rect 146956 718 147187 720
rect 146956 716 146962 718
rect 146201 715 146267 716
rect 147121 715 147187 718
rect 148358 716 148364 780
rect 148428 778 148434 780
rect 148501 778 148567 781
rect 148428 776 148567 778
rect 148428 720 148506 776
rect 148562 720 148567 776
rect 148428 718 148567 720
rect 148428 716 148434 718
rect 148501 715 148567 718
rect 149094 716 149100 780
rect 149164 778 149170 780
rect 149697 778 149763 781
rect 149164 776 149763 778
rect 149164 720 149702 776
rect 149758 720 149763 776
rect 149164 718 149763 720
rect 149164 716 149170 718
rect 149697 715 149763 718
rect 150566 716 150572 780
rect 150636 778 150642 780
rect 150985 778 151051 781
rect 150636 776 151051 778
rect 150636 720 150990 776
rect 151046 720 151051 776
rect 150636 718 151051 720
rect 150636 716 150642 718
rect 150985 715 151051 718
rect 151302 716 151308 780
rect 151372 778 151378 780
rect 151629 778 151695 781
rect 151372 776 151695 778
rect 151372 720 151634 776
rect 151690 720 151695 776
rect 151372 718 151695 720
rect 151372 716 151378 718
rect 151629 715 151695 718
rect 152038 716 152044 780
rect 152108 778 152114 780
rect 152273 778 152339 781
rect 152108 776 152339 778
rect 152108 720 152278 776
rect 152334 720 152339 776
rect 152108 718 152339 720
rect 152108 716 152114 718
rect 152273 715 152339 718
rect 152774 716 152780 780
rect 152844 778 152850 780
rect 153193 778 153259 781
rect 152844 776 153259 778
rect 152844 720 153198 776
rect 153254 720 153259 776
rect 152844 718 153259 720
rect 152844 716 152850 718
rect 153193 715 153259 718
rect 154246 716 154252 780
rect 154316 778 154322 780
rect 154573 778 154639 781
rect 154316 776 154639 778
rect 154316 720 154578 776
rect 154634 720 154639 776
rect 154316 718 154639 720
rect 154316 716 154322 718
rect 154573 715 154639 718
rect 156781 778 156847 781
rect 169293 778 169359 781
rect 248370 778 248430 854
rect 258073 851 258139 854
rect 257889 778 257955 781
rect 156781 776 169218 778
rect 156781 720 156786 776
rect 156842 720 169218 776
rect 156781 718 169218 720
rect 156781 715 156847 718
rect 82721 640 113466 642
rect 82721 584 82726 640
rect 82782 584 113466 640
rect 82721 582 113466 584
rect 114185 644 114251 645
rect 114185 640 114232 644
rect 114296 642 114302 644
rect 114185 584 114190 640
rect 82721 579 82787 582
rect 114185 580 114232 584
rect 114296 582 114342 642
rect 114296 580 114302 582
rect 114962 580 114968 644
rect 115032 642 115038 644
rect 115197 642 115263 645
rect 115749 644 115815 645
rect 115698 642 115704 644
rect 115032 640 115263 642
rect 115032 584 115202 640
rect 115258 584 115263 640
rect 115032 582 115263 584
rect 115658 582 115704 642
rect 115768 640 115815 644
rect 115810 584 115815 640
rect 115032 580 115038 582
rect 114185 579 114251 580
rect 115197 579 115263 582
rect 115698 580 115704 582
rect 115768 580 115815 584
rect 116434 580 116440 644
rect 116504 642 116510 644
rect 116669 642 116735 645
rect 116504 640 116735 642
rect 116504 584 116674 640
rect 116730 584 116735 640
rect 116504 582 116735 584
rect 116504 580 116510 582
rect 115749 579 115815 580
rect 116669 579 116735 582
rect 117906 580 117912 644
rect 117976 642 117982 644
rect 118049 642 118115 645
rect 118693 644 118759 645
rect 118642 642 118648 644
rect 117976 640 118115 642
rect 117976 584 118054 640
rect 118110 584 118115 640
rect 117976 582 118115 584
rect 118602 582 118648 642
rect 118712 640 118759 644
rect 118754 584 118759 640
rect 117976 580 117982 582
rect 118049 579 118115 582
rect 118642 580 118648 582
rect 118712 580 118759 584
rect 118693 579 118759 580
rect 119337 644 119403 645
rect 119337 640 119384 644
rect 119448 642 119454 644
rect 119337 584 119342 640
rect 119337 580 119384 584
rect 119448 582 119494 642
rect 119448 580 119454 582
rect 120114 580 120120 644
rect 120184 642 120190 644
rect 120349 642 120415 645
rect 120184 640 120415 642
rect 120184 584 120354 640
rect 120410 584 120415 640
rect 120184 582 120415 584
rect 120184 580 120190 582
rect 119337 579 119403 580
rect 120349 579 120415 582
rect 120850 580 120856 644
rect 120920 642 120926 644
rect 121085 642 121151 645
rect 120920 640 121151 642
rect 120920 584 121090 640
rect 121146 584 121151 640
rect 120920 582 121151 584
rect 120920 580 120926 582
rect 121085 579 121151 582
rect 121586 580 121592 644
rect 121656 642 121662 644
rect 121821 642 121887 645
rect 121656 640 121887 642
rect 121656 584 121826 640
rect 121882 584 121887 640
rect 121656 582 121887 584
rect 121656 580 121662 582
rect 121821 579 121887 582
rect 122322 580 122328 644
rect 122392 642 122398 644
rect 122649 642 122715 645
rect 123109 644 123175 645
rect 123058 642 123064 644
rect 122392 640 122715 642
rect 122392 584 122654 640
rect 122710 584 122715 640
rect 122392 582 122715 584
rect 123018 582 123064 642
rect 123128 640 123175 644
rect 123170 584 123175 640
rect 122392 580 122398 582
rect 122649 579 122715 582
rect 123058 580 123064 582
rect 123128 580 123175 584
rect 123794 580 123800 644
rect 123864 642 123870 644
rect 123937 642 124003 645
rect 123864 640 124003 642
rect 123864 584 123942 640
rect 123998 584 124003 640
rect 123864 582 124003 584
rect 123864 580 123870 582
rect 123109 579 123175 580
rect 123937 579 124003 582
rect 124530 580 124536 644
rect 124600 642 124606 644
rect 124765 642 124831 645
rect 125317 644 125383 645
rect 125266 642 125272 644
rect 124600 640 124831 642
rect 124600 584 124770 640
rect 124826 584 124831 640
rect 124600 582 124831 584
rect 125226 582 125272 642
rect 125336 640 125383 644
rect 125378 584 125383 640
rect 124600 580 124606 582
rect 124765 579 124831 582
rect 125266 580 125272 582
rect 125336 580 125383 584
rect 126002 580 126008 644
rect 126072 642 126078 644
rect 126329 642 126395 645
rect 126789 644 126855 645
rect 126738 642 126744 644
rect 126072 640 126395 642
rect 126072 584 126334 640
rect 126390 584 126395 640
rect 126072 582 126395 584
rect 126698 582 126744 642
rect 126808 640 126855 644
rect 126850 584 126855 640
rect 126072 580 126078 582
rect 125317 579 125383 580
rect 126329 579 126395 582
rect 126738 580 126744 582
rect 126808 580 126855 584
rect 127474 580 127480 644
rect 127544 642 127550 644
rect 127801 642 127867 645
rect 127544 640 127867 642
rect 127544 584 127806 640
rect 127862 584 127867 640
rect 127544 582 127867 584
rect 127544 580 127550 582
rect 126789 579 126855 580
rect 127801 579 127867 582
rect 128946 580 128952 644
rect 129016 642 129022 644
rect 129273 642 129339 645
rect 129016 640 129339 642
rect 129016 584 129278 640
rect 129334 584 129339 640
rect 129016 582 129339 584
rect 129016 580 129022 582
rect 129273 579 129339 582
rect 129682 580 129688 644
rect 129752 642 129758 644
rect 130009 642 130075 645
rect 129752 640 130075 642
rect 129752 584 130014 640
rect 130070 584 130075 640
rect 129752 582 130075 584
rect 129752 580 129758 582
rect 130009 579 130075 582
rect 131154 580 131160 644
rect 131224 642 131230 644
rect 131573 642 131639 645
rect 131224 640 131639 642
rect 131224 584 131578 640
rect 131634 584 131639 640
rect 131224 582 131639 584
rect 131224 580 131230 582
rect 131573 579 131639 582
rect 131890 580 131896 644
rect 131960 642 131966 644
rect 132125 642 132191 645
rect 131960 640 132191 642
rect 131960 584 132130 640
rect 132186 584 132191 640
rect 131960 582 132191 584
rect 131960 580 131966 582
rect 132125 579 132191 582
rect 132626 580 132632 644
rect 132696 642 132702 644
rect 132953 642 133019 645
rect 132696 640 133019 642
rect 132696 584 132958 640
rect 133014 584 133019 640
rect 132696 582 133019 584
rect 132696 580 132702 582
rect 132953 579 133019 582
rect 133362 580 133368 644
rect 133432 642 133438 644
rect 133689 642 133755 645
rect 133432 640 133755 642
rect 133432 584 133694 640
rect 133750 584 133755 640
rect 133432 582 133755 584
rect 133432 580 133438 582
rect 133689 579 133755 582
rect 134098 580 134104 644
rect 134168 642 134174 644
rect 134425 642 134491 645
rect 134168 640 134491 642
rect 134168 584 134430 640
rect 134486 584 134491 640
rect 134168 582 134491 584
rect 134168 580 134174 582
rect 134425 579 134491 582
rect 138054 580 138060 644
rect 138124 642 138130 644
rect 138749 642 138815 645
rect 138124 640 138815 642
rect 138124 584 138754 640
rect 138810 584 138815 640
rect 138124 582 138815 584
rect 138124 580 138130 582
rect 138749 579 138815 582
rect 141734 580 141740 644
rect 141804 642 141810 644
rect 142061 642 142127 645
rect 141804 640 142127 642
rect 141804 584 142066 640
rect 142122 584 142127 640
rect 141804 582 142127 584
rect 141804 580 141810 582
rect 142061 579 142127 582
rect 147622 580 147628 644
rect 147692 642 147698 644
rect 148409 642 148475 645
rect 147692 640 148475 642
rect 147692 584 148414 640
rect 148470 584 148475 640
rect 147692 582 148475 584
rect 147692 580 147698 582
rect 148409 579 148475 582
rect 153510 580 153516 644
rect 153580 642 153586 644
rect 154205 642 154271 645
rect 153580 640 154271 642
rect 153580 584 154210 640
rect 154266 584 154271 640
rect 153580 582 154271 584
rect 153580 580 153586 582
rect 154205 579 154271 582
rect 158662 580 158668 644
rect 158732 642 158738 644
rect 158805 642 158871 645
rect 158732 640 158871 642
rect 158732 584 158810 640
rect 158866 584 158871 640
rect 158732 582 158871 584
rect 158732 580 158738 582
rect 158805 579 158871 582
rect 160870 580 160876 644
rect 160940 642 160946 644
rect 161289 642 161355 645
rect 160940 640 161355 642
rect 160940 584 161294 640
rect 161350 584 161355 640
rect 160940 582 161355 584
rect 160940 580 160946 582
rect 161289 579 161355 582
rect 162342 580 162348 644
rect 162412 642 162418 644
rect 162485 642 162551 645
rect 162412 640 162551 642
rect 162412 584 162490 640
rect 162546 584 162551 640
rect 162412 582 162551 584
rect 162412 580 162418 582
rect 162485 579 162551 582
rect 164550 580 164556 644
rect 164620 642 164626 644
rect 164693 642 164759 645
rect 164620 640 164759 642
rect 164620 584 164698 640
rect 164754 584 164759 640
rect 164620 582 164759 584
rect 164620 580 164626 582
rect 164693 579 164759 582
rect 167494 580 167500 644
rect 167564 642 167570 644
rect 168005 642 168071 645
rect 169017 644 169083 645
rect 168966 642 168972 644
rect 167564 640 168071 642
rect 167564 584 168010 640
rect 168066 584 168071 640
rect 167564 582 168071 584
rect 168926 582 168972 642
rect 169036 640 169083 644
rect 169078 584 169083 640
rect 167564 580 167570 582
rect 168005 579 168071 582
rect 168966 580 168972 582
rect 169036 580 169083 584
rect 169158 642 169218 718
rect 169293 776 248430 778
rect 169293 720 169298 776
rect 169354 720 248430 776
rect 169293 718 248430 720
rect 249750 776 257955 778
rect 249750 720 257894 776
rect 257950 720 257955 776
rect 249750 718 257955 720
rect 169293 715 169359 718
rect 249750 642 249810 718
rect 257889 715 257955 718
rect 169158 582 249810 642
rect 250018 580 250024 644
rect 250088 642 250094 644
rect 250161 642 250227 645
rect 251541 644 251607 645
rect 252277 644 252343 645
rect 251490 642 251496 644
rect 250088 640 250227 642
rect 250088 584 250166 640
rect 250222 584 250227 640
rect 250088 582 250227 584
rect 251450 582 251496 642
rect 251560 640 251607 644
rect 252226 642 252232 644
rect 251602 584 251607 640
rect 250088 580 250094 582
rect 169017 579 169083 580
rect 250161 579 250227 582
rect 251490 580 251496 582
rect 251560 580 251607 584
rect 252186 582 252232 642
rect 252296 640 252343 644
rect 252338 584 252343 640
rect 252226 580 252232 582
rect 252296 580 252343 584
rect 252962 580 252968 644
rect 253032 642 253038 644
rect 253473 642 253539 645
rect 253032 640 253539 642
rect 253032 584 253478 640
rect 253534 584 253539 640
rect 253032 582 253539 584
rect 253032 580 253038 582
rect 251541 579 251607 580
rect 252277 579 252343 580
rect 253473 579 253539 582
rect 253698 580 253704 644
rect 253768 642 253774 644
rect 253841 642 253907 645
rect 255221 644 255287 645
rect 255170 642 255176 644
rect 253768 640 253907 642
rect 253768 584 253846 640
rect 253902 584 253907 640
rect 253768 582 253907 584
rect 255130 582 255176 642
rect 255240 640 255287 644
rect 255282 584 255287 640
rect 253768 580 253774 582
rect 253841 579 253907 582
rect 255170 580 255176 582
rect 255240 580 255287 584
rect 255906 580 255912 644
rect 255976 642 255982 644
rect 256417 642 256483 645
rect 256693 644 256759 645
rect 257429 644 257495 645
rect 256642 642 256648 644
rect 255976 640 256483 642
rect 255976 584 256422 640
rect 256478 584 256483 640
rect 255976 582 256483 584
rect 256602 582 256648 642
rect 256712 640 256759 644
rect 257378 642 257384 644
rect 256754 584 256759 640
rect 255976 580 255982 582
rect 255221 579 255287 580
rect 256417 579 256483 582
rect 256642 580 256648 582
rect 256712 580 256759 584
rect 257338 582 257384 642
rect 257448 640 257495 644
rect 257490 584 257495 640
rect 257378 580 257384 582
rect 257448 580 257495 584
rect 258850 580 258856 644
rect 258920 642 258926 644
rect 259177 642 259243 645
rect 258920 640 259243 642
rect 258920 584 259182 640
rect 259238 584 259243 640
rect 258920 582 259243 584
rect 258920 580 258926 582
rect 256693 579 256759 580
rect 257429 579 257495 580
rect 259177 579 259243 582
rect 259586 580 259592 644
rect 259656 642 259662 644
rect 259913 642 259979 645
rect 259656 640 259979 642
rect 259656 584 259918 640
rect 259974 584 259979 640
rect 259656 582 259979 584
rect 259656 580 259662 582
rect 259913 579 259979 582
rect 260322 580 260328 644
rect 260392 642 260398 644
rect 260465 642 260531 645
rect 260392 640 260531 642
rect 260392 584 260470 640
rect 260526 584 260531 640
rect 260392 582 260531 584
rect 260392 580 260398 582
rect 260465 579 260531 582
rect 261058 580 261064 644
rect 261128 642 261134 644
rect 261753 642 261819 645
rect 261128 640 261819 642
rect 261128 584 261758 640
rect 261814 584 261819 640
rect 261128 582 261819 584
rect 261128 580 261134 582
rect 261753 579 261819 582
rect 262489 644 262555 645
rect 263225 644 263291 645
rect 262489 640 262536 644
rect 262600 642 262606 644
rect 262489 584 262494 640
rect 262489 580 262536 584
rect 262600 582 262646 642
rect 263225 640 263272 644
rect 263336 642 263342 644
rect 263225 584 263230 640
rect 262600 580 262606 582
rect 263225 580 263272 584
rect 263336 582 263382 642
rect 263336 580 263342 582
rect 264002 580 264008 644
rect 264072 642 264078 644
rect 264329 642 264395 645
rect 264072 640 264395 642
rect 264072 584 264334 640
rect 264390 584 264395 640
rect 264072 582 264395 584
rect 264072 580 264078 582
rect 262489 579 262555 580
rect 263225 579 263291 580
rect 264329 579 264395 582
rect 265341 642 265407 645
rect 265474 642 265480 644
rect 265341 640 265480 642
rect 265341 584 265346 640
rect 265402 584 265480 640
rect 265341 582 265480 584
rect 265341 579 265407 582
rect 265474 580 265480 582
rect 265544 580 265550 644
rect 266077 642 266143 645
rect 266905 644 266971 645
rect 267641 644 267707 645
rect 268377 644 268443 645
rect 266210 642 266216 644
rect 266077 640 266216 642
rect 266077 584 266082 640
rect 266138 584 266216 640
rect 266077 582 266216 584
rect 266077 579 266143 582
rect 266210 580 266216 582
rect 266280 580 266286 644
rect 266905 640 266952 644
rect 267016 642 267022 644
rect 266905 584 266910 640
rect 266905 580 266952 584
rect 267016 582 267062 642
rect 267641 640 267688 644
rect 267752 642 267758 644
rect 267641 584 267646 640
rect 267016 580 267022 582
rect 267641 580 267688 584
rect 267752 582 267794 642
rect 268377 640 268424 644
rect 268488 642 268494 644
rect 268377 584 268382 640
rect 267752 580 267758 582
rect 268377 580 268424 584
rect 268488 582 268534 642
rect 268488 580 268494 582
rect 266905 579 266971 580
rect 267641 579 267707 580
rect 268377 579 268443 580
rect 28022 444 28028 508
rect 28092 506 28098 508
rect 28717 506 28783 509
rect 28092 504 28783 506
rect 28092 448 28722 504
rect 28778 448 28783 504
rect 28092 446 28783 448
rect 28092 444 28098 446
rect 28717 443 28783 446
rect 29494 444 29500 508
rect 29564 506 29570 508
rect 29913 506 29979 509
rect 29564 504 29979 506
rect 29564 448 29918 504
rect 29974 448 29979 504
rect 29564 446 29979 448
rect 29564 444 29570 446
rect 29913 443 29979 446
rect 31702 444 31708 508
rect 31772 506 31778 508
rect 32489 506 32555 509
rect 31772 504 32555 506
rect 31772 448 32494 504
rect 32550 448 32555 504
rect 31772 446 32555 448
rect 31772 444 31778 446
rect 32489 443 32555 446
rect 65834 444 65840 508
rect 65904 506 65910 508
rect 66161 506 66227 509
rect 65904 504 66227 506
rect 65904 448 66166 504
rect 66222 448 66227 504
rect 65904 446 66227 448
rect 65904 444 65910 446
rect 66161 443 66227 446
rect 66570 444 66576 508
rect 66640 506 66646 508
rect 67541 506 67607 509
rect 66640 504 67607 506
rect 66640 448 67546 504
rect 67602 448 67607 504
rect 66640 446 67607 448
rect 66640 444 66646 446
rect 67541 443 67607 446
rect 83917 506 83983 509
rect 96521 506 96587 509
rect 100017 508 100083 509
rect 103237 508 103303 509
rect 97022 506 97028 508
rect 83917 504 94514 506
rect 83917 448 83922 504
rect 83978 448 94514 504
rect 83917 446 94514 448
rect 83917 443 83983 446
rect 30966 308 30972 372
rect 31036 370 31042 372
rect 31569 370 31635 373
rect 31036 368 31635 370
rect 31036 312 31574 368
rect 31630 312 31635 368
rect 31036 310 31635 312
rect 31036 308 31042 310
rect 31569 307 31635 310
rect 34421 370 34487 373
rect 34922 370 34928 372
rect 34421 368 34928 370
rect 34421 312 34426 368
rect 34482 312 34928 368
rect 34421 310 34928 312
rect 34421 307 34487 310
rect 34922 308 34928 310
rect 34992 308 34998 372
rect 38837 370 38903 373
rect 39338 370 39344 372
rect 38837 368 39344 370
rect 38837 312 38842 368
rect 38898 312 39344 368
rect 38837 310 39344 312
rect 38837 307 38903 310
rect 39338 308 39344 310
rect 39408 308 39414 372
rect 89662 308 89668 372
rect 89732 370 89738 372
rect 90817 370 90883 373
rect 89732 368 90883 370
rect 89732 312 90822 368
rect 90878 312 90883 368
rect 89732 310 90883 312
rect 89732 308 89738 310
rect 90817 307 90883 310
rect 91134 308 91140 372
rect 91204 370 91210 372
rect 91737 370 91803 373
rect 91204 368 91803 370
rect 91204 312 91742 368
rect 91798 312 91803 368
rect 91204 310 91803 312
rect 91204 308 91210 310
rect 91737 307 91803 310
rect 92606 308 92612 372
rect 92676 370 92682 372
rect 93025 370 93091 373
rect 92676 368 93091 370
rect 92676 312 93030 368
rect 93086 312 93091 368
rect 92676 310 93091 312
rect 94454 370 94514 446
rect 96521 504 97028 506
rect 96521 448 96526 504
rect 96582 448 97028 504
rect 96521 446 97028 448
rect 96521 443 96587 446
rect 97022 444 97028 446
rect 97092 444 97098 508
rect 99966 506 99972 508
rect 99926 446 99972 506
rect 100036 504 100083 508
rect 103186 506 103192 508
rect 100078 448 100083 504
rect 99966 444 99972 446
rect 100036 444 100083 448
rect 103146 446 103192 506
rect 103256 504 103303 508
rect 103298 448 103303 504
rect 103186 444 103192 446
rect 103256 444 103303 448
rect 100017 443 100083 444
rect 103237 443 103303 444
rect 103881 508 103947 509
rect 104709 508 104775 509
rect 103881 504 103928 508
rect 103992 506 103998 508
rect 104658 506 104664 508
rect 103881 448 103886 504
rect 103881 444 103928 448
rect 103992 446 104038 506
rect 104618 446 104664 506
rect 104728 504 104775 508
rect 104770 448 104775 504
rect 103992 444 103998 446
rect 104658 444 104664 446
rect 104728 444 104775 448
rect 105394 444 105400 508
rect 105464 506 105470 508
rect 105629 506 105695 509
rect 106181 508 106247 509
rect 106130 506 106136 508
rect 105464 504 105695 506
rect 105464 448 105634 504
rect 105690 448 105695 504
rect 105464 446 105695 448
rect 106090 446 106136 506
rect 106200 504 106247 508
rect 106242 448 106247 504
rect 105464 444 105470 446
rect 103881 443 103947 444
rect 104709 443 104775 444
rect 105629 443 105695 446
rect 106130 444 106136 446
rect 106200 444 106247 448
rect 106866 444 106872 508
rect 106936 506 106942 508
rect 107101 506 107167 509
rect 106936 504 107167 506
rect 106936 448 107106 504
rect 107162 448 107167 504
rect 106936 446 107167 448
rect 106936 444 106942 446
rect 106181 443 106247 444
rect 107101 443 107167 446
rect 107602 444 107608 508
rect 107672 506 107678 508
rect 107745 506 107811 509
rect 108389 508 108455 509
rect 108338 506 108344 508
rect 107672 504 107811 506
rect 107672 448 107750 504
rect 107806 448 107811 504
rect 107672 446 107811 448
rect 108298 446 108344 506
rect 108408 504 108455 508
rect 108450 448 108455 504
rect 107672 444 107678 446
rect 107745 443 107811 446
rect 108338 444 108344 446
rect 108408 444 108455 448
rect 108389 443 108455 444
rect 109033 508 109099 509
rect 109033 504 109080 508
rect 109144 506 109150 508
rect 109033 448 109038 504
rect 109033 444 109080 448
rect 109144 446 109190 506
rect 109144 444 109150 446
rect 109810 444 109816 508
rect 109880 506 109886 508
rect 110045 506 110111 509
rect 109880 504 110111 506
rect 109880 448 110050 504
rect 110106 448 110111 504
rect 109880 446 110111 448
rect 109880 444 109886 446
rect 109033 443 109099 444
rect 110045 443 110111 446
rect 110546 444 110552 508
rect 110616 506 110622 508
rect 110781 506 110847 509
rect 110616 504 110847 506
rect 110616 448 110786 504
rect 110842 448 110847 504
rect 110616 446 110847 448
rect 110616 444 110622 446
rect 110781 443 110847 446
rect 111282 444 111288 508
rect 111352 506 111358 508
rect 111517 506 111583 509
rect 111352 504 111583 506
rect 111352 448 111522 504
rect 111578 448 111583 504
rect 111352 446 111583 448
rect 111352 444 111358 446
rect 111517 443 111583 446
rect 112018 444 112024 508
rect 112088 506 112094 508
rect 112253 506 112319 509
rect 112088 504 112319 506
rect 112088 448 112258 504
rect 112314 448 112319 504
rect 112088 446 112319 448
rect 112088 444 112094 446
rect 112253 443 112319 446
rect 112754 444 112760 508
rect 112824 506 112830 508
rect 112897 506 112963 509
rect 120441 506 120507 509
rect 112824 504 112963 506
rect 112824 448 112902 504
rect 112958 448 112963 504
rect 112824 446 112963 448
rect 112824 444 112830 446
rect 112897 443 112963 446
rect 113130 504 120507 506
rect 113130 448 120446 504
rect 120502 448 120507 504
rect 113130 446 120507 448
rect 98729 370 98795 373
rect 94454 368 98795 370
rect 94454 312 98734 368
rect 98790 312 98795 368
rect 94454 310 98795 312
rect 92676 308 92682 310
rect 93025 307 93091 310
rect 98729 307 98795 310
rect 87045 234 87111 237
rect 113130 234 113190 446
rect 120441 443 120507 446
rect 124029 506 124095 509
rect 124029 504 132510 506
rect 124029 448 124034 504
rect 124090 448 132510 504
rect 124029 446 132510 448
rect 124029 443 124095 446
rect 113541 372 113607 373
rect 113490 370 113496 372
rect 113450 310 113496 370
rect 113560 368 113607 372
rect 113602 312 113607 368
rect 113490 308 113496 310
rect 113560 308 113607 312
rect 130418 308 130424 372
rect 130488 370 130494 372
rect 130837 370 130903 373
rect 130488 368 130903 370
rect 130488 312 130842 368
rect 130898 312 130903 368
rect 130488 310 130903 312
rect 132450 370 132510 446
rect 139526 444 139532 508
rect 139596 506 139602 508
rect 140681 506 140747 509
rect 139596 504 140747 506
rect 139596 448 140686 504
rect 140742 448 140747 504
rect 139596 446 140747 448
rect 139596 444 139602 446
rect 140681 443 140747 446
rect 158621 506 158687 509
rect 234613 506 234679 509
rect 158621 504 234679 506
rect 158621 448 158626 504
rect 158682 448 234618 504
rect 234674 448 234679 504
rect 158621 446 234679 448
rect 158621 443 158687 446
rect 234613 443 234679 446
rect 234889 506 234955 509
rect 241237 508 241303 509
rect 241973 508 242039 509
rect 243445 508 243511 509
rect 244917 508 244983 509
rect 235022 506 235028 508
rect 234889 504 235028 506
rect 234889 448 234894 504
rect 234950 448 235028 504
rect 234889 446 235028 448
rect 234889 443 234955 446
rect 235022 444 235028 446
rect 235092 444 235098 508
rect 241186 506 241192 508
rect 241146 446 241192 506
rect 241256 504 241303 508
rect 241922 506 241928 508
rect 241298 448 241303 504
rect 241186 444 241192 446
rect 241256 444 241303 448
rect 241882 446 241928 506
rect 241992 504 242039 508
rect 243394 506 243400 508
rect 242034 448 242039 504
rect 241922 444 241928 446
rect 241992 444 242039 448
rect 243354 446 243400 506
rect 243464 504 243511 508
rect 244866 506 244872 508
rect 243506 448 243511 504
rect 243394 444 243400 446
rect 243464 444 243511 448
rect 244826 446 244872 506
rect 244936 504 244983 508
rect 244978 448 244983 504
rect 244866 444 244872 446
rect 244936 444 244983 448
rect 245602 444 245608 508
rect 245672 506 245678 508
rect 246113 506 246179 509
rect 246389 508 246455 509
rect 246338 506 246344 508
rect 245672 504 246179 506
rect 245672 448 246118 504
rect 246174 448 246179 504
rect 245672 446 246179 448
rect 246298 446 246344 506
rect 246408 504 246455 508
rect 246450 448 246455 504
rect 245672 444 245678 446
rect 241237 443 241303 444
rect 241973 443 242039 444
rect 243445 443 243511 444
rect 244917 443 244983 444
rect 246113 443 246179 446
rect 246338 444 246344 446
rect 246408 444 246455 448
rect 246389 443 246455 444
rect 248321 506 248387 509
rect 261845 508 261911 509
rect 248546 506 248552 508
rect 248321 504 248552 506
rect 248321 448 248326 504
rect 248382 448 248552 504
rect 248321 446 248552 448
rect 248321 443 248387 446
rect 248546 444 248552 446
rect 248616 444 248622 508
rect 261794 506 261800 508
rect 261754 446 261800 506
rect 261864 504 261911 508
rect 268886 506 268946 1262
rect 271781 1186 271847 1189
rect 271781 1184 272504 1186
rect 271781 1128 271786 1184
rect 271842 1128 272504 1184
rect 271781 1126 272504 1128
rect 271781 1123 271847 1126
rect 271333 1120 271649 1121
rect 271333 1056 271339 1120
rect 271403 1056 271419 1120
rect 271483 1056 271499 1120
rect 271563 1056 271579 1120
rect 271643 1056 271649 1120
rect 271333 1055 271649 1056
rect 271830 990 272504 1050
rect 269021 914 269087 917
rect 271830 914 271890 990
rect 269021 912 271890 914
rect 269021 856 269026 912
rect 269082 856 271890 912
rect 269021 854 271890 856
rect 269021 851 269087 854
rect 269890 580 269896 644
rect 269960 642 269966 644
rect 270309 642 270375 645
rect 269960 640 270375 642
rect 269960 584 270314 640
rect 270370 584 270375 640
rect 269960 582 270375 584
rect 269960 580 269966 582
rect 270309 579 270375 582
rect 261906 448 261911 504
rect 261794 444 261800 446
rect 261864 444 261911 448
rect 261845 443 261911 444
rect 267690 446 268946 506
rect 160093 370 160159 373
rect 132450 368 160159 370
rect 132450 312 160098 368
rect 160154 312 160159 368
rect 132450 310 160159 312
rect 130488 308 130494 310
rect 113541 307 113607 308
rect 130837 307 130903 310
rect 160093 307 160159 310
rect 163313 370 163379 373
rect 218881 372 218947 373
rect 219617 372 219683 373
rect 218830 370 218836 372
rect 163313 368 215310 370
rect 163313 312 163318 368
rect 163374 312 215310 368
rect 163313 310 215310 312
rect 218790 310 218836 370
rect 218900 368 218947 372
rect 219566 370 219572 372
rect 218942 312 218947 368
rect 163313 307 163379 310
rect 87045 232 113190 234
rect 87045 176 87050 232
rect 87106 176 113190 232
rect 87045 174 113190 176
rect 215250 234 215310 310
rect 218830 308 218836 310
rect 218900 308 218947 312
rect 219526 310 219572 370
rect 219636 368 219683 372
rect 219678 312 219683 368
rect 219566 308 219572 310
rect 219636 308 219683 312
rect 221774 308 221780 372
rect 221844 370 221850 372
rect 222285 370 222351 373
rect 224861 370 224927 373
rect 221844 368 222351 370
rect 221844 312 222290 368
rect 222346 312 222351 368
rect 221844 310 222351 312
rect 221844 308 221850 310
rect 218881 307 218947 308
rect 219617 307 219683 308
rect 222285 307 222351 310
rect 222518 368 224927 370
rect 222518 312 224866 368
rect 224922 312 224927 368
rect 222518 310 224927 312
rect 222518 234 222578 310
rect 224861 307 224927 310
rect 229093 372 229159 373
rect 229829 372 229895 373
rect 229093 368 229140 372
rect 229204 370 229210 372
rect 229093 312 229098 368
rect 229093 308 229140 312
rect 229204 310 229250 370
rect 229829 368 229876 372
rect 229940 370 229946 372
rect 229829 312 229834 368
rect 229204 308 229210 310
rect 229829 308 229876 312
rect 229940 310 229986 370
rect 229940 308 229946 310
rect 230606 308 230612 372
rect 230676 370 230682 372
rect 230841 370 230907 373
rect 230676 368 230907 370
rect 230676 312 230846 368
rect 230902 312 230907 368
rect 230676 310 230907 312
rect 230676 308 230682 310
rect 229093 307 229159 308
rect 229829 307 229895 308
rect 230841 307 230907 310
rect 233417 370 233483 373
rect 233550 370 233556 372
rect 233417 368 233556 370
rect 233417 312 233422 368
rect 233478 312 233556 368
rect 233417 310 233556 312
rect 233417 307 233483 310
rect 233550 308 233556 310
rect 233620 308 233626 372
rect 234153 370 234219 373
rect 234286 370 234292 372
rect 234153 368 234292 370
rect 234153 312 234158 368
rect 234214 312 234292 368
rect 234153 310 234292 312
rect 234153 307 234219 310
rect 234286 308 234292 310
rect 234356 308 234362 372
rect 239581 370 239647 373
rect 234570 368 239647 370
rect 234570 312 239586 368
rect 239642 312 239647 368
rect 234570 310 239647 312
rect 215250 174 222578 234
rect 224033 234 224099 237
rect 234570 234 234630 310
rect 239581 307 239647 310
rect 239714 308 239720 372
rect 239784 370 239790 372
rect 239949 370 240015 373
rect 239784 368 240015 370
rect 239784 312 239954 368
rect 240010 312 240015 368
rect 239784 310 240015 312
rect 239784 308 239790 310
rect 239949 307 240015 310
rect 240450 308 240456 372
rect 240520 370 240526 372
rect 240961 370 241027 373
rect 240520 368 241027 370
rect 240520 312 240966 368
rect 241022 312 241027 368
rect 240520 310 241027 312
rect 240520 308 240526 310
rect 240961 307 241027 310
rect 254434 308 254440 372
rect 254504 370 254510 372
rect 255129 370 255195 373
rect 267690 370 267750 446
rect 269154 444 269160 508
rect 269224 506 269230 508
rect 270033 506 270099 509
rect 269224 504 270099 506
rect 269224 448 270038 504
rect 270094 448 270099 504
rect 269224 446 270099 448
rect 269224 444 269230 446
rect 270033 443 270099 446
rect 254504 368 255195 370
rect 254504 312 255134 368
rect 255190 312 255195 368
rect 254504 310 255195 312
rect 254504 308 254510 310
rect 255129 307 255195 310
rect 263550 310 267750 370
rect 270769 370 270835 373
rect 271362 370 271368 372
rect 270769 368 271368 370
rect 270769 312 270774 368
rect 270830 312 271368 368
rect 270769 310 271368 312
rect 263550 234 263610 310
rect 270769 307 270835 310
rect 271362 308 271368 310
rect 271432 308 271438 372
rect 224033 232 234630 234
rect 224033 176 224038 232
rect 224094 176 234630 232
rect 224033 174 234630 176
rect 239446 174 263610 234
rect 87045 171 87111 174
rect 224033 171 224099 174
rect 180885 98 180951 101
rect 224769 98 224835 101
rect 180885 96 224835 98
rect 180885 40 180890 96
rect 180946 40 224774 96
rect 224830 40 224835 96
rect 180885 38 224835 40
rect 180885 35 180951 38
rect 224769 35 224835 38
rect 224953 98 225019 101
rect 239446 98 239506 174
rect 224953 96 239506 98
rect 224953 40 224958 96
rect 225014 40 239506 96
rect 224953 38 239506 40
rect 239581 98 239647 101
rect 271781 98 271847 101
rect 239581 96 271847 98
rect 239581 40 239586 96
rect 239642 40 271786 96
rect 271842 40 271847 96
rect 239581 38 271847 40
rect 224953 35 225019 38
rect 239581 35 239647 38
rect 271781 35 271847 38
<< via3 >>
rect 9628 10568 9692 10572
rect 9628 10512 9678 10568
rect 9678 10512 9692 10568
rect 9628 10508 9692 10512
rect 20668 10568 20732 10572
rect 20668 10512 20718 10568
rect 20718 10512 20732 10568
rect 20668 10508 20732 10512
rect 71268 10568 71332 10572
rect 71268 10512 71318 10568
rect 71318 10512 71332 10568
rect 71268 10508 71332 10512
rect 74212 10568 74276 10572
rect 74212 10512 74262 10568
rect 74262 10512 74276 10568
rect 74212 10508 74276 10512
rect 84516 10568 84580 10572
rect 84516 10512 84566 10568
rect 84566 10512 84580 10568
rect 84516 10508 84580 10512
rect 86724 10568 86788 10572
rect 86724 10512 86774 10568
rect 86774 10512 86788 10568
rect 86724 10508 86788 10512
rect 207796 10508 207860 10572
rect 218100 10508 218164 10572
rect 54064 10372 54128 10436
rect 72004 10432 72068 10436
rect 72004 10376 72054 10432
rect 72054 10376 72068 10432
rect 72004 10372 72068 10376
rect 77156 10432 77220 10436
rect 77156 10376 77206 10432
rect 77206 10376 77220 10432
rect 77156 10372 77220 10376
rect 82308 10432 82372 10436
rect 82308 10376 82358 10432
rect 82358 10376 82372 10432
rect 82308 10372 82372 10376
rect 83780 10432 83844 10436
rect 83780 10376 83830 10432
rect 83830 10376 83844 10432
rect 83780 10372 83844 10376
rect 125272 10432 125336 10436
rect 125272 10376 125322 10432
rect 125322 10376 125336 10432
rect 125272 10372 125336 10376
rect 128216 10372 128280 10436
rect 147628 10372 147692 10436
rect 181760 10432 181824 10436
rect 181760 10376 181810 10432
rect 181810 10376 181824 10432
rect 181760 10372 181824 10376
rect 190592 10372 190656 10436
rect 193536 10372 193600 10436
rect 198688 10372 198752 10436
rect 200896 10432 200960 10436
rect 200896 10376 200946 10432
rect 200946 10376 200960 10432
rect 200896 10372 200960 10376
rect 202368 10372 202432 10436
rect 210004 10372 210068 10436
rect 211476 10372 211540 10436
rect 221044 10372 221108 10436
rect 261064 10372 261128 10436
rect 264744 10372 264808 10436
rect 31708 10296 31772 10300
rect 31708 10240 31758 10296
rect 31758 10240 31772 10296
rect 31708 10236 31772 10240
rect 34928 10236 34992 10300
rect 35664 10296 35728 10300
rect 35664 10240 35678 10296
rect 35678 10240 35728 10296
rect 35664 10236 35728 10240
rect 36400 10236 36464 10300
rect 37136 10236 37200 10300
rect 37872 10236 37936 10300
rect 38608 10236 38672 10300
rect 39344 10236 39408 10300
rect 40080 10236 40144 10300
rect 40816 10296 40880 10300
rect 40816 10240 40830 10296
rect 40830 10240 40880 10296
rect 40816 10236 40880 10240
rect 41552 10236 41616 10300
rect 42288 10236 42352 10300
rect 43024 10236 43088 10300
rect 43760 10236 43824 10300
rect 44496 10236 44560 10300
rect 45232 10236 45296 10300
rect 45968 10296 46032 10300
rect 45968 10240 45982 10296
rect 45982 10240 46032 10296
rect 45968 10236 46032 10240
rect 46704 10236 46768 10300
rect 47440 10236 47504 10300
rect 48176 10296 48240 10300
rect 48176 10240 48226 10296
rect 48226 10240 48240 10296
rect 48176 10236 48240 10240
rect 48912 10236 48976 10300
rect 49648 10236 49712 10300
rect 50384 10236 50448 10300
rect 51120 10236 51184 10300
rect 51856 10236 51920 10300
rect 52592 10236 52656 10300
rect 53328 10236 53392 10300
rect 54800 10296 54864 10300
rect 54800 10240 54814 10296
rect 54814 10240 54864 10296
rect 54800 10236 54864 10240
rect 55536 10296 55600 10300
rect 55536 10240 55550 10296
rect 55550 10240 55600 10296
rect 55536 10236 55600 10240
rect 56272 10296 56336 10300
rect 56272 10240 56286 10296
rect 56286 10240 56336 10296
rect 56272 10236 56336 10240
rect 57008 10296 57072 10300
rect 57008 10240 57058 10296
rect 57058 10240 57072 10296
rect 57008 10236 57072 10240
rect 57744 10296 57808 10300
rect 57744 10240 57794 10296
rect 57794 10240 57808 10296
rect 57744 10236 57808 10240
rect 58480 10236 58544 10300
rect 59216 10296 59280 10300
rect 59216 10240 59266 10296
rect 59266 10240 59280 10296
rect 59216 10236 59280 10240
rect 59952 10296 60016 10300
rect 59952 10240 60002 10296
rect 60002 10240 60016 10296
rect 59952 10236 60016 10240
rect 60688 10236 60752 10300
rect 61424 10236 61488 10300
rect 62160 10236 62224 10300
rect 62896 10236 62960 10300
rect 63632 10236 63696 10300
rect 64368 10236 64432 10300
rect 65104 10236 65168 10300
rect 65840 10236 65904 10300
rect 66576 10236 66640 10300
rect 89668 10236 89732 10300
rect 103192 10296 103256 10300
rect 103192 10240 103242 10296
rect 103242 10240 103256 10296
rect 103192 10236 103256 10240
rect 103928 10296 103992 10300
rect 103928 10240 103942 10296
rect 103942 10240 103992 10296
rect 103928 10236 103992 10240
rect 104664 10236 104728 10300
rect 105400 10236 105464 10300
rect 106136 10236 106200 10300
rect 106872 10236 106936 10300
rect 107608 10236 107672 10300
rect 108344 10296 108408 10300
rect 108344 10240 108394 10296
rect 108394 10240 108408 10296
rect 108344 10236 108408 10240
rect 109080 10296 109144 10300
rect 109080 10240 109094 10296
rect 109094 10240 109144 10296
rect 109080 10236 109144 10240
rect 109816 10236 109880 10300
rect 110552 10236 110616 10300
rect 111288 10236 111352 10300
rect 112024 10236 112088 10300
rect 112760 10236 112824 10300
rect 113496 10296 113560 10300
rect 113496 10240 113546 10296
rect 113546 10240 113560 10296
rect 113496 10236 113560 10240
rect 114232 10296 114296 10300
rect 114232 10240 114246 10296
rect 114246 10240 114296 10296
rect 114232 10236 114296 10240
rect 114968 10236 115032 10300
rect 115704 10236 115768 10300
rect 116440 10236 116504 10300
rect 117176 10236 117240 10300
rect 117912 10236 117976 10300
rect 118648 10296 118712 10300
rect 118648 10240 118698 10296
rect 118698 10240 118712 10296
rect 118648 10236 118712 10240
rect 119384 10296 119448 10300
rect 119384 10240 119398 10296
rect 119398 10240 119448 10296
rect 119384 10236 119448 10240
rect 120120 10236 120184 10300
rect 120856 10236 120920 10300
rect 121592 10236 121656 10300
rect 122328 10236 122392 10300
rect 123064 10236 123128 10300
rect 123800 10236 123864 10300
rect 124536 10236 124600 10300
rect 126008 10236 126072 10300
rect 126744 10296 126808 10300
rect 126744 10240 126794 10296
rect 126794 10240 126808 10296
rect 126744 10236 126808 10240
rect 127480 10236 127544 10300
rect 128952 10236 129016 10300
rect 129688 10296 129752 10300
rect 129688 10240 129702 10296
rect 129702 10240 129752 10296
rect 129688 10236 129752 10240
rect 130424 10296 130488 10300
rect 130424 10240 130474 10296
rect 130474 10240 130488 10296
rect 130424 10236 130488 10240
rect 131160 10236 131224 10300
rect 131896 10236 131960 10300
rect 132632 10236 132696 10300
rect 133368 10236 133432 10300
rect 134104 10236 134168 10300
rect 134840 10296 134904 10300
rect 134840 10240 134890 10296
rect 134890 10240 134904 10296
rect 134840 10236 134904 10240
rect 138060 10236 138124 10300
rect 142476 10236 142540 10300
rect 153516 10236 153580 10300
rect 157196 10296 157260 10300
rect 157196 10240 157246 10296
rect 157246 10240 157260 10296
rect 157196 10236 157260 10240
rect 171456 10236 171520 10300
rect 172192 10236 172256 10300
rect 172928 10236 172992 10300
rect 173664 10296 173728 10300
rect 173664 10240 173714 10296
rect 173714 10240 173728 10296
rect 173664 10236 173728 10240
rect 174400 10296 174464 10300
rect 174400 10240 174450 10296
rect 174450 10240 174464 10296
rect 174400 10236 174464 10240
rect 175136 10296 175200 10300
rect 175136 10240 175186 10296
rect 175186 10240 175200 10296
rect 175136 10236 175200 10240
rect 175872 10296 175936 10300
rect 175872 10240 175922 10296
rect 175922 10240 175936 10296
rect 175872 10236 175936 10240
rect 176608 10236 176672 10300
rect 177344 10236 177408 10300
rect 178080 10236 178144 10300
rect 178816 10236 178880 10300
rect 179552 10296 179616 10300
rect 179552 10240 179602 10296
rect 179602 10240 179616 10296
rect 179552 10236 179616 10240
rect 180288 10296 180352 10300
rect 180288 10240 180338 10296
rect 180338 10240 180352 10296
rect 180288 10236 180352 10240
rect 181024 10236 181088 10300
rect 182496 10296 182560 10300
rect 182496 10240 182546 10296
rect 182546 10240 182560 10296
rect 182496 10236 182560 10240
rect 183232 10296 183296 10300
rect 183232 10240 183282 10296
rect 183282 10240 183296 10296
rect 183232 10236 183296 10240
rect 183968 10236 184032 10300
rect 184704 10296 184768 10300
rect 184704 10240 184754 10296
rect 184754 10240 184768 10296
rect 184704 10236 184768 10240
rect 185440 10296 185504 10300
rect 185440 10240 185490 10296
rect 185490 10240 185504 10296
rect 185440 10236 185504 10240
rect 186176 10296 186240 10300
rect 186176 10240 186226 10296
rect 186226 10240 186240 10296
rect 186176 10236 186240 10240
rect 186912 10296 186976 10300
rect 186912 10240 186962 10296
rect 186962 10240 186976 10296
rect 186912 10236 186976 10240
rect 187648 10296 187712 10300
rect 187648 10240 187698 10296
rect 187698 10240 187712 10296
rect 187648 10236 187712 10240
rect 188384 10296 188448 10300
rect 188384 10240 188434 10296
rect 188434 10240 188448 10296
rect 188384 10236 188448 10240
rect 189120 10236 189184 10300
rect 189856 10296 189920 10300
rect 189856 10240 189906 10296
rect 189906 10240 189920 10296
rect 189856 10236 189920 10240
rect 191328 10296 191392 10300
rect 191328 10240 191378 10296
rect 191378 10240 191392 10296
rect 191328 10236 191392 10240
rect 192064 10236 192128 10300
rect 192800 10296 192864 10300
rect 192800 10240 192850 10296
rect 192850 10240 192864 10296
rect 192800 10236 192864 10240
rect 194272 10296 194336 10300
rect 194272 10240 194322 10296
rect 194322 10240 194336 10296
rect 194272 10236 194336 10240
rect 195008 10236 195072 10300
rect 195744 10296 195808 10300
rect 195744 10240 195794 10296
rect 195794 10240 195808 10296
rect 195744 10236 195808 10240
rect 196480 10296 196544 10300
rect 196480 10240 196530 10296
rect 196530 10240 196544 10296
rect 196480 10236 196544 10240
rect 197216 10296 197280 10300
rect 197216 10240 197266 10296
rect 197266 10240 197280 10296
rect 197216 10236 197280 10240
rect 197952 10296 198016 10300
rect 197952 10240 198002 10296
rect 198002 10240 198016 10296
rect 197952 10236 198016 10240
rect 199424 10236 199488 10300
rect 200160 10236 200224 10300
rect 201632 10236 201696 10300
rect 203104 10236 203168 10300
rect 215156 10236 215220 10300
rect 220308 10236 220372 10300
rect 221780 10236 221844 10300
rect 222516 10236 222580 10300
rect 239720 10296 239784 10300
rect 239720 10240 239734 10296
rect 239734 10240 239784 10296
rect 239720 10236 239784 10240
rect 240456 10236 240520 10300
rect 241192 10296 241256 10300
rect 241192 10240 241242 10296
rect 241242 10240 241256 10296
rect 241192 10236 241256 10240
rect 241928 10296 241992 10300
rect 241928 10240 241978 10296
rect 241978 10240 241992 10296
rect 241928 10236 241992 10240
rect 242664 10296 242728 10300
rect 242664 10240 242714 10296
rect 242714 10240 242728 10296
rect 242664 10236 242728 10240
rect 243400 10296 243464 10300
rect 243400 10240 243450 10296
rect 243450 10240 243464 10296
rect 243400 10236 243464 10240
rect 244136 10296 244200 10300
rect 244136 10240 244186 10296
rect 244186 10240 244200 10296
rect 244136 10236 244200 10240
rect 244872 10296 244936 10300
rect 244872 10240 244922 10296
rect 244922 10240 244936 10296
rect 244872 10236 244936 10240
rect 245608 10236 245672 10300
rect 246344 10296 246408 10300
rect 246344 10240 246394 10296
rect 246394 10240 246408 10296
rect 246344 10236 246408 10240
rect 247080 10236 247144 10300
rect 247816 10296 247880 10300
rect 247816 10240 247866 10296
rect 247866 10240 247880 10296
rect 247816 10236 247880 10240
rect 248552 10236 248616 10300
rect 249288 10296 249352 10300
rect 249288 10240 249338 10296
rect 249338 10240 249352 10296
rect 249288 10236 249352 10240
rect 250024 10296 250088 10300
rect 250024 10240 250074 10296
rect 250074 10240 250088 10296
rect 250024 10236 250088 10240
rect 250760 10296 250824 10300
rect 250760 10240 250810 10296
rect 250810 10240 250824 10296
rect 250760 10236 250824 10240
rect 251496 10296 251560 10300
rect 251496 10240 251546 10296
rect 251546 10240 251560 10296
rect 251496 10236 251560 10240
rect 252232 10296 252296 10300
rect 252232 10240 252282 10296
rect 252282 10240 252296 10296
rect 252232 10236 252296 10240
rect 252968 10236 253032 10300
rect 253704 10236 253768 10300
rect 254440 10296 254504 10300
rect 254440 10240 254490 10296
rect 254490 10240 254504 10296
rect 254440 10236 254504 10240
rect 255176 10296 255240 10300
rect 255176 10240 255226 10296
rect 255226 10240 255240 10296
rect 255176 10236 255240 10240
rect 255912 10236 255976 10300
rect 256648 10296 256712 10300
rect 256648 10240 256698 10296
rect 256698 10240 256712 10296
rect 256648 10236 256712 10240
rect 257384 10236 257448 10300
rect 258120 10236 258184 10300
rect 258856 10236 258920 10300
rect 259592 10236 259656 10300
rect 260328 10236 260392 10300
rect 261800 10296 261864 10300
rect 261800 10240 261814 10296
rect 261814 10240 261864 10296
rect 261800 10236 261864 10240
rect 262536 10296 262600 10300
rect 262536 10240 262550 10296
rect 262550 10240 262600 10296
rect 262536 10236 262600 10240
rect 263272 10296 263336 10300
rect 263272 10240 263286 10296
rect 263286 10240 263336 10296
rect 263272 10236 263336 10240
rect 264008 10236 264072 10300
rect 265480 10236 265544 10300
rect 1532 10100 1596 10164
rect 2268 10100 2332 10164
rect 3740 10100 3804 10164
rect 4476 10100 4540 10164
rect 5212 10100 5276 10164
rect 5948 10100 6012 10164
rect 6684 10100 6748 10164
rect 7420 10100 7484 10164
rect 8892 10100 8956 10164
rect 11836 10100 11900 10164
rect 12572 10100 12636 10164
rect 14044 10100 14108 10164
rect 14780 10100 14844 10164
rect 15516 10100 15580 10164
rect 16252 10100 16316 10164
rect 16988 10100 17052 10164
rect 17724 10100 17788 10164
rect 18460 10100 18524 10164
rect 22140 10100 22204 10164
rect 138796 10160 138860 10164
rect 138796 10104 138846 10160
rect 138846 10104 138860 10160
rect 138796 10100 138860 10104
rect 140268 10100 140332 10164
rect 141004 10100 141068 10164
rect 141740 10100 141804 10164
rect 143212 10100 143276 10164
rect 143948 10100 144012 10164
rect 145420 10100 145484 10164
rect 146156 10160 146220 10164
rect 146156 10104 146206 10160
rect 146206 10104 146220 10160
rect 146156 10100 146220 10104
rect 146892 10100 146956 10164
rect 148364 10100 148428 10164
rect 149100 10100 149164 10164
rect 150572 10100 150636 10164
rect 151308 10100 151372 10164
rect 152044 10100 152108 10164
rect 152780 10100 152844 10164
rect 154252 10100 154316 10164
rect 206324 10100 206388 10164
rect 207060 10100 207124 10164
rect 208532 10100 208596 10164
rect 209268 10160 209332 10164
rect 209268 10104 209318 10160
rect 209318 10104 209332 10160
rect 209268 10100 209332 10104
rect 210740 10160 210804 10164
rect 210740 10104 210790 10160
rect 210790 10104 210804 10160
rect 210740 10100 210804 10104
rect 212948 10100 213012 10164
rect 213684 10100 213748 10164
rect 214420 10100 214484 10164
rect 215892 10100 215956 10164
rect 217364 10100 217428 10164
rect 218836 10100 218900 10164
rect 219572 10100 219636 10164
rect 223252 10160 223316 10164
rect 223252 10104 223302 10160
rect 223302 10104 223316 10160
rect 223252 10100 223316 10104
rect 3004 9828 3068 9892
rect 8156 9888 8220 9892
rect 8156 9832 8206 9888
rect 8206 9832 8220 9888
rect 8156 9828 8220 9832
rect 10364 9828 10428 9892
rect 11100 9828 11164 9892
rect 13308 9828 13372 9892
rect 21404 9888 21468 9892
rect 21404 9832 21454 9888
rect 21454 9832 21468 9888
rect 21404 9828 21468 9832
rect 85252 9828 85316 9892
rect 85988 9828 86052 9892
rect 139532 9828 139596 9892
rect 144684 9888 144748 9892
rect 144684 9832 144734 9888
rect 144734 9832 144748 9888
rect 144684 9828 144748 9832
rect 149836 9828 149900 9892
rect 154988 9828 155052 9892
rect 216628 9828 216692 9892
rect 68548 9820 68612 9824
rect 68548 9764 68552 9820
rect 68552 9764 68608 9820
rect 68608 9764 68612 9820
rect 68548 9760 68612 9764
rect 68628 9820 68692 9824
rect 68628 9764 68632 9820
rect 68632 9764 68688 9820
rect 68688 9764 68692 9820
rect 68628 9760 68692 9764
rect 68708 9820 68772 9824
rect 68708 9764 68712 9820
rect 68712 9764 68768 9820
rect 68768 9764 68772 9820
rect 68708 9760 68772 9764
rect 68788 9820 68852 9824
rect 68788 9764 68792 9820
rect 68792 9764 68848 9820
rect 68848 9764 68852 9820
rect 68788 9760 68852 9764
rect 136145 9820 136209 9824
rect 136145 9764 136149 9820
rect 136149 9764 136205 9820
rect 136205 9764 136209 9820
rect 136145 9760 136209 9764
rect 136225 9820 136289 9824
rect 136225 9764 136229 9820
rect 136229 9764 136285 9820
rect 136285 9764 136289 9820
rect 136225 9760 136289 9764
rect 136305 9820 136369 9824
rect 136305 9764 136309 9820
rect 136309 9764 136365 9820
rect 136365 9764 136369 9820
rect 136305 9760 136369 9764
rect 136385 9820 136449 9824
rect 136385 9764 136389 9820
rect 136389 9764 136445 9820
rect 136445 9764 136449 9820
rect 136385 9760 136449 9764
rect 203742 9820 203806 9824
rect 203742 9764 203746 9820
rect 203746 9764 203802 9820
rect 203802 9764 203806 9820
rect 203742 9760 203806 9764
rect 203822 9820 203886 9824
rect 203822 9764 203826 9820
rect 203826 9764 203882 9820
rect 203882 9764 203886 9820
rect 203822 9760 203886 9764
rect 203902 9820 203966 9824
rect 203902 9764 203906 9820
rect 203906 9764 203962 9820
rect 203962 9764 203966 9820
rect 203902 9760 203966 9764
rect 203982 9820 204046 9824
rect 203982 9764 203986 9820
rect 203986 9764 204042 9820
rect 204042 9764 204046 9820
rect 203982 9760 204046 9764
rect 271339 9820 271403 9824
rect 271339 9764 271343 9820
rect 271343 9764 271399 9820
rect 271399 9764 271403 9820
rect 271339 9760 271403 9764
rect 271419 9820 271483 9824
rect 271419 9764 271423 9820
rect 271423 9764 271479 9820
rect 271479 9764 271483 9820
rect 271419 9760 271483 9764
rect 271499 9820 271563 9824
rect 271499 9764 271503 9820
rect 271503 9764 271559 9820
rect 271559 9764 271563 9820
rect 271499 9760 271563 9764
rect 271579 9820 271643 9824
rect 271579 9764 271583 9820
rect 271583 9764 271639 9820
rect 271639 9764 271643 9820
rect 271579 9760 271643 9764
rect 76420 9752 76484 9756
rect 76420 9696 76470 9752
rect 76470 9696 76484 9752
rect 76420 9692 76484 9696
rect 79364 9752 79428 9756
rect 79364 9696 79414 9752
rect 79414 9696 79428 9752
rect 79364 9692 79428 9696
rect 81572 9752 81636 9756
rect 81572 9696 81622 9752
rect 81622 9696 81636 9752
rect 81572 9692 81636 9696
rect 93348 9692 93412 9756
rect 95556 9692 95620 9756
rect 96292 9752 96356 9756
rect 96292 9696 96342 9752
rect 96342 9696 96356 9752
rect 96292 9692 96356 9696
rect 97764 9692 97828 9756
rect 100708 9752 100772 9756
rect 100708 9696 100722 9752
rect 100722 9696 100772 9752
rect 100708 9692 100772 9696
rect 155724 9692 155788 9756
rect 156460 9692 156524 9756
rect 157932 9752 157996 9756
rect 157932 9696 157982 9752
rect 157982 9696 157996 9752
rect 157932 9692 157996 9696
rect 159404 9752 159468 9756
rect 159404 9696 159454 9752
rect 159454 9696 159468 9752
rect 159404 9692 159468 9696
rect 163820 9752 163884 9756
rect 163820 9696 163870 9752
rect 163870 9696 163884 9752
rect 163820 9692 163884 9696
rect 225460 9692 225524 9756
rect 229876 9752 229940 9756
rect 229876 9696 229890 9752
rect 229890 9696 229940 9752
rect 229876 9692 229940 9696
rect 231348 9692 231412 9756
rect 233556 9752 233620 9756
rect 233556 9696 233570 9752
rect 233570 9696 233620 9752
rect 233556 9692 233620 9696
rect 234292 9752 234356 9756
rect 234292 9696 234342 9752
rect 234342 9696 234356 9752
rect 234292 9692 234356 9696
rect 235028 9752 235092 9756
rect 235028 9696 235078 9752
rect 235078 9696 235092 9752
rect 235028 9692 235092 9696
rect 25820 9616 25884 9620
rect 25820 9560 25870 9616
rect 25870 9560 25884 9616
rect 25820 9556 25884 9560
rect 32444 9556 32508 9620
rect 69060 9616 69124 9620
rect 69060 9560 69110 9616
rect 69110 9560 69124 9616
rect 69060 9556 69124 9560
rect 70532 9556 70596 9620
rect 72740 9556 72804 9620
rect 75684 9556 75748 9620
rect 77892 9556 77956 9620
rect 80836 9556 80900 9620
rect 83044 9556 83108 9620
rect 137324 9616 137388 9620
rect 137324 9560 137374 9616
rect 137374 9560 137388 9616
rect 137324 9556 137388 9560
rect 205588 9556 205652 9620
rect 28764 9480 28828 9484
rect 28764 9424 28814 9480
rect 28814 9424 28828 9480
rect 28764 9420 28828 9424
rect 158668 9420 158732 9484
rect 228404 9420 228468 9484
rect 34750 9276 34814 9280
rect 34750 9220 34754 9276
rect 34754 9220 34810 9276
rect 34810 9220 34814 9276
rect 34750 9216 34814 9220
rect 34830 9276 34894 9280
rect 34830 9220 34834 9276
rect 34834 9220 34890 9276
rect 34890 9220 34894 9276
rect 34830 9216 34894 9220
rect 34910 9276 34974 9280
rect 34910 9220 34914 9276
rect 34914 9220 34970 9276
rect 34970 9220 34974 9276
rect 34910 9216 34974 9220
rect 34990 9276 35054 9280
rect 34990 9220 34994 9276
rect 34994 9220 35050 9276
rect 35050 9220 35054 9276
rect 34990 9216 35054 9220
rect 102347 9276 102411 9280
rect 102347 9220 102351 9276
rect 102351 9220 102407 9276
rect 102407 9220 102411 9276
rect 102347 9216 102411 9220
rect 102427 9276 102491 9280
rect 102427 9220 102431 9276
rect 102431 9220 102487 9276
rect 102487 9220 102491 9276
rect 102427 9216 102491 9220
rect 102507 9276 102571 9280
rect 102507 9220 102511 9276
rect 102511 9220 102567 9276
rect 102567 9220 102571 9276
rect 102507 9216 102571 9220
rect 102587 9276 102651 9280
rect 102587 9220 102591 9276
rect 102591 9220 102647 9276
rect 102647 9220 102651 9276
rect 102587 9216 102651 9220
rect 169944 9276 170008 9280
rect 169944 9220 169948 9276
rect 169948 9220 170004 9276
rect 170004 9220 170008 9276
rect 169944 9216 170008 9220
rect 170024 9276 170088 9280
rect 170024 9220 170028 9276
rect 170028 9220 170084 9276
rect 170084 9220 170088 9276
rect 170024 9216 170088 9220
rect 170104 9276 170168 9280
rect 170104 9220 170108 9276
rect 170108 9220 170164 9276
rect 170164 9220 170168 9276
rect 170104 9216 170168 9220
rect 170184 9276 170248 9280
rect 170184 9220 170188 9276
rect 170188 9220 170244 9276
rect 170244 9220 170248 9276
rect 170184 9216 170248 9220
rect 237541 9276 237605 9280
rect 237541 9220 237545 9276
rect 237545 9220 237601 9276
rect 237601 9220 237605 9276
rect 237541 9216 237605 9220
rect 237621 9276 237685 9280
rect 237621 9220 237625 9276
rect 237625 9220 237681 9276
rect 237681 9220 237685 9276
rect 237621 9216 237685 9220
rect 237701 9276 237765 9280
rect 237701 9220 237705 9276
rect 237705 9220 237761 9276
rect 237761 9220 237765 9276
rect 237701 9216 237765 9220
rect 237781 9276 237845 9280
rect 237781 9220 237785 9276
rect 237785 9220 237841 9276
rect 237841 9220 237845 9276
rect 237781 9216 237845 9220
rect 796 9148 860 9212
rect 88196 9148 88260 9212
rect 168972 9208 169036 9212
rect 168972 9152 169022 9208
rect 169022 9152 169036 9208
rect 168972 9148 169036 9152
rect 223988 9148 224052 9212
rect 235764 9148 235828 9212
rect 237236 9208 237300 9212
rect 237236 9152 237286 9208
rect 237286 9152 237300 9208
rect 237236 9148 237300 9152
rect 69796 9012 69860 9076
rect 73476 9072 73540 9076
rect 73476 9016 73490 9072
rect 73490 9016 73540 9072
rect 73476 9012 73540 9016
rect 74948 9012 75012 9076
rect 78628 9072 78692 9076
rect 78628 9016 78642 9072
rect 78642 9016 78692 9072
rect 78628 9012 78692 9016
rect 80100 9012 80164 9076
rect 91140 8740 91204 8804
rect 262076 8740 262140 8804
rect 68548 8732 68612 8736
rect 68548 8676 68552 8732
rect 68552 8676 68608 8732
rect 68608 8676 68612 8732
rect 68548 8672 68612 8676
rect 68628 8732 68692 8736
rect 68628 8676 68632 8732
rect 68632 8676 68688 8732
rect 68688 8676 68692 8732
rect 68628 8672 68692 8676
rect 68708 8732 68772 8736
rect 68708 8676 68712 8732
rect 68712 8676 68768 8732
rect 68768 8676 68772 8732
rect 68708 8672 68772 8676
rect 68788 8732 68852 8736
rect 68788 8676 68792 8732
rect 68792 8676 68848 8732
rect 68848 8676 68852 8732
rect 68788 8672 68852 8676
rect 136145 8732 136209 8736
rect 136145 8676 136149 8732
rect 136149 8676 136205 8732
rect 136205 8676 136209 8732
rect 136145 8672 136209 8676
rect 136225 8732 136289 8736
rect 136225 8676 136229 8732
rect 136229 8676 136285 8732
rect 136285 8676 136289 8732
rect 136225 8672 136289 8676
rect 136305 8732 136369 8736
rect 136305 8676 136309 8732
rect 136309 8676 136365 8732
rect 136365 8676 136369 8732
rect 136305 8672 136369 8676
rect 136385 8732 136449 8736
rect 136385 8676 136389 8732
rect 136389 8676 136445 8732
rect 136445 8676 136449 8732
rect 136385 8672 136449 8676
rect 203742 8732 203806 8736
rect 203742 8676 203746 8732
rect 203746 8676 203802 8732
rect 203802 8676 203806 8732
rect 203742 8672 203806 8676
rect 203822 8732 203886 8736
rect 203822 8676 203826 8732
rect 203826 8676 203882 8732
rect 203882 8676 203886 8732
rect 203822 8672 203886 8676
rect 203902 8732 203966 8736
rect 203902 8676 203906 8732
rect 203906 8676 203962 8732
rect 203962 8676 203966 8732
rect 203902 8672 203966 8676
rect 203982 8732 204046 8736
rect 203982 8676 203986 8732
rect 203986 8676 204042 8732
rect 204042 8676 204046 8732
rect 203982 8672 204046 8676
rect 271339 8732 271403 8736
rect 271339 8676 271343 8732
rect 271343 8676 271399 8732
rect 271399 8676 271403 8732
rect 271339 8672 271403 8676
rect 271419 8732 271483 8736
rect 271419 8676 271423 8732
rect 271423 8676 271479 8732
rect 271479 8676 271483 8732
rect 271419 8672 271483 8676
rect 271499 8732 271563 8736
rect 271499 8676 271503 8732
rect 271503 8676 271559 8732
rect 271559 8676 271563 8732
rect 271499 8672 271563 8676
rect 271579 8732 271643 8736
rect 271579 8676 271583 8732
rect 271583 8676 271639 8732
rect 271639 8676 271643 8732
rect 271579 8672 271643 8676
rect 24348 8604 24412 8668
rect 29500 8604 29564 8668
rect 30236 8664 30300 8668
rect 30236 8608 30250 8664
rect 30250 8608 30300 8664
rect 30236 8604 30300 8608
rect 30972 8604 31036 8668
rect 87460 8604 87524 8668
rect 90404 8664 90468 8668
rect 90404 8608 90454 8664
rect 90454 8608 90468 8664
rect 90404 8604 90468 8608
rect 91876 8664 91940 8668
rect 91876 8608 91926 8664
rect 91926 8608 91940 8664
rect 91876 8604 91940 8608
rect 94084 8604 94148 8668
rect 94820 8664 94884 8668
rect 94820 8608 94870 8664
rect 94870 8608 94884 8664
rect 94820 8604 94884 8608
rect 97028 8604 97092 8668
rect 98500 8604 98564 8668
rect 99972 8604 100036 8668
rect 226196 8604 226260 8668
rect 226932 8604 226996 8668
rect 227668 8604 227732 8668
rect 229140 8664 229204 8668
rect 229140 8608 229154 8664
rect 229154 8608 229204 8664
rect 229140 8604 229204 8608
rect 232084 8604 232148 8668
rect 232820 8664 232884 8668
rect 232820 8608 232870 8664
rect 232870 8608 232884 8664
rect 232820 8604 232884 8608
rect 236500 8604 236564 8668
rect 161612 8468 161676 8532
rect 26556 8332 26620 8396
rect 28028 8332 28092 8396
rect 92612 8332 92676 8396
rect 160140 8332 160204 8396
rect 160876 8332 160940 8396
rect 162348 8332 162412 8396
rect 163084 8332 163148 8396
rect 164556 8332 164620 8396
rect 165292 8332 165356 8396
rect 166028 8332 166092 8396
rect 167500 8332 167564 8396
rect 224724 8392 224788 8396
rect 224724 8336 224774 8392
rect 224774 8336 224788 8392
rect 224724 8332 224788 8336
rect 230612 8332 230676 8396
rect 263180 8332 263244 8396
rect 99236 8256 99300 8260
rect 99236 8200 99286 8256
rect 99286 8200 99300 8256
rect 99236 8196 99300 8200
rect 166764 8256 166828 8260
rect 166764 8200 166814 8256
rect 166814 8200 166828 8256
rect 166764 8196 166828 8200
rect 266492 8392 266556 8396
rect 266492 8336 266506 8392
rect 266506 8336 266556 8392
rect 266492 8332 266556 8336
rect 34750 8188 34814 8192
rect 34750 8132 34754 8188
rect 34754 8132 34810 8188
rect 34810 8132 34814 8188
rect 34750 8128 34814 8132
rect 34830 8188 34894 8192
rect 34830 8132 34834 8188
rect 34834 8132 34890 8188
rect 34890 8132 34894 8188
rect 34830 8128 34894 8132
rect 34910 8188 34974 8192
rect 34910 8132 34914 8188
rect 34914 8132 34970 8188
rect 34970 8132 34974 8188
rect 34910 8128 34974 8132
rect 34990 8188 35054 8192
rect 34990 8132 34994 8188
rect 34994 8132 35050 8188
rect 35050 8132 35054 8188
rect 34990 8128 35054 8132
rect 102347 8188 102411 8192
rect 102347 8132 102351 8188
rect 102351 8132 102407 8188
rect 102407 8132 102411 8188
rect 102347 8128 102411 8132
rect 102427 8188 102491 8192
rect 102427 8132 102431 8188
rect 102431 8132 102487 8188
rect 102487 8132 102491 8188
rect 102427 8128 102491 8132
rect 102507 8188 102571 8192
rect 102507 8132 102511 8188
rect 102511 8132 102567 8188
rect 102567 8132 102571 8188
rect 102507 8128 102571 8132
rect 102587 8188 102651 8192
rect 102587 8132 102591 8188
rect 102591 8132 102647 8188
rect 102647 8132 102651 8188
rect 102587 8128 102651 8132
rect 169944 8188 170008 8192
rect 169944 8132 169948 8188
rect 169948 8132 170004 8188
rect 170004 8132 170008 8188
rect 169944 8128 170008 8132
rect 170024 8188 170088 8192
rect 170024 8132 170028 8188
rect 170028 8132 170084 8188
rect 170084 8132 170088 8188
rect 170024 8128 170088 8132
rect 170104 8188 170168 8192
rect 170104 8132 170108 8188
rect 170108 8132 170164 8188
rect 170164 8132 170168 8188
rect 170104 8128 170168 8132
rect 170184 8188 170248 8192
rect 170184 8132 170188 8188
rect 170188 8132 170244 8188
rect 170244 8132 170248 8188
rect 170184 8128 170248 8132
rect 237541 8188 237605 8192
rect 237541 8132 237545 8188
rect 237545 8132 237601 8188
rect 237601 8132 237605 8188
rect 237541 8128 237605 8132
rect 237621 8188 237685 8192
rect 237621 8132 237625 8188
rect 237625 8132 237681 8188
rect 237681 8132 237685 8188
rect 237621 8128 237685 8132
rect 237701 8188 237765 8192
rect 237701 8132 237705 8188
rect 237705 8132 237761 8188
rect 237761 8132 237765 8188
rect 237701 8128 237765 8132
rect 237781 8188 237845 8192
rect 237781 8132 237785 8188
rect 237785 8132 237841 8188
rect 237841 8132 237845 8188
rect 237781 8128 237845 8132
rect 88932 8060 88996 8124
rect 168236 8060 168300 8124
rect 27292 7788 27356 7852
rect 68548 7644 68612 7648
rect 68548 7588 68552 7644
rect 68552 7588 68608 7644
rect 68608 7588 68612 7644
rect 68548 7584 68612 7588
rect 68628 7644 68692 7648
rect 68628 7588 68632 7644
rect 68632 7588 68688 7644
rect 68688 7588 68692 7644
rect 68628 7584 68692 7588
rect 68708 7644 68772 7648
rect 68708 7588 68712 7644
rect 68712 7588 68768 7644
rect 68768 7588 68772 7644
rect 68708 7584 68772 7588
rect 68788 7644 68852 7648
rect 68788 7588 68792 7644
rect 68792 7588 68848 7644
rect 68848 7588 68852 7644
rect 68788 7584 68852 7588
rect 136145 7644 136209 7648
rect 136145 7588 136149 7644
rect 136149 7588 136205 7644
rect 136205 7588 136209 7644
rect 136145 7584 136209 7588
rect 136225 7644 136289 7648
rect 136225 7588 136229 7644
rect 136229 7588 136285 7644
rect 136285 7588 136289 7644
rect 136225 7584 136289 7588
rect 136305 7644 136369 7648
rect 136305 7588 136309 7644
rect 136309 7588 136365 7644
rect 136365 7588 136369 7644
rect 136305 7584 136369 7588
rect 136385 7644 136449 7648
rect 136385 7588 136389 7644
rect 136389 7588 136445 7644
rect 136445 7588 136449 7644
rect 136385 7584 136449 7588
rect 203742 7644 203806 7648
rect 203742 7588 203746 7644
rect 203746 7588 203802 7644
rect 203802 7588 203806 7644
rect 203742 7584 203806 7588
rect 203822 7644 203886 7648
rect 203822 7588 203826 7644
rect 203826 7588 203882 7644
rect 203882 7588 203886 7644
rect 203822 7584 203886 7588
rect 203902 7644 203966 7648
rect 203902 7588 203906 7644
rect 203906 7588 203962 7644
rect 203962 7588 203966 7644
rect 203902 7584 203966 7588
rect 203982 7644 204046 7648
rect 203982 7588 203986 7644
rect 203986 7588 204042 7644
rect 204042 7588 204046 7644
rect 203982 7584 204046 7588
rect 267412 7652 267476 7716
rect 271339 7644 271403 7648
rect 271339 7588 271343 7644
rect 271343 7588 271399 7644
rect 271399 7588 271403 7644
rect 271339 7584 271403 7588
rect 271419 7644 271483 7648
rect 271419 7588 271423 7644
rect 271423 7588 271479 7644
rect 271479 7588 271483 7644
rect 271419 7584 271483 7588
rect 271499 7644 271563 7648
rect 271499 7588 271503 7644
rect 271503 7588 271559 7644
rect 271559 7588 271563 7644
rect 271499 7584 271563 7588
rect 271579 7644 271643 7648
rect 271579 7588 271583 7644
rect 271583 7588 271639 7644
rect 271639 7588 271643 7644
rect 271579 7584 271643 7588
rect 267964 7516 268028 7580
rect 34750 7100 34814 7104
rect 34750 7044 34754 7100
rect 34754 7044 34810 7100
rect 34810 7044 34814 7100
rect 34750 7040 34814 7044
rect 34830 7100 34894 7104
rect 34830 7044 34834 7100
rect 34834 7044 34890 7100
rect 34890 7044 34894 7100
rect 34830 7040 34894 7044
rect 34910 7100 34974 7104
rect 34910 7044 34914 7100
rect 34914 7044 34970 7100
rect 34970 7044 34974 7100
rect 34910 7040 34974 7044
rect 34990 7100 35054 7104
rect 34990 7044 34994 7100
rect 34994 7044 35050 7100
rect 35050 7044 35054 7100
rect 34990 7040 35054 7044
rect 102347 7100 102411 7104
rect 102347 7044 102351 7100
rect 102351 7044 102407 7100
rect 102407 7044 102411 7100
rect 102347 7040 102411 7044
rect 102427 7100 102491 7104
rect 102427 7044 102431 7100
rect 102431 7044 102487 7100
rect 102487 7044 102491 7100
rect 102427 7040 102491 7044
rect 102507 7100 102571 7104
rect 102507 7044 102511 7100
rect 102511 7044 102567 7100
rect 102567 7044 102571 7100
rect 102507 7040 102571 7044
rect 102587 7100 102651 7104
rect 102587 7044 102591 7100
rect 102591 7044 102647 7100
rect 102647 7044 102651 7100
rect 102587 7040 102651 7044
rect 169944 7100 170008 7104
rect 169944 7044 169948 7100
rect 169948 7044 170004 7100
rect 170004 7044 170008 7100
rect 169944 7040 170008 7044
rect 170024 7100 170088 7104
rect 170024 7044 170028 7100
rect 170028 7044 170084 7100
rect 170084 7044 170088 7100
rect 170024 7040 170088 7044
rect 170104 7100 170168 7104
rect 170104 7044 170108 7100
rect 170108 7044 170164 7100
rect 170164 7044 170168 7100
rect 170104 7040 170168 7044
rect 170184 7100 170248 7104
rect 170184 7044 170188 7100
rect 170188 7044 170244 7100
rect 170244 7044 170248 7100
rect 170184 7040 170248 7044
rect 237541 7100 237605 7104
rect 237541 7044 237545 7100
rect 237545 7044 237601 7100
rect 237601 7044 237605 7100
rect 237541 7040 237605 7044
rect 237621 7100 237685 7104
rect 237621 7044 237625 7100
rect 237625 7044 237681 7100
rect 237681 7044 237685 7100
rect 237621 7040 237685 7044
rect 237701 7100 237765 7104
rect 237701 7044 237705 7100
rect 237705 7044 237761 7100
rect 237761 7044 237765 7100
rect 237701 7040 237765 7044
rect 237781 7100 237845 7104
rect 237781 7044 237785 7100
rect 237785 7044 237841 7100
rect 237841 7044 237845 7100
rect 237781 7040 237845 7044
rect 19196 6896 19260 6900
rect 19196 6840 19246 6896
rect 19246 6840 19260 6896
rect 19196 6836 19260 6840
rect 19932 6896 19996 6900
rect 19932 6840 19982 6896
rect 19982 6840 19996 6896
rect 19932 6836 19996 6840
rect 22876 6836 22940 6900
rect 23612 6836 23676 6900
rect 25084 6836 25148 6900
rect 212212 6836 212276 6900
rect 266124 6700 266188 6764
rect 267596 6700 267660 6764
rect 68548 6556 68612 6560
rect 68548 6500 68552 6556
rect 68552 6500 68608 6556
rect 68608 6500 68612 6556
rect 68548 6496 68612 6500
rect 68628 6556 68692 6560
rect 68628 6500 68632 6556
rect 68632 6500 68688 6556
rect 68688 6500 68692 6556
rect 68628 6496 68692 6500
rect 68708 6556 68772 6560
rect 68708 6500 68712 6556
rect 68712 6500 68768 6556
rect 68768 6500 68772 6556
rect 68708 6496 68772 6500
rect 68788 6556 68852 6560
rect 68788 6500 68792 6556
rect 68792 6500 68848 6556
rect 68848 6500 68852 6556
rect 68788 6496 68852 6500
rect 216628 6564 216692 6628
rect 136145 6556 136209 6560
rect 136145 6500 136149 6556
rect 136149 6500 136205 6556
rect 136205 6500 136209 6556
rect 136145 6496 136209 6500
rect 136225 6556 136289 6560
rect 136225 6500 136229 6556
rect 136229 6500 136285 6556
rect 136285 6500 136289 6556
rect 136225 6496 136289 6500
rect 136305 6556 136369 6560
rect 136305 6500 136309 6556
rect 136309 6500 136365 6556
rect 136365 6500 136369 6556
rect 136305 6496 136369 6500
rect 136385 6556 136449 6560
rect 136385 6500 136389 6556
rect 136389 6500 136445 6556
rect 136445 6500 136449 6556
rect 136385 6496 136449 6500
rect 203742 6556 203806 6560
rect 203742 6500 203746 6556
rect 203746 6500 203802 6556
rect 203802 6500 203806 6556
rect 203742 6496 203806 6500
rect 203822 6556 203886 6560
rect 203822 6500 203826 6556
rect 203826 6500 203882 6556
rect 203882 6500 203886 6556
rect 203822 6496 203886 6500
rect 203902 6556 203966 6560
rect 203902 6500 203906 6556
rect 203906 6500 203962 6556
rect 203962 6500 203966 6556
rect 203902 6496 203966 6500
rect 203982 6556 204046 6560
rect 203982 6500 203986 6556
rect 203986 6500 204042 6556
rect 204042 6500 204046 6556
rect 203982 6496 204046 6500
rect 271339 6556 271403 6560
rect 271339 6500 271343 6556
rect 271343 6500 271399 6556
rect 271399 6500 271403 6556
rect 271339 6496 271403 6500
rect 271419 6556 271483 6560
rect 271419 6500 271423 6556
rect 271423 6500 271479 6556
rect 271479 6500 271483 6556
rect 271419 6496 271483 6500
rect 271499 6556 271563 6560
rect 271499 6500 271503 6556
rect 271503 6500 271559 6556
rect 271559 6500 271563 6556
rect 271499 6496 271563 6500
rect 271579 6556 271643 6560
rect 271579 6500 271583 6556
rect 271583 6500 271639 6556
rect 271639 6500 271643 6556
rect 271579 6496 271643 6500
rect 262076 6156 262140 6220
rect 268148 6156 268212 6220
rect 34750 6012 34814 6016
rect 34750 5956 34754 6012
rect 34754 5956 34810 6012
rect 34810 5956 34814 6012
rect 34750 5952 34814 5956
rect 34830 6012 34894 6016
rect 34830 5956 34834 6012
rect 34834 5956 34890 6012
rect 34890 5956 34894 6012
rect 34830 5952 34894 5956
rect 34910 6012 34974 6016
rect 34910 5956 34914 6012
rect 34914 5956 34970 6012
rect 34970 5956 34974 6012
rect 34910 5952 34974 5956
rect 34990 6012 35054 6016
rect 34990 5956 34994 6012
rect 34994 5956 35050 6012
rect 35050 5956 35054 6012
rect 34990 5952 35054 5956
rect 102347 6012 102411 6016
rect 102347 5956 102351 6012
rect 102351 5956 102407 6012
rect 102407 5956 102411 6012
rect 102347 5952 102411 5956
rect 102427 6012 102491 6016
rect 102427 5956 102431 6012
rect 102431 5956 102487 6012
rect 102487 5956 102491 6012
rect 102427 5952 102491 5956
rect 102507 6012 102571 6016
rect 102507 5956 102511 6012
rect 102511 5956 102567 6012
rect 102567 5956 102571 6012
rect 102507 5952 102571 5956
rect 102587 6012 102651 6016
rect 102587 5956 102591 6012
rect 102591 5956 102647 6012
rect 102647 5956 102651 6012
rect 102587 5952 102651 5956
rect 169944 6012 170008 6016
rect 169944 5956 169948 6012
rect 169948 5956 170004 6012
rect 170004 5956 170008 6012
rect 169944 5952 170008 5956
rect 170024 6012 170088 6016
rect 170024 5956 170028 6012
rect 170028 5956 170084 6012
rect 170084 5956 170088 6012
rect 170024 5952 170088 5956
rect 170104 6012 170168 6016
rect 170104 5956 170108 6012
rect 170108 5956 170164 6012
rect 170164 5956 170168 6012
rect 170104 5952 170168 5956
rect 170184 6012 170248 6016
rect 170184 5956 170188 6012
rect 170188 5956 170244 6012
rect 170244 5956 170248 6012
rect 170184 5952 170248 5956
rect 237541 6012 237605 6016
rect 237541 5956 237545 6012
rect 237545 5956 237601 6012
rect 237601 5956 237605 6012
rect 237541 5952 237605 5956
rect 237621 6012 237685 6016
rect 237621 5956 237625 6012
rect 237625 5956 237681 6012
rect 237681 5956 237685 6012
rect 237621 5952 237685 5956
rect 237701 6012 237765 6016
rect 237701 5956 237705 6012
rect 237705 5956 237761 6012
rect 237761 5956 237765 6012
rect 237701 5952 237765 5956
rect 237781 6012 237845 6016
rect 237781 5956 237785 6012
rect 237785 5956 237841 6012
rect 237841 5956 237845 6012
rect 237781 5952 237845 5956
rect 271092 5748 271156 5812
rect 230612 5476 230676 5540
rect 266860 5672 266924 5676
rect 266860 5616 266910 5672
rect 266910 5616 266924 5672
rect 266860 5612 266924 5616
rect 267780 5672 267844 5676
rect 267780 5616 267794 5672
rect 267794 5616 267844 5672
rect 267780 5612 267844 5616
rect 268332 5612 268396 5676
rect 269252 5612 269316 5676
rect 269804 5612 269868 5676
rect 270540 5672 270604 5676
rect 270540 5616 270554 5672
rect 270554 5616 270604 5672
rect 270540 5612 270604 5616
rect 68548 5468 68612 5472
rect 68548 5412 68552 5468
rect 68552 5412 68608 5468
rect 68608 5412 68612 5468
rect 68548 5408 68612 5412
rect 68628 5468 68692 5472
rect 68628 5412 68632 5468
rect 68632 5412 68688 5468
rect 68688 5412 68692 5468
rect 68628 5408 68692 5412
rect 68708 5468 68772 5472
rect 68708 5412 68712 5468
rect 68712 5412 68768 5468
rect 68768 5412 68772 5468
rect 68708 5408 68772 5412
rect 68788 5468 68852 5472
rect 68788 5412 68792 5468
rect 68792 5412 68848 5468
rect 68848 5412 68852 5468
rect 68788 5408 68852 5412
rect 136145 5468 136209 5472
rect 136145 5412 136149 5468
rect 136149 5412 136205 5468
rect 136205 5412 136209 5468
rect 136145 5408 136209 5412
rect 136225 5468 136289 5472
rect 136225 5412 136229 5468
rect 136229 5412 136285 5468
rect 136285 5412 136289 5468
rect 136225 5408 136289 5412
rect 136305 5468 136369 5472
rect 136305 5412 136309 5468
rect 136309 5412 136365 5468
rect 136365 5412 136369 5468
rect 136305 5408 136369 5412
rect 136385 5468 136449 5472
rect 136385 5412 136389 5468
rect 136389 5412 136445 5468
rect 136445 5412 136449 5468
rect 136385 5408 136449 5412
rect 203742 5468 203806 5472
rect 203742 5412 203746 5468
rect 203746 5412 203802 5468
rect 203802 5412 203806 5468
rect 203742 5408 203806 5412
rect 203822 5468 203886 5472
rect 203822 5412 203826 5468
rect 203826 5412 203882 5468
rect 203882 5412 203886 5468
rect 203822 5408 203886 5412
rect 203902 5468 203966 5472
rect 203902 5412 203906 5468
rect 203906 5412 203962 5468
rect 203962 5412 203966 5468
rect 203902 5408 203966 5412
rect 203982 5468 204046 5472
rect 203982 5412 203986 5468
rect 203986 5412 204042 5468
rect 204042 5412 204046 5468
rect 203982 5408 204046 5412
rect 271339 5468 271403 5472
rect 271339 5412 271343 5468
rect 271343 5412 271399 5468
rect 271399 5412 271403 5468
rect 271339 5408 271403 5412
rect 271419 5468 271483 5472
rect 271419 5412 271423 5468
rect 271423 5412 271479 5468
rect 271479 5412 271483 5468
rect 271419 5408 271483 5412
rect 271499 5468 271563 5472
rect 271499 5412 271503 5468
rect 271503 5412 271559 5468
rect 271559 5412 271563 5468
rect 271499 5408 271563 5412
rect 271579 5468 271643 5472
rect 271579 5412 271583 5468
rect 271583 5412 271639 5468
rect 271639 5412 271643 5468
rect 271579 5408 271643 5412
rect 263180 5264 263244 5268
rect 263180 5208 263230 5264
rect 263230 5208 263244 5264
rect 263180 5204 263244 5208
rect 230612 5068 230676 5132
rect 34750 4924 34814 4928
rect 34750 4868 34754 4924
rect 34754 4868 34810 4924
rect 34810 4868 34814 4924
rect 34750 4864 34814 4868
rect 34830 4924 34894 4928
rect 34830 4868 34834 4924
rect 34834 4868 34890 4924
rect 34890 4868 34894 4924
rect 34830 4864 34894 4868
rect 34910 4924 34974 4928
rect 34910 4868 34914 4924
rect 34914 4868 34970 4924
rect 34970 4868 34974 4924
rect 34910 4864 34974 4868
rect 34990 4924 35054 4928
rect 34990 4868 34994 4924
rect 34994 4868 35050 4924
rect 35050 4868 35054 4924
rect 34990 4864 35054 4868
rect 102347 4924 102411 4928
rect 102347 4868 102351 4924
rect 102351 4868 102407 4924
rect 102407 4868 102411 4924
rect 102347 4864 102411 4868
rect 102427 4924 102491 4928
rect 102427 4868 102431 4924
rect 102431 4868 102487 4924
rect 102487 4868 102491 4924
rect 102427 4864 102491 4868
rect 102507 4924 102571 4928
rect 102507 4868 102511 4924
rect 102511 4868 102567 4924
rect 102567 4868 102571 4924
rect 102507 4864 102571 4868
rect 102587 4924 102651 4928
rect 102587 4868 102591 4924
rect 102591 4868 102647 4924
rect 102647 4868 102651 4924
rect 102587 4864 102651 4868
rect 169944 4924 170008 4928
rect 169944 4868 169948 4924
rect 169948 4868 170004 4924
rect 170004 4868 170008 4924
rect 169944 4864 170008 4868
rect 170024 4924 170088 4928
rect 170024 4868 170028 4924
rect 170028 4868 170084 4924
rect 170084 4868 170088 4924
rect 170024 4864 170088 4868
rect 170104 4924 170168 4928
rect 170104 4868 170108 4924
rect 170108 4868 170164 4924
rect 170164 4868 170168 4924
rect 170104 4864 170168 4868
rect 170184 4924 170248 4928
rect 170184 4868 170188 4924
rect 170188 4868 170244 4924
rect 170244 4868 170248 4924
rect 170184 4864 170248 4868
rect 237541 4924 237605 4928
rect 237541 4868 237545 4924
rect 237545 4868 237601 4924
rect 237601 4868 237605 4924
rect 237541 4864 237605 4868
rect 237621 4924 237685 4928
rect 237621 4868 237625 4924
rect 237625 4868 237681 4924
rect 237681 4868 237685 4924
rect 237621 4864 237685 4868
rect 237701 4924 237765 4928
rect 237701 4868 237705 4924
rect 237705 4868 237761 4924
rect 237761 4868 237765 4924
rect 237701 4864 237765 4868
rect 237781 4924 237845 4928
rect 237781 4868 237785 4924
rect 237785 4868 237841 4924
rect 237841 4868 237845 4924
rect 237781 4864 237845 4868
rect 68548 4380 68612 4384
rect 68548 4324 68552 4380
rect 68552 4324 68608 4380
rect 68608 4324 68612 4380
rect 68548 4320 68612 4324
rect 68628 4380 68692 4384
rect 68628 4324 68632 4380
rect 68632 4324 68688 4380
rect 68688 4324 68692 4380
rect 68628 4320 68692 4324
rect 68708 4380 68772 4384
rect 68708 4324 68712 4380
rect 68712 4324 68768 4380
rect 68768 4324 68772 4380
rect 68708 4320 68772 4324
rect 68788 4380 68852 4384
rect 68788 4324 68792 4380
rect 68792 4324 68848 4380
rect 68848 4324 68852 4380
rect 68788 4320 68852 4324
rect 136145 4380 136209 4384
rect 136145 4324 136149 4380
rect 136149 4324 136205 4380
rect 136205 4324 136209 4380
rect 136145 4320 136209 4324
rect 136225 4380 136289 4384
rect 136225 4324 136229 4380
rect 136229 4324 136285 4380
rect 136285 4324 136289 4380
rect 136225 4320 136289 4324
rect 136305 4380 136369 4384
rect 136305 4324 136309 4380
rect 136309 4324 136365 4380
rect 136365 4324 136369 4380
rect 136305 4320 136369 4324
rect 136385 4380 136449 4384
rect 136385 4324 136389 4380
rect 136389 4324 136445 4380
rect 136445 4324 136449 4380
rect 136385 4320 136449 4324
rect 203742 4380 203806 4384
rect 203742 4324 203746 4380
rect 203746 4324 203802 4380
rect 203802 4324 203806 4380
rect 203742 4320 203806 4324
rect 203822 4380 203886 4384
rect 203822 4324 203826 4380
rect 203826 4324 203882 4380
rect 203882 4324 203886 4380
rect 203822 4320 203886 4324
rect 203902 4380 203966 4384
rect 203902 4324 203906 4380
rect 203906 4324 203962 4380
rect 203962 4324 203966 4380
rect 203902 4320 203966 4324
rect 203982 4380 204046 4384
rect 203982 4324 203986 4380
rect 203986 4324 204042 4380
rect 204042 4324 204046 4380
rect 203982 4320 204046 4324
rect 271339 4380 271403 4384
rect 271339 4324 271343 4380
rect 271343 4324 271399 4380
rect 271399 4324 271403 4380
rect 271339 4320 271403 4324
rect 271419 4380 271483 4384
rect 271419 4324 271423 4380
rect 271423 4324 271479 4380
rect 271479 4324 271483 4380
rect 271419 4320 271483 4324
rect 271499 4380 271563 4384
rect 271499 4324 271503 4380
rect 271503 4324 271559 4380
rect 271559 4324 271563 4380
rect 271499 4320 271563 4324
rect 271579 4380 271643 4384
rect 271579 4324 271583 4380
rect 271583 4324 271639 4380
rect 271639 4324 271643 4380
rect 271579 4320 271643 4324
rect 34750 3836 34814 3840
rect 34750 3780 34754 3836
rect 34754 3780 34810 3836
rect 34810 3780 34814 3836
rect 34750 3776 34814 3780
rect 34830 3836 34894 3840
rect 34830 3780 34834 3836
rect 34834 3780 34890 3836
rect 34890 3780 34894 3836
rect 34830 3776 34894 3780
rect 34910 3836 34974 3840
rect 34910 3780 34914 3836
rect 34914 3780 34970 3836
rect 34970 3780 34974 3836
rect 34910 3776 34974 3780
rect 34990 3836 35054 3840
rect 34990 3780 34994 3836
rect 34994 3780 35050 3836
rect 35050 3780 35054 3836
rect 34990 3776 35054 3780
rect 102347 3836 102411 3840
rect 102347 3780 102351 3836
rect 102351 3780 102407 3836
rect 102407 3780 102411 3836
rect 102347 3776 102411 3780
rect 102427 3836 102491 3840
rect 102427 3780 102431 3836
rect 102431 3780 102487 3836
rect 102487 3780 102491 3836
rect 102427 3776 102491 3780
rect 102507 3836 102571 3840
rect 102507 3780 102511 3836
rect 102511 3780 102567 3836
rect 102567 3780 102571 3836
rect 102507 3776 102571 3780
rect 102587 3836 102651 3840
rect 102587 3780 102591 3836
rect 102591 3780 102647 3836
rect 102647 3780 102651 3836
rect 102587 3776 102651 3780
rect 169944 3836 170008 3840
rect 169944 3780 169948 3836
rect 169948 3780 170004 3836
rect 170004 3780 170008 3836
rect 169944 3776 170008 3780
rect 170024 3836 170088 3840
rect 170024 3780 170028 3836
rect 170028 3780 170084 3836
rect 170084 3780 170088 3836
rect 170024 3776 170088 3780
rect 170104 3836 170168 3840
rect 170104 3780 170108 3836
rect 170108 3780 170164 3836
rect 170164 3780 170168 3836
rect 170104 3776 170168 3780
rect 170184 3836 170248 3840
rect 170184 3780 170188 3836
rect 170188 3780 170244 3836
rect 170244 3780 170248 3836
rect 170184 3776 170248 3780
rect 237541 3836 237605 3840
rect 237541 3780 237545 3836
rect 237545 3780 237601 3836
rect 237601 3780 237605 3836
rect 237541 3776 237605 3780
rect 237621 3836 237685 3840
rect 237621 3780 237625 3836
rect 237625 3780 237681 3836
rect 237681 3780 237685 3836
rect 237621 3776 237685 3780
rect 237701 3836 237765 3840
rect 237701 3780 237705 3836
rect 237705 3780 237761 3836
rect 237761 3780 237765 3836
rect 237701 3776 237765 3780
rect 237781 3836 237845 3840
rect 237781 3780 237785 3836
rect 237785 3780 237841 3836
rect 237841 3780 237845 3836
rect 237781 3776 237845 3780
rect 215340 3708 215404 3772
rect 267596 3708 267660 3772
rect 24348 3300 24412 3364
rect 68548 3292 68612 3296
rect 68548 3236 68552 3292
rect 68552 3236 68608 3292
rect 68608 3236 68612 3292
rect 68548 3232 68612 3236
rect 68628 3292 68692 3296
rect 68628 3236 68632 3292
rect 68632 3236 68688 3292
rect 68688 3236 68692 3292
rect 68628 3232 68692 3236
rect 68708 3292 68772 3296
rect 68708 3236 68712 3292
rect 68712 3236 68768 3292
rect 68768 3236 68772 3292
rect 68708 3232 68772 3236
rect 68788 3292 68852 3296
rect 68788 3236 68792 3292
rect 68792 3236 68848 3292
rect 68848 3236 68852 3292
rect 68788 3232 68852 3236
rect 136145 3292 136209 3296
rect 136145 3236 136149 3292
rect 136149 3236 136205 3292
rect 136205 3236 136209 3292
rect 136145 3232 136209 3236
rect 136225 3292 136289 3296
rect 136225 3236 136229 3292
rect 136229 3236 136285 3292
rect 136285 3236 136289 3292
rect 136225 3232 136289 3236
rect 136305 3292 136369 3296
rect 136305 3236 136309 3292
rect 136309 3236 136365 3292
rect 136365 3236 136369 3292
rect 136305 3232 136369 3236
rect 136385 3292 136449 3296
rect 136385 3236 136389 3292
rect 136389 3236 136445 3292
rect 136445 3236 136449 3292
rect 136385 3232 136449 3236
rect 203742 3292 203806 3296
rect 203742 3236 203746 3292
rect 203746 3236 203802 3292
rect 203802 3236 203806 3292
rect 203742 3232 203806 3236
rect 203822 3292 203886 3296
rect 203822 3236 203826 3292
rect 203826 3236 203882 3292
rect 203882 3236 203886 3292
rect 203822 3232 203886 3236
rect 203902 3292 203966 3296
rect 203902 3236 203906 3292
rect 203906 3236 203962 3292
rect 203962 3236 203966 3292
rect 203902 3232 203966 3236
rect 203982 3292 204046 3296
rect 203982 3236 203986 3292
rect 203986 3236 204042 3292
rect 204042 3236 204046 3292
rect 203982 3232 204046 3236
rect 271339 3292 271403 3296
rect 271339 3236 271343 3292
rect 271343 3236 271399 3292
rect 271399 3236 271403 3292
rect 271339 3232 271403 3236
rect 271419 3292 271483 3296
rect 271419 3236 271423 3292
rect 271423 3236 271479 3292
rect 271479 3236 271483 3292
rect 271419 3232 271483 3236
rect 271499 3292 271563 3296
rect 271499 3236 271503 3292
rect 271503 3236 271559 3292
rect 271559 3236 271563 3292
rect 271499 3232 271563 3236
rect 271579 3292 271643 3296
rect 271579 3236 271583 3292
rect 271583 3236 271639 3292
rect 271639 3236 271643 3292
rect 271579 3232 271643 3236
rect 267964 3164 268028 3228
rect 19196 2952 19260 2956
rect 19196 2896 19246 2952
rect 19246 2896 19260 2952
rect 19196 2892 19260 2896
rect 22876 2952 22940 2956
rect 22876 2896 22926 2952
rect 22926 2896 22940 2952
rect 22876 2892 22940 2896
rect 19932 2816 19996 2820
rect 19932 2760 19982 2816
rect 19982 2760 19996 2816
rect 19932 2756 19996 2760
rect 22140 2756 22204 2820
rect 25084 2756 25148 2820
rect 60044 2756 60108 2820
rect 157196 2816 157260 2820
rect 157196 2760 157246 2816
rect 157246 2760 157260 2816
rect 157196 2756 157260 2760
rect 159404 2756 159468 2820
rect 189948 2756 190012 2820
rect 191420 2756 191484 2820
rect 202460 2756 202524 2820
rect 223252 2816 223316 2820
rect 223252 2760 223302 2816
rect 223302 2760 223316 2816
rect 223252 2756 223316 2760
rect 224724 2756 224788 2820
rect 226196 2816 226260 2820
rect 226196 2760 226246 2816
rect 226246 2760 226260 2816
rect 226196 2756 226260 2760
rect 235764 2756 235828 2820
rect 258028 2816 258092 2820
rect 258028 2760 258078 2816
rect 258078 2760 258092 2816
rect 258028 2756 258092 2760
rect 270540 2816 270604 2820
rect 270540 2760 270554 2816
rect 270554 2760 270604 2816
rect 270540 2756 270604 2760
rect 34750 2748 34814 2752
rect 34750 2692 34754 2748
rect 34754 2692 34810 2748
rect 34810 2692 34814 2748
rect 34750 2688 34814 2692
rect 34830 2748 34894 2752
rect 34830 2692 34834 2748
rect 34834 2692 34890 2748
rect 34890 2692 34894 2748
rect 34830 2688 34894 2692
rect 34910 2748 34974 2752
rect 34910 2692 34914 2748
rect 34914 2692 34970 2748
rect 34970 2692 34974 2748
rect 34910 2688 34974 2692
rect 34990 2748 35054 2752
rect 34990 2692 34994 2748
rect 34994 2692 35050 2748
rect 35050 2692 35054 2748
rect 34990 2688 35054 2692
rect 102347 2748 102411 2752
rect 102347 2692 102351 2748
rect 102351 2692 102407 2748
rect 102407 2692 102411 2748
rect 102347 2688 102411 2692
rect 102427 2748 102491 2752
rect 102427 2692 102431 2748
rect 102431 2692 102487 2748
rect 102487 2692 102491 2748
rect 102427 2688 102491 2692
rect 102507 2748 102571 2752
rect 102507 2692 102511 2748
rect 102511 2692 102567 2748
rect 102567 2692 102571 2748
rect 102507 2688 102571 2692
rect 102587 2748 102651 2752
rect 102587 2692 102591 2748
rect 102591 2692 102647 2748
rect 102647 2692 102651 2748
rect 102587 2688 102651 2692
rect 169944 2748 170008 2752
rect 169944 2692 169948 2748
rect 169948 2692 170004 2748
rect 170004 2692 170008 2748
rect 169944 2688 170008 2692
rect 170024 2748 170088 2752
rect 170024 2692 170028 2748
rect 170028 2692 170084 2748
rect 170084 2692 170088 2748
rect 170024 2688 170088 2692
rect 170104 2748 170168 2752
rect 170104 2692 170108 2748
rect 170108 2692 170164 2748
rect 170164 2692 170168 2748
rect 170104 2688 170168 2692
rect 170184 2748 170248 2752
rect 170184 2692 170188 2748
rect 170188 2692 170244 2748
rect 170244 2692 170248 2748
rect 170184 2688 170248 2692
rect 237541 2748 237605 2752
rect 237541 2692 237545 2748
rect 237545 2692 237601 2748
rect 237601 2692 237605 2748
rect 237541 2688 237605 2692
rect 237621 2748 237685 2752
rect 237621 2692 237625 2748
rect 237625 2692 237681 2748
rect 237681 2692 237685 2748
rect 237621 2688 237685 2692
rect 237701 2748 237765 2752
rect 237701 2692 237705 2748
rect 237705 2692 237761 2748
rect 237761 2692 237765 2748
rect 237701 2688 237765 2692
rect 237781 2748 237845 2752
rect 237781 2692 237785 2748
rect 237785 2692 237841 2748
rect 237841 2692 237845 2748
rect 237781 2688 237845 2692
rect 266492 2620 266556 2684
rect 223620 2484 223684 2548
rect 267964 2484 268028 2548
rect 216628 2348 216692 2412
rect 224172 2212 224236 2276
rect 68548 2204 68612 2208
rect 68548 2148 68552 2204
rect 68552 2148 68608 2204
rect 68608 2148 68612 2204
rect 68548 2144 68612 2148
rect 68628 2204 68692 2208
rect 68628 2148 68632 2204
rect 68632 2148 68688 2204
rect 68688 2148 68692 2204
rect 68628 2144 68692 2148
rect 68708 2204 68772 2208
rect 68708 2148 68712 2204
rect 68712 2148 68768 2204
rect 68768 2148 68772 2204
rect 68708 2144 68772 2148
rect 68788 2204 68852 2208
rect 68788 2148 68792 2204
rect 68792 2148 68848 2204
rect 68848 2148 68852 2204
rect 68788 2144 68852 2148
rect 136145 2204 136209 2208
rect 136145 2148 136149 2204
rect 136149 2148 136205 2204
rect 136205 2148 136209 2204
rect 136145 2144 136209 2148
rect 136225 2204 136289 2208
rect 136225 2148 136229 2204
rect 136229 2148 136285 2204
rect 136285 2148 136289 2204
rect 136225 2144 136289 2148
rect 136305 2204 136369 2208
rect 136305 2148 136309 2204
rect 136309 2148 136365 2204
rect 136365 2148 136369 2204
rect 136305 2144 136369 2148
rect 136385 2204 136449 2208
rect 136385 2148 136389 2204
rect 136389 2148 136445 2204
rect 136445 2148 136449 2204
rect 136385 2144 136449 2148
rect 203742 2204 203806 2208
rect 203742 2148 203746 2204
rect 203746 2148 203802 2204
rect 203802 2148 203806 2204
rect 203742 2144 203806 2148
rect 203822 2204 203886 2208
rect 203822 2148 203826 2204
rect 203826 2148 203882 2204
rect 203882 2148 203886 2204
rect 203822 2144 203886 2148
rect 203902 2204 203966 2208
rect 203902 2148 203906 2204
rect 203906 2148 203962 2204
rect 203962 2148 203966 2204
rect 203902 2144 203966 2148
rect 203982 2204 204046 2208
rect 203982 2148 203986 2204
rect 203986 2148 204042 2204
rect 204042 2148 204046 2204
rect 203982 2144 204046 2148
rect 271339 2204 271403 2208
rect 271339 2148 271343 2204
rect 271343 2148 271399 2204
rect 271399 2148 271403 2204
rect 271339 2144 271403 2148
rect 271419 2204 271483 2208
rect 271419 2148 271423 2204
rect 271423 2148 271479 2204
rect 271479 2148 271483 2204
rect 271419 2144 271483 2148
rect 271499 2204 271563 2208
rect 271499 2148 271503 2204
rect 271503 2148 271559 2204
rect 271559 2148 271563 2204
rect 271499 2144 271563 2148
rect 271579 2204 271643 2208
rect 271579 2148 271583 2204
rect 271583 2148 271639 2204
rect 271639 2148 271643 2204
rect 271579 2144 271643 2148
rect 21404 1668 21468 1732
rect 215340 1668 215404 1732
rect 267412 1668 267476 1732
rect 34750 1660 34814 1664
rect 34750 1604 34754 1660
rect 34754 1604 34810 1660
rect 34810 1604 34814 1660
rect 34750 1600 34814 1604
rect 34830 1660 34894 1664
rect 34830 1604 34834 1660
rect 34834 1604 34890 1660
rect 34890 1604 34894 1660
rect 34830 1600 34894 1604
rect 34910 1660 34974 1664
rect 34910 1604 34914 1660
rect 34914 1604 34970 1660
rect 34970 1604 34974 1660
rect 34910 1600 34974 1604
rect 34990 1660 35054 1664
rect 34990 1604 34994 1660
rect 34994 1604 35050 1660
rect 35050 1604 35054 1660
rect 34990 1600 35054 1604
rect 102347 1660 102411 1664
rect 102347 1604 102351 1660
rect 102351 1604 102407 1660
rect 102407 1604 102411 1660
rect 102347 1600 102411 1604
rect 102427 1660 102491 1664
rect 102427 1604 102431 1660
rect 102431 1604 102487 1660
rect 102487 1604 102491 1660
rect 102427 1600 102491 1604
rect 102507 1660 102571 1664
rect 102507 1604 102511 1660
rect 102511 1604 102567 1660
rect 102567 1604 102571 1660
rect 102507 1600 102571 1604
rect 102587 1660 102651 1664
rect 102587 1604 102591 1660
rect 102591 1604 102647 1660
rect 102647 1604 102651 1660
rect 102587 1600 102651 1604
rect 169944 1660 170008 1664
rect 169944 1604 169948 1660
rect 169948 1604 170004 1660
rect 170004 1604 170008 1660
rect 169944 1600 170008 1604
rect 170024 1660 170088 1664
rect 170024 1604 170028 1660
rect 170028 1604 170084 1660
rect 170084 1604 170088 1660
rect 170024 1600 170088 1604
rect 170104 1660 170168 1664
rect 170104 1604 170108 1660
rect 170108 1604 170164 1660
rect 170164 1604 170168 1660
rect 170104 1600 170168 1604
rect 170184 1660 170248 1664
rect 170184 1604 170188 1660
rect 170188 1604 170244 1660
rect 170244 1604 170248 1660
rect 170184 1600 170248 1604
rect 237541 1660 237605 1664
rect 237541 1604 237545 1660
rect 237545 1604 237601 1660
rect 237601 1604 237605 1660
rect 237541 1600 237605 1604
rect 237621 1660 237685 1664
rect 237621 1604 237625 1660
rect 237625 1604 237681 1660
rect 237681 1604 237685 1660
rect 237621 1600 237685 1604
rect 237701 1660 237765 1664
rect 237701 1604 237705 1660
rect 237705 1604 237761 1660
rect 237761 1604 237765 1660
rect 237701 1600 237765 1604
rect 237781 1660 237845 1664
rect 237781 1604 237785 1660
rect 237785 1604 237841 1660
rect 237841 1604 237845 1660
rect 237781 1600 237845 1604
rect 59308 1592 59372 1596
rect 59308 1536 59358 1592
rect 59358 1536 59372 1592
rect 59308 1532 59372 1536
rect 80100 1592 80164 1596
rect 80100 1536 80114 1592
rect 80114 1536 80164 1592
rect 80100 1532 80164 1536
rect 81572 1532 81636 1596
rect 83044 1592 83108 1596
rect 83044 1536 83058 1592
rect 83058 1536 83108 1592
rect 83044 1532 83108 1536
rect 83780 1592 83844 1596
rect 83780 1536 83794 1592
rect 83794 1536 83844 1592
rect 83780 1532 83844 1536
rect 99236 1532 99300 1596
rect 796 1456 860 1460
rect 796 1400 846 1456
rect 846 1400 860 1456
rect 796 1396 860 1400
rect 16252 1396 16316 1460
rect 20668 1396 20732 1460
rect 32444 1396 32508 1460
rect 53972 1456 54036 1460
rect 53972 1400 53986 1456
rect 53986 1400 54036 1456
rect 53972 1396 54036 1400
rect 117268 1456 117332 1460
rect 117268 1400 117318 1456
rect 117318 1400 117332 1456
rect 117268 1396 117332 1400
rect 128308 1456 128372 1460
rect 128308 1400 128358 1456
rect 128358 1400 128372 1456
rect 128308 1396 128372 1400
rect 134932 1396 134996 1460
rect 137324 1396 137388 1460
rect 144684 1396 144748 1460
rect 155724 1396 155788 1460
rect 156460 1396 156524 1460
rect 157932 1456 157996 1460
rect 157932 1400 157946 1456
rect 157946 1400 157996 1456
rect 157932 1396 157996 1400
rect 163820 1396 163884 1460
rect 168236 1396 168300 1460
rect 186268 1456 186332 1460
rect 186268 1400 186318 1456
rect 186318 1400 186332 1456
rect 186268 1396 186332 1400
rect 194364 1396 194428 1460
rect 195836 1396 195900 1460
rect 201724 1532 201788 1596
rect 216628 1456 216692 1460
rect 216628 1400 216678 1456
rect 216678 1400 216692 1456
rect 216628 1396 216692 1400
rect 220308 1396 220372 1460
rect 223988 1456 224052 1460
rect 223988 1400 224038 1456
rect 224038 1400 224052 1456
rect 223988 1396 224052 1400
rect 225460 1396 225524 1460
rect 237236 1456 237300 1460
rect 237236 1400 237286 1456
rect 237286 1400 237300 1456
rect 237236 1396 237300 1400
rect 242756 1396 242820 1460
rect 244044 1396 244108 1460
rect 247908 1396 247972 1460
rect 249380 1396 249444 1460
rect 250852 1396 250916 1460
rect 264836 1396 264900 1460
rect 1532 1320 1596 1324
rect 1532 1264 1582 1320
rect 1582 1264 1596 1320
rect 1532 1260 1596 1264
rect 25820 1260 25884 1324
rect 26556 1260 26620 1324
rect 27292 1260 27356 1324
rect 71268 1320 71332 1324
rect 71268 1264 71318 1320
rect 71318 1264 71332 1320
rect 71268 1260 71332 1264
rect 73476 1320 73540 1324
rect 73476 1264 73526 1320
rect 73526 1264 73540 1320
rect 73476 1260 73540 1264
rect 76420 1320 76484 1324
rect 76420 1264 76470 1320
rect 76470 1264 76484 1320
rect 76420 1260 76484 1264
rect 77892 1320 77956 1324
rect 77892 1264 77942 1320
rect 77942 1264 77956 1320
rect 77892 1260 77956 1264
rect 79364 1320 79428 1324
rect 79364 1264 79414 1320
rect 79414 1264 79428 1320
rect 79364 1260 79428 1264
rect 82308 1260 82372 1324
rect 87460 1320 87524 1324
rect 87460 1264 87510 1320
rect 87510 1264 87524 1320
rect 87460 1260 87524 1264
rect 88932 1260 88996 1324
rect 140268 1260 140332 1324
rect 154988 1260 155052 1324
rect 176700 1320 176764 1324
rect 176700 1264 176714 1320
rect 176714 1264 176764 1320
rect 176700 1260 176764 1264
rect 179644 1320 179708 1324
rect 179644 1264 179658 1320
rect 179658 1264 179708 1320
rect 179644 1260 179708 1264
rect 181852 1320 181916 1324
rect 181852 1264 181902 1320
rect 181902 1264 181916 1320
rect 181852 1260 181916 1264
rect 187004 1320 187068 1324
rect 187004 1264 187018 1320
rect 187018 1264 187068 1320
rect 187004 1260 187068 1264
rect 199516 1260 199580 1324
rect 210740 1260 210804 1324
rect 222516 1260 222580 1324
rect 226932 1260 226996 1324
rect 227668 1260 227732 1324
rect 2268 1048 2332 1052
rect 2268 992 2318 1048
rect 2318 992 2332 1048
rect 2268 988 2332 992
rect 4476 1048 4540 1052
rect 4476 992 4526 1048
rect 4526 992 4540 1048
rect 4476 988 4540 992
rect 6684 988 6748 1052
rect 14044 1048 14108 1052
rect 14044 992 14094 1048
rect 14094 992 14108 1048
rect 14044 988 14108 992
rect 68548 1116 68612 1120
rect 68548 1060 68552 1116
rect 68552 1060 68608 1116
rect 68608 1060 68612 1116
rect 68548 1056 68612 1060
rect 68628 1116 68692 1120
rect 68628 1060 68632 1116
rect 68632 1060 68688 1116
rect 68688 1060 68692 1116
rect 68628 1056 68692 1060
rect 68708 1116 68772 1120
rect 68708 1060 68712 1116
rect 68712 1060 68768 1116
rect 68768 1060 68772 1116
rect 68708 1056 68772 1060
rect 68788 1116 68852 1120
rect 68788 1060 68792 1116
rect 68792 1060 68848 1116
rect 68848 1060 68852 1116
rect 68788 1056 68852 1060
rect 70532 1048 70596 1052
rect 70532 992 70582 1048
rect 70582 992 70596 1048
rect 70532 988 70596 992
rect 72004 1048 72068 1052
rect 72004 992 72054 1048
rect 72054 992 72068 1048
rect 72004 988 72068 992
rect 74212 1048 74276 1052
rect 74212 992 74262 1048
rect 74262 992 74276 1048
rect 74212 988 74276 992
rect 75684 1048 75748 1052
rect 75684 992 75734 1048
rect 75734 992 75748 1048
rect 75684 988 75748 992
rect 77156 1048 77220 1052
rect 77156 992 77206 1048
rect 77206 992 77220 1048
rect 77156 988 77220 992
rect 85988 988 86052 1052
rect 88196 1124 88260 1188
rect 94084 1124 94148 1188
rect 94820 1124 94884 1188
rect 95556 1124 95620 1188
rect 96292 1124 96356 1188
rect 160140 1124 160204 1188
rect 161612 1124 161676 1188
rect 163084 1124 163148 1188
rect 165292 1184 165356 1188
rect 165292 1128 165342 1184
rect 165342 1128 165356 1184
rect 165292 1124 165356 1128
rect 166028 1184 166092 1188
rect 166028 1128 166078 1184
rect 166078 1128 166092 1184
rect 166028 1124 166092 1128
rect 166764 1184 166828 1188
rect 166764 1128 166814 1184
rect 166814 1128 166828 1184
rect 166764 1124 166828 1128
rect 136145 1116 136209 1120
rect 136145 1060 136149 1116
rect 136149 1060 136205 1116
rect 136205 1060 136209 1116
rect 136145 1056 136209 1060
rect 136225 1116 136289 1120
rect 136225 1060 136229 1116
rect 136229 1060 136285 1116
rect 136285 1060 136289 1116
rect 136225 1056 136289 1060
rect 136305 1116 136369 1120
rect 136305 1060 136309 1116
rect 136309 1060 136365 1116
rect 136365 1060 136369 1116
rect 136305 1056 136369 1060
rect 136385 1116 136449 1120
rect 136385 1060 136389 1116
rect 136389 1060 136445 1116
rect 136445 1060 136449 1116
rect 136385 1056 136449 1060
rect 142476 988 142540 1052
rect 149836 988 149900 1052
rect 190684 1124 190748 1188
rect 198044 1124 198108 1188
rect 200988 1124 201052 1188
rect 228404 1184 228468 1188
rect 228404 1128 228454 1184
rect 228454 1128 228468 1184
rect 228404 1124 228468 1128
rect 231348 1184 231412 1188
rect 231348 1128 231362 1184
rect 231362 1128 231412 1184
rect 231348 1124 231412 1128
rect 232084 1184 232148 1188
rect 232084 1128 232098 1184
rect 232098 1128 232148 1184
rect 232084 1124 232148 1128
rect 232820 1184 232884 1188
rect 232820 1128 232834 1184
rect 232834 1128 232884 1184
rect 232820 1124 232884 1128
rect 236500 1124 236564 1188
rect 247172 1124 247236 1188
rect 203742 1116 203806 1120
rect 203742 1060 203746 1116
rect 203746 1060 203802 1116
rect 203802 1060 203806 1116
rect 203742 1056 203806 1060
rect 203822 1116 203886 1120
rect 203822 1060 203826 1116
rect 203826 1060 203882 1116
rect 203882 1060 203886 1116
rect 203822 1056 203886 1060
rect 203902 1116 203966 1120
rect 203902 1060 203906 1116
rect 203906 1060 203962 1116
rect 203962 1060 203966 1116
rect 203902 1056 203966 1060
rect 203982 1116 204046 1120
rect 203982 1060 203986 1116
rect 203986 1060 204042 1116
rect 204042 1060 204046 1116
rect 203982 1056 204046 1060
rect 183324 1048 183388 1052
rect 183324 992 183338 1048
rect 183338 992 183388 1048
rect 183324 988 183388 992
rect 184796 1048 184860 1052
rect 184796 992 184810 1048
rect 184810 992 184860 1048
rect 184796 988 184860 992
rect 187740 988 187804 1052
rect 189212 988 189276 1052
rect 210004 988 210068 1052
rect 211476 988 211540 1052
rect 100708 852 100772 916
rect 3004 776 3068 780
rect 3004 720 3018 776
rect 3018 720 3068 776
rect 3004 716 3068 720
rect 5212 776 5276 780
rect 5212 720 5226 776
rect 5226 720 5276 776
rect 5212 716 5276 720
rect 5948 716 6012 780
rect 7420 716 7484 780
rect 8892 716 8956 780
rect 14780 776 14844 780
rect 14780 720 14830 776
rect 14830 720 14844 776
rect 14780 716 14844 720
rect 15516 716 15580 780
rect 69060 776 69124 780
rect 69060 720 69110 776
rect 69110 720 69124 776
rect 69060 716 69124 720
rect 69796 716 69860 780
rect 78628 776 78692 780
rect 78628 720 78642 776
rect 78642 720 78692 776
rect 78628 716 78692 720
rect 80836 716 80900 780
rect 84516 776 84580 780
rect 84516 720 84530 776
rect 84530 720 84580 776
rect 84516 716 84580 720
rect 85252 716 85316 780
rect 86724 776 86788 780
rect 86724 720 86774 776
rect 86774 720 86788 776
rect 86724 716 86788 720
rect 90404 716 90468 780
rect 91876 716 91940 780
rect 93348 716 93412 780
rect 97764 716 97828 780
rect 98500 776 98564 780
rect 171548 852 171612 916
rect 172284 912 172348 916
rect 172284 856 172298 912
rect 172298 856 172348 912
rect 172284 852 172348 856
rect 173020 912 173084 916
rect 173020 856 173034 912
rect 173034 856 173084 912
rect 173020 852 173084 856
rect 173756 912 173820 916
rect 173756 856 173806 912
rect 173806 856 173820 912
rect 173756 852 173820 856
rect 174492 912 174556 916
rect 174492 856 174506 912
rect 174506 856 174556 912
rect 174492 852 174556 856
rect 175228 912 175292 916
rect 175228 856 175242 912
rect 175242 856 175292 912
rect 175228 852 175292 856
rect 175964 852 176028 916
rect 177436 852 177500 916
rect 178172 852 178236 916
rect 178908 852 178972 916
rect 180380 852 180444 916
rect 181116 852 181180 916
rect 182588 912 182652 916
rect 182588 856 182602 912
rect 182602 856 182652 912
rect 182588 852 182652 856
rect 184060 852 184124 916
rect 185532 912 185596 916
rect 185532 856 185582 912
rect 185582 856 185596 912
rect 185532 852 185596 856
rect 188476 912 188540 916
rect 188476 856 188526 912
rect 188526 856 188540 912
rect 188476 852 188540 856
rect 192156 852 192220 916
rect 192892 912 192956 916
rect 192892 856 192942 912
rect 192942 856 192956 912
rect 192892 852 192956 856
rect 193628 912 193692 916
rect 193628 856 193678 912
rect 193678 856 193692 912
rect 193628 852 193692 856
rect 195100 852 195164 916
rect 196572 912 196636 916
rect 196572 856 196622 912
rect 196622 856 196636 912
rect 196572 852 196636 856
rect 197308 912 197372 916
rect 197308 856 197322 912
rect 197322 856 197372 912
rect 197308 852 197372 856
rect 198780 852 198844 916
rect 200252 852 200316 916
rect 203196 852 203260 916
rect 205772 912 205836 916
rect 205772 856 205822 912
rect 205822 856 205836 912
rect 205772 852 205836 856
rect 206324 852 206388 916
rect 207060 852 207124 916
rect 207796 852 207860 916
rect 208532 852 208596 916
rect 209268 852 209332 916
rect 212212 912 212276 916
rect 212212 856 212262 912
rect 212262 856 212276 912
rect 212212 852 212276 856
rect 212948 852 213012 916
rect 213684 912 213748 916
rect 213684 856 213734 912
rect 213734 856 213748 912
rect 213684 852 213748 856
rect 214420 912 214484 916
rect 214420 856 214470 912
rect 214470 856 214484 912
rect 214420 852 214484 856
rect 215156 912 215220 916
rect 215156 856 215170 912
rect 215170 856 215220 912
rect 215156 852 215220 856
rect 215892 852 215956 916
rect 217364 912 217428 916
rect 217364 856 217414 912
rect 217414 856 217428 912
rect 217364 852 217428 856
rect 218100 852 218164 916
rect 221044 852 221108 916
rect 98500 720 98514 776
rect 98514 720 98564 776
rect 98500 716 98564 720
rect 138796 776 138860 780
rect 138796 720 138846 776
rect 138846 720 138860 776
rect 3740 580 3804 644
rect 8156 640 8220 644
rect 8156 584 8206 640
rect 8206 584 8220 640
rect 8156 580 8220 584
rect 9628 640 9692 644
rect 9628 584 9642 640
rect 9642 584 9692 640
rect 9628 580 9692 584
rect 10364 580 10428 644
rect 11100 580 11164 644
rect 11836 580 11900 644
rect 12572 580 12636 644
rect 13308 580 13372 644
rect 16988 580 17052 644
rect 17724 580 17788 644
rect 18460 580 18524 644
rect 23612 580 23676 644
rect 28764 580 28828 644
rect 30236 580 30300 644
rect 35664 640 35728 644
rect 35664 584 35678 640
rect 35678 584 35728 640
rect 35664 580 35728 584
rect 36400 580 36464 644
rect 37136 580 37200 644
rect 37872 580 37936 644
rect 38608 640 38672 644
rect 38608 584 38622 640
rect 38622 584 38672 640
rect 38608 580 38672 584
rect 40080 580 40144 644
rect 40816 640 40880 644
rect 40816 584 40830 640
rect 40830 584 40880 640
rect 40816 580 40880 584
rect 41552 580 41616 644
rect 42288 580 42352 644
rect 43024 580 43088 644
rect 43760 580 43824 644
rect 44496 580 44560 644
rect 45232 580 45296 644
rect 45968 640 46032 644
rect 45968 584 45982 640
rect 45982 584 46032 640
rect 45968 580 46032 584
rect 46704 580 46768 644
rect 47440 580 47504 644
rect 48176 580 48240 644
rect 48912 580 48976 644
rect 49648 580 49712 644
rect 50384 580 50448 644
rect 51120 640 51184 644
rect 51120 584 51134 640
rect 51134 584 51184 640
rect 51120 580 51184 584
rect 51856 580 51920 644
rect 52592 580 52656 644
rect 53328 640 53392 644
rect 53328 584 53378 640
rect 53378 584 53392 640
rect 53328 580 53392 584
rect 54800 640 54864 644
rect 54800 584 54850 640
rect 54850 584 54864 640
rect 54800 580 54864 584
rect 55536 580 55600 644
rect 56272 640 56336 644
rect 56272 584 56286 640
rect 56286 584 56336 640
rect 56272 580 56336 584
rect 57008 640 57072 644
rect 57008 584 57058 640
rect 57058 584 57072 640
rect 57008 580 57072 584
rect 57744 640 57808 644
rect 57744 584 57794 640
rect 57794 584 57808 640
rect 57744 580 57808 584
rect 58480 580 58544 644
rect 60688 580 60752 644
rect 61424 580 61488 644
rect 62160 580 62224 644
rect 62896 640 62960 644
rect 62896 584 62946 640
rect 62946 584 62960 640
rect 62896 580 62960 584
rect 63632 580 63696 644
rect 64368 580 64432 644
rect 65104 580 65168 644
rect 72740 580 72804 644
rect 74948 580 75012 644
rect 138796 716 138860 720
rect 141004 716 141068 780
rect 143212 716 143276 780
rect 143948 716 144012 780
rect 145420 716 145484 780
rect 146156 776 146220 780
rect 146156 720 146206 776
rect 146206 720 146220 776
rect 146156 716 146220 720
rect 146892 716 146956 780
rect 148364 716 148428 780
rect 149100 716 149164 780
rect 150572 716 150636 780
rect 151308 716 151372 780
rect 152044 716 152108 780
rect 152780 716 152844 780
rect 154252 716 154316 780
rect 114232 640 114296 644
rect 114232 584 114246 640
rect 114246 584 114296 640
rect 114232 580 114296 584
rect 114968 580 115032 644
rect 115704 640 115768 644
rect 115704 584 115754 640
rect 115754 584 115768 640
rect 115704 580 115768 584
rect 116440 580 116504 644
rect 117912 580 117976 644
rect 118648 640 118712 644
rect 118648 584 118698 640
rect 118698 584 118712 640
rect 118648 580 118712 584
rect 119384 640 119448 644
rect 119384 584 119398 640
rect 119398 584 119448 640
rect 119384 580 119448 584
rect 120120 580 120184 644
rect 120856 580 120920 644
rect 121592 580 121656 644
rect 122328 580 122392 644
rect 123064 640 123128 644
rect 123064 584 123114 640
rect 123114 584 123128 640
rect 123064 580 123128 584
rect 123800 580 123864 644
rect 124536 580 124600 644
rect 125272 640 125336 644
rect 125272 584 125322 640
rect 125322 584 125336 640
rect 125272 580 125336 584
rect 126008 580 126072 644
rect 126744 640 126808 644
rect 126744 584 126794 640
rect 126794 584 126808 640
rect 126744 580 126808 584
rect 127480 580 127544 644
rect 128952 580 129016 644
rect 129688 580 129752 644
rect 131160 580 131224 644
rect 131896 580 131960 644
rect 132632 580 132696 644
rect 133368 580 133432 644
rect 134104 580 134168 644
rect 138060 580 138124 644
rect 141740 580 141804 644
rect 147628 580 147692 644
rect 153516 580 153580 644
rect 158668 580 158732 644
rect 160876 580 160940 644
rect 162348 580 162412 644
rect 164556 580 164620 644
rect 167500 580 167564 644
rect 168972 640 169036 644
rect 168972 584 169022 640
rect 169022 584 169036 640
rect 168972 580 169036 584
rect 250024 580 250088 644
rect 251496 640 251560 644
rect 251496 584 251546 640
rect 251546 584 251560 640
rect 251496 580 251560 584
rect 252232 640 252296 644
rect 252232 584 252282 640
rect 252282 584 252296 640
rect 252232 580 252296 584
rect 252968 580 253032 644
rect 253704 580 253768 644
rect 255176 640 255240 644
rect 255176 584 255226 640
rect 255226 584 255240 640
rect 255176 580 255240 584
rect 255912 580 255976 644
rect 256648 640 256712 644
rect 256648 584 256698 640
rect 256698 584 256712 640
rect 256648 580 256712 584
rect 257384 640 257448 644
rect 257384 584 257434 640
rect 257434 584 257448 640
rect 257384 580 257448 584
rect 258856 580 258920 644
rect 259592 580 259656 644
rect 260328 580 260392 644
rect 261064 580 261128 644
rect 262536 640 262600 644
rect 262536 584 262550 640
rect 262550 584 262600 640
rect 262536 580 262600 584
rect 263272 640 263336 644
rect 263272 584 263286 640
rect 263286 584 263336 640
rect 263272 580 263336 584
rect 264008 580 264072 644
rect 265480 580 265544 644
rect 266216 580 266280 644
rect 266952 640 267016 644
rect 266952 584 266966 640
rect 266966 584 267016 640
rect 266952 580 267016 584
rect 267688 640 267752 644
rect 267688 584 267702 640
rect 267702 584 267752 640
rect 267688 580 267752 584
rect 268424 640 268488 644
rect 268424 584 268438 640
rect 268438 584 268488 640
rect 268424 580 268488 584
rect 28028 444 28092 508
rect 29500 444 29564 508
rect 31708 444 31772 508
rect 65840 444 65904 508
rect 66576 444 66640 508
rect 30972 308 31036 372
rect 34928 308 34992 372
rect 39344 308 39408 372
rect 89668 308 89732 372
rect 91140 308 91204 372
rect 92612 308 92676 372
rect 97028 444 97092 508
rect 99972 504 100036 508
rect 99972 448 100022 504
rect 100022 448 100036 504
rect 99972 444 100036 448
rect 103192 504 103256 508
rect 103192 448 103242 504
rect 103242 448 103256 504
rect 103192 444 103256 448
rect 103928 504 103992 508
rect 103928 448 103942 504
rect 103942 448 103992 504
rect 103928 444 103992 448
rect 104664 504 104728 508
rect 104664 448 104714 504
rect 104714 448 104728 504
rect 104664 444 104728 448
rect 105400 444 105464 508
rect 106136 504 106200 508
rect 106136 448 106186 504
rect 106186 448 106200 504
rect 106136 444 106200 448
rect 106872 444 106936 508
rect 107608 444 107672 508
rect 108344 504 108408 508
rect 108344 448 108394 504
rect 108394 448 108408 504
rect 108344 444 108408 448
rect 109080 504 109144 508
rect 109080 448 109094 504
rect 109094 448 109144 504
rect 109080 444 109144 448
rect 109816 444 109880 508
rect 110552 444 110616 508
rect 111288 444 111352 508
rect 112024 444 112088 508
rect 112760 444 112824 508
rect 113496 368 113560 372
rect 113496 312 113546 368
rect 113546 312 113560 368
rect 113496 308 113560 312
rect 130424 308 130488 372
rect 139532 444 139596 508
rect 235028 444 235092 508
rect 241192 504 241256 508
rect 241192 448 241242 504
rect 241242 448 241256 504
rect 241192 444 241256 448
rect 241928 504 241992 508
rect 241928 448 241978 504
rect 241978 448 241992 504
rect 241928 444 241992 448
rect 243400 504 243464 508
rect 243400 448 243450 504
rect 243450 448 243464 504
rect 243400 444 243464 448
rect 244872 504 244936 508
rect 244872 448 244922 504
rect 244922 448 244936 504
rect 244872 444 244936 448
rect 245608 444 245672 508
rect 246344 504 246408 508
rect 246344 448 246394 504
rect 246394 448 246408 504
rect 246344 444 246408 448
rect 248552 444 248616 508
rect 261800 504 261864 508
rect 271339 1116 271403 1120
rect 271339 1060 271343 1116
rect 271343 1060 271399 1116
rect 271399 1060 271403 1116
rect 271339 1056 271403 1060
rect 271419 1116 271483 1120
rect 271419 1060 271423 1116
rect 271423 1060 271479 1116
rect 271479 1060 271483 1116
rect 271419 1056 271483 1060
rect 271499 1116 271563 1120
rect 271499 1060 271503 1116
rect 271503 1060 271559 1116
rect 271559 1060 271563 1116
rect 271499 1056 271563 1060
rect 271579 1116 271643 1120
rect 271579 1060 271583 1116
rect 271583 1060 271639 1116
rect 271639 1060 271643 1116
rect 271579 1056 271643 1060
rect 269896 580 269960 644
rect 261800 448 261850 504
rect 261850 448 261864 504
rect 261800 444 261864 448
rect 218836 368 218900 372
rect 218836 312 218886 368
rect 218886 312 218900 368
rect 218836 308 218900 312
rect 219572 368 219636 372
rect 219572 312 219622 368
rect 219622 312 219636 368
rect 219572 308 219636 312
rect 221780 308 221844 372
rect 229140 368 229204 372
rect 229140 312 229154 368
rect 229154 312 229204 368
rect 229140 308 229204 312
rect 229876 368 229940 372
rect 229876 312 229890 368
rect 229890 312 229940 368
rect 229876 308 229940 312
rect 230612 308 230676 372
rect 233556 308 233620 372
rect 234292 308 234356 372
rect 239720 308 239784 372
rect 240456 308 240520 372
rect 254440 308 254504 372
rect 269160 444 269224 508
rect 271368 308 271432 372
<< metal4 >>
rect 798 9213 858 10880
rect 1534 10165 1594 10880
rect 2270 10165 2330 10880
rect 1531 10164 1597 10165
rect 1531 10100 1532 10164
rect 1596 10100 1597 10164
rect 1531 10099 1597 10100
rect 2267 10164 2333 10165
rect 2267 10100 2268 10164
rect 2332 10100 2333 10164
rect 2267 10099 2333 10100
rect 3006 9893 3066 10880
rect 3742 10165 3802 10880
rect 4478 10165 4538 10880
rect 5214 10165 5274 10880
rect 5950 10165 6010 10880
rect 6686 10165 6746 10880
rect 7422 10165 7482 10880
rect 3739 10164 3805 10165
rect 3739 10100 3740 10164
rect 3804 10100 3805 10164
rect 3739 10099 3805 10100
rect 4475 10164 4541 10165
rect 4475 10100 4476 10164
rect 4540 10100 4541 10164
rect 4475 10099 4541 10100
rect 5211 10164 5277 10165
rect 5211 10100 5212 10164
rect 5276 10100 5277 10164
rect 5211 10099 5277 10100
rect 5947 10164 6013 10165
rect 5947 10100 5948 10164
rect 6012 10100 6013 10164
rect 5947 10099 6013 10100
rect 6683 10164 6749 10165
rect 6683 10100 6684 10164
rect 6748 10100 6749 10164
rect 6683 10099 6749 10100
rect 7419 10164 7485 10165
rect 7419 10100 7420 10164
rect 7484 10100 7485 10164
rect 7419 10099 7485 10100
rect 8158 9893 8218 10880
rect 8894 10165 8954 10880
rect 9630 10573 9690 10880
rect 9627 10572 9693 10573
rect 9627 10508 9628 10572
rect 9692 10508 9693 10572
rect 9627 10507 9693 10508
rect 8891 10164 8957 10165
rect 8891 10100 8892 10164
rect 8956 10100 8957 10164
rect 8891 10099 8957 10100
rect 10366 9893 10426 10880
rect 11102 9893 11162 10880
rect 11838 10165 11898 10880
rect 12574 10165 12634 10880
rect 11835 10164 11901 10165
rect 11835 10100 11836 10164
rect 11900 10100 11901 10164
rect 11835 10099 11901 10100
rect 12571 10164 12637 10165
rect 12571 10100 12572 10164
rect 12636 10100 12637 10164
rect 12571 10099 12637 10100
rect 13310 9893 13370 10880
rect 14046 10165 14106 10880
rect 14782 10165 14842 10880
rect 15518 10165 15578 10880
rect 16254 10165 16314 10880
rect 16990 10165 17050 10880
rect 17726 10165 17786 10880
rect 18462 10165 18522 10880
rect 14043 10164 14109 10165
rect 14043 10100 14044 10164
rect 14108 10100 14109 10164
rect 14043 10099 14109 10100
rect 14779 10164 14845 10165
rect 14779 10100 14780 10164
rect 14844 10100 14845 10164
rect 14779 10099 14845 10100
rect 15515 10164 15581 10165
rect 15515 10100 15516 10164
rect 15580 10100 15581 10164
rect 15515 10099 15581 10100
rect 16251 10164 16317 10165
rect 16251 10100 16252 10164
rect 16316 10100 16317 10164
rect 16251 10099 16317 10100
rect 16987 10164 17053 10165
rect 16987 10100 16988 10164
rect 17052 10100 17053 10164
rect 16987 10099 17053 10100
rect 17723 10164 17789 10165
rect 17723 10100 17724 10164
rect 17788 10100 17789 10164
rect 17723 10099 17789 10100
rect 18459 10164 18525 10165
rect 18459 10100 18460 10164
rect 18524 10100 18525 10164
rect 18459 10099 18525 10100
rect 3003 9892 3069 9893
rect 3003 9828 3004 9892
rect 3068 9828 3069 9892
rect 3003 9827 3069 9828
rect 8155 9892 8221 9893
rect 8155 9828 8156 9892
rect 8220 9828 8221 9892
rect 8155 9827 8221 9828
rect 10363 9892 10429 9893
rect 10363 9828 10364 9892
rect 10428 9828 10429 9892
rect 10363 9827 10429 9828
rect 11099 9892 11165 9893
rect 11099 9828 11100 9892
rect 11164 9828 11165 9892
rect 11099 9827 11165 9828
rect 13307 9892 13373 9893
rect 13307 9828 13308 9892
rect 13372 9828 13373 9892
rect 13307 9827 13373 9828
rect 795 9212 861 9213
rect 795 9148 796 9212
rect 860 9148 861 9212
rect 795 9147 861 9148
rect 19198 6901 19258 10880
rect 19934 6901 19994 10880
rect 20670 10573 20730 10880
rect 20667 10572 20733 10573
rect 20667 10508 20668 10572
rect 20732 10508 20733 10572
rect 20667 10507 20733 10508
rect 21406 9893 21466 10880
rect 22142 10165 22202 10880
rect 22139 10164 22205 10165
rect 22139 10100 22140 10164
rect 22204 10100 22205 10164
rect 22139 10099 22205 10100
rect 21403 9892 21469 9893
rect 21403 9828 21404 9892
rect 21468 9828 21469 9892
rect 21403 9827 21469 9828
rect 22878 6901 22938 10880
rect 23614 6901 23674 10880
rect 24350 8669 24410 10880
rect 24347 8668 24413 8669
rect 24347 8604 24348 8668
rect 24412 8604 24413 8668
rect 24347 8603 24413 8604
rect 25086 6901 25146 10880
rect 25822 9621 25882 10880
rect 25819 9620 25885 9621
rect 25819 9556 25820 9620
rect 25884 9556 25885 9620
rect 25819 9555 25885 9556
rect 26558 8397 26618 10880
rect 26555 8396 26621 8397
rect 26555 8332 26556 8396
rect 26620 8332 26621 8396
rect 26555 8331 26621 8332
rect 27294 7853 27354 10880
rect 28030 8397 28090 10880
rect 28766 9485 28826 10880
rect 28763 9484 28829 9485
rect 28763 9420 28764 9484
rect 28828 9420 28829 9484
rect 28763 9419 28829 9420
rect 29502 8669 29562 10880
rect 30238 8669 30298 10880
rect 30974 8669 31034 10880
rect 31710 10301 31770 10880
rect 31707 10300 31773 10301
rect 31707 10236 31708 10300
rect 31772 10236 31773 10300
rect 31707 10235 31773 10236
rect 32446 9621 32506 10880
rect 34930 10301 34990 10880
rect 35666 10301 35726 10880
rect 36402 10301 36462 10880
rect 37138 10301 37198 10880
rect 37874 10301 37934 10880
rect 38610 10301 38670 10880
rect 39346 10301 39406 10880
rect 40082 10301 40142 10880
rect 40818 10301 40878 10880
rect 41554 10301 41614 10880
rect 42290 10301 42350 10880
rect 43026 10301 43086 10880
rect 43762 10301 43822 10880
rect 44498 10301 44558 10880
rect 45234 10301 45294 10880
rect 45970 10301 46030 10880
rect 46706 10301 46766 10880
rect 47442 10301 47502 10880
rect 48178 10301 48238 10880
rect 48914 10301 48974 10880
rect 49650 10301 49710 10880
rect 50386 10301 50446 10880
rect 51122 10301 51182 10880
rect 51858 10301 51918 10880
rect 52594 10301 52654 10880
rect 53330 10301 53390 10880
rect 54066 10437 54126 10880
rect 54063 10436 54129 10437
rect 54063 10372 54064 10436
rect 54128 10372 54129 10436
rect 54063 10371 54129 10372
rect 54802 10301 54862 10880
rect 55538 10301 55598 10880
rect 56274 10301 56334 10880
rect 57010 10301 57070 10880
rect 57746 10301 57806 10880
rect 58482 10301 58542 10880
rect 59218 10301 59278 10880
rect 59954 10301 60014 10880
rect 60690 10301 60750 10880
rect 61426 10301 61486 10880
rect 62162 10301 62222 10880
rect 62898 10301 62958 10880
rect 63634 10301 63694 10880
rect 64370 10301 64430 10880
rect 65106 10301 65166 10880
rect 65842 10301 65902 10880
rect 66578 10301 66638 10880
rect 34927 10300 34993 10301
rect 34927 10236 34928 10300
rect 34992 10236 34993 10300
rect 34927 10235 34993 10236
rect 35663 10300 35729 10301
rect 35663 10236 35664 10300
rect 35728 10236 35729 10300
rect 35663 10235 35729 10236
rect 36399 10300 36465 10301
rect 36399 10236 36400 10300
rect 36464 10236 36465 10300
rect 36399 10235 36465 10236
rect 37135 10300 37201 10301
rect 37135 10236 37136 10300
rect 37200 10236 37201 10300
rect 37135 10235 37201 10236
rect 37871 10300 37937 10301
rect 37871 10236 37872 10300
rect 37936 10236 37937 10300
rect 37871 10235 37937 10236
rect 38607 10300 38673 10301
rect 38607 10236 38608 10300
rect 38672 10236 38673 10300
rect 38607 10235 38673 10236
rect 39343 10300 39409 10301
rect 39343 10236 39344 10300
rect 39408 10236 39409 10300
rect 39343 10235 39409 10236
rect 40079 10300 40145 10301
rect 40079 10236 40080 10300
rect 40144 10236 40145 10300
rect 40079 10235 40145 10236
rect 40815 10300 40881 10301
rect 40815 10236 40816 10300
rect 40880 10236 40881 10300
rect 40815 10235 40881 10236
rect 41551 10300 41617 10301
rect 41551 10236 41552 10300
rect 41616 10236 41617 10300
rect 41551 10235 41617 10236
rect 42287 10300 42353 10301
rect 42287 10236 42288 10300
rect 42352 10236 42353 10300
rect 42287 10235 42353 10236
rect 43023 10300 43089 10301
rect 43023 10236 43024 10300
rect 43088 10236 43089 10300
rect 43023 10235 43089 10236
rect 43759 10300 43825 10301
rect 43759 10236 43760 10300
rect 43824 10236 43825 10300
rect 43759 10235 43825 10236
rect 44495 10300 44561 10301
rect 44495 10236 44496 10300
rect 44560 10236 44561 10300
rect 44495 10235 44561 10236
rect 45231 10300 45297 10301
rect 45231 10236 45232 10300
rect 45296 10236 45297 10300
rect 45231 10235 45297 10236
rect 45967 10300 46033 10301
rect 45967 10236 45968 10300
rect 46032 10236 46033 10300
rect 45967 10235 46033 10236
rect 46703 10300 46769 10301
rect 46703 10236 46704 10300
rect 46768 10236 46769 10300
rect 46703 10235 46769 10236
rect 47439 10300 47505 10301
rect 47439 10236 47440 10300
rect 47504 10236 47505 10300
rect 47439 10235 47505 10236
rect 48175 10300 48241 10301
rect 48175 10236 48176 10300
rect 48240 10236 48241 10300
rect 48175 10235 48241 10236
rect 48911 10300 48977 10301
rect 48911 10236 48912 10300
rect 48976 10236 48977 10300
rect 48911 10235 48977 10236
rect 49647 10300 49713 10301
rect 49647 10236 49648 10300
rect 49712 10236 49713 10300
rect 49647 10235 49713 10236
rect 50383 10300 50449 10301
rect 50383 10236 50384 10300
rect 50448 10236 50449 10300
rect 50383 10235 50449 10236
rect 51119 10300 51185 10301
rect 51119 10236 51120 10300
rect 51184 10236 51185 10300
rect 51119 10235 51185 10236
rect 51855 10300 51921 10301
rect 51855 10236 51856 10300
rect 51920 10236 51921 10300
rect 51855 10235 51921 10236
rect 52591 10300 52657 10301
rect 52591 10236 52592 10300
rect 52656 10236 52657 10300
rect 52591 10235 52657 10236
rect 53327 10300 53393 10301
rect 53327 10236 53328 10300
rect 53392 10236 53393 10300
rect 53327 10235 53393 10236
rect 54799 10300 54865 10301
rect 54799 10236 54800 10300
rect 54864 10236 54865 10300
rect 54799 10235 54865 10236
rect 55535 10300 55601 10301
rect 55535 10236 55536 10300
rect 55600 10236 55601 10300
rect 55535 10235 55601 10236
rect 56271 10300 56337 10301
rect 56271 10236 56272 10300
rect 56336 10236 56337 10300
rect 56271 10235 56337 10236
rect 57007 10300 57073 10301
rect 57007 10236 57008 10300
rect 57072 10236 57073 10300
rect 57007 10235 57073 10236
rect 57743 10300 57809 10301
rect 57743 10236 57744 10300
rect 57808 10236 57809 10300
rect 57743 10235 57809 10236
rect 58479 10300 58545 10301
rect 58479 10236 58480 10300
rect 58544 10236 58545 10300
rect 58479 10235 58545 10236
rect 59215 10300 59281 10301
rect 59215 10236 59216 10300
rect 59280 10236 59281 10300
rect 59215 10235 59281 10236
rect 59951 10300 60017 10301
rect 59951 10236 59952 10300
rect 60016 10236 60017 10300
rect 59951 10235 60017 10236
rect 60687 10300 60753 10301
rect 60687 10236 60688 10300
rect 60752 10236 60753 10300
rect 60687 10235 60753 10236
rect 61423 10300 61489 10301
rect 61423 10236 61424 10300
rect 61488 10236 61489 10300
rect 61423 10235 61489 10236
rect 62159 10300 62225 10301
rect 62159 10236 62160 10300
rect 62224 10236 62225 10300
rect 62159 10235 62225 10236
rect 62895 10300 62961 10301
rect 62895 10236 62896 10300
rect 62960 10236 62961 10300
rect 62895 10235 62961 10236
rect 63631 10300 63697 10301
rect 63631 10236 63632 10300
rect 63696 10236 63697 10300
rect 63631 10235 63697 10236
rect 64367 10300 64433 10301
rect 64367 10236 64368 10300
rect 64432 10236 64433 10300
rect 64367 10235 64433 10236
rect 65103 10300 65169 10301
rect 65103 10236 65104 10300
rect 65168 10236 65169 10300
rect 65103 10235 65169 10236
rect 65839 10300 65905 10301
rect 65839 10236 65840 10300
rect 65904 10236 65905 10300
rect 65839 10235 65905 10236
rect 66575 10300 66641 10301
rect 66575 10236 66576 10300
rect 66640 10236 66641 10300
rect 66575 10235 66641 10236
rect 32443 9620 32509 9621
rect 32443 9556 32444 9620
rect 32508 9556 32509 9620
rect 32443 9555 32509 9556
rect 34742 9280 35062 9840
rect 34742 9216 34750 9280
rect 34814 9216 34830 9280
rect 34894 9216 34910 9280
rect 34974 9216 34990 9280
rect 35054 9216 35062 9280
rect 29499 8668 29565 8669
rect 29499 8604 29500 8668
rect 29564 8604 29565 8668
rect 29499 8603 29565 8604
rect 30235 8668 30301 8669
rect 30235 8604 30236 8668
rect 30300 8604 30301 8668
rect 30235 8603 30301 8604
rect 30971 8668 31037 8669
rect 30971 8604 30972 8668
rect 31036 8604 31037 8668
rect 30971 8603 31037 8604
rect 28027 8396 28093 8397
rect 28027 8332 28028 8396
rect 28092 8332 28093 8396
rect 28027 8331 28093 8332
rect 34742 8192 35062 9216
rect 34742 8128 34750 8192
rect 34814 8128 34830 8192
rect 34894 8128 34910 8192
rect 34974 8128 34990 8192
rect 35054 8128 35062 8192
rect 27291 7852 27357 7853
rect 27291 7788 27292 7852
rect 27356 7788 27357 7852
rect 27291 7787 27357 7788
rect 34742 7104 35062 8128
rect 34742 7040 34750 7104
rect 34814 7040 34830 7104
rect 34894 7040 34910 7104
rect 34974 7040 34990 7104
rect 35054 7040 35062 7104
rect 19195 6900 19261 6901
rect 19195 6836 19196 6900
rect 19260 6836 19261 6900
rect 19195 6835 19261 6836
rect 19931 6900 19997 6901
rect 19931 6836 19932 6900
rect 19996 6836 19997 6900
rect 19931 6835 19997 6836
rect 22875 6900 22941 6901
rect 22875 6836 22876 6900
rect 22940 6836 22941 6900
rect 22875 6835 22941 6836
rect 23611 6900 23677 6901
rect 23611 6836 23612 6900
rect 23676 6836 23677 6900
rect 23611 6835 23677 6836
rect 25083 6900 25149 6901
rect 25083 6836 25084 6900
rect 25148 6836 25149 6900
rect 25083 6835 25149 6836
rect 34742 6016 35062 7040
rect 34742 5952 34750 6016
rect 34814 5952 34830 6016
rect 34894 5952 34910 6016
rect 34974 5952 34990 6016
rect 35054 5952 35062 6016
rect 34742 4928 35062 5952
rect 34742 4864 34750 4928
rect 34814 4864 34830 4928
rect 34894 4864 34910 4928
rect 34974 4864 34990 4928
rect 35054 4864 35062 4928
rect 34742 3840 35062 4864
rect 34742 3776 34750 3840
rect 34814 3776 34830 3840
rect 34894 3776 34910 3840
rect 34974 3776 34990 3840
rect 35054 3776 35062 3840
rect 24347 3364 24413 3365
rect 24347 3300 24348 3364
rect 24412 3300 24413 3364
rect 24347 3299 24413 3300
rect 19195 2956 19261 2957
rect 19195 2892 19196 2956
rect 19260 2892 19261 2956
rect 19195 2891 19261 2892
rect 22875 2956 22941 2957
rect 22875 2892 22876 2956
rect 22940 2892 22941 2956
rect 22875 2891 22941 2892
rect 795 1460 861 1461
rect 795 1396 796 1460
rect 860 1396 861 1460
rect 795 1395 861 1396
rect 16251 1460 16317 1461
rect 16251 1396 16252 1460
rect 16316 1396 16317 1460
rect 16251 1395 16317 1396
rect 798 0 858 1395
rect 1531 1324 1597 1325
rect 1531 1260 1532 1324
rect 1596 1260 1597 1324
rect 1531 1259 1597 1260
rect 1534 0 1594 1259
rect 2267 1052 2333 1053
rect 2267 988 2268 1052
rect 2332 988 2333 1052
rect 2267 987 2333 988
rect 4475 1052 4541 1053
rect 4475 988 4476 1052
rect 4540 988 4541 1052
rect 4475 987 4541 988
rect 6683 1052 6749 1053
rect 6683 988 6684 1052
rect 6748 988 6749 1052
rect 6683 987 6749 988
rect 14043 1052 14109 1053
rect 14043 988 14044 1052
rect 14108 988 14109 1052
rect 14043 987 14109 988
rect 2270 0 2330 987
rect 3003 780 3069 781
rect 3003 716 3004 780
rect 3068 716 3069 780
rect 3003 715 3069 716
rect 3006 0 3066 715
rect 3739 644 3805 645
rect 3739 580 3740 644
rect 3804 580 3805 644
rect 3739 579 3805 580
rect 3742 0 3802 579
rect 4478 0 4538 987
rect 5211 780 5277 781
rect 5211 716 5212 780
rect 5276 716 5277 780
rect 5211 715 5277 716
rect 5947 780 6013 781
rect 5947 716 5948 780
rect 6012 716 6013 780
rect 5947 715 6013 716
rect 5214 0 5274 715
rect 5950 0 6010 715
rect 6686 0 6746 987
rect 7419 780 7485 781
rect 7419 716 7420 780
rect 7484 716 7485 780
rect 7419 715 7485 716
rect 8891 780 8957 781
rect 8891 716 8892 780
rect 8956 716 8957 780
rect 8891 715 8957 716
rect 7422 0 7482 715
rect 8155 644 8221 645
rect 8155 580 8156 644
rect 8220 580 8221 644
rect 8155 579 8221 580
rect 8158 0 8218 579
rect 8894 0 8954 715
rect 9627 644 9693 645
rect 9627 580 9628 644
rect 9692 580 9693 644
rect 9627 579 9693 580
rect 10363 644 10429 645
rect 10363 580 10364 644
rect 10428 580 10429 644
rect 10363 579 10429 580
rect 11099 644 11165 645
rect 11099 580 11100 644
rect 11164 580 11165 644
rect 11099 579 11165 580
rect 11835 644 11901 645
rect 11835 580 11836 644
rect 11900 580 11901 644
rect 11835 579 11901 580
rect 12571 644 12637 645
rect 12571 580 12572 644
rect 12636 580 12637 644
rect 12571 579 12637 580
rect 13307 644 13373 645
rect 13307 580 13308 644
rect 13372 580 13373 644
rect 13307 579 13373 580
rect 9630 0 9690 579
rect 10366 0 10426 579
rect 11102 0 11162 579
rect 11838 0 11898 579
rect 12574 0 12634 579
rect 13310 0 13370 579
rect 14046 0 14106 987
rect 14779 780 14845 781
rect 14779 716 14780 780
rect 14844 716 14845 780
rect 14779 715 14845 716
rect 15515 780 15581 781
rect 15515 716 15516 780
rect 15580 716 15581 780
rect 15515 715 15581 716
rect 14782 0 14842 715
rect 15518 0 15578 715
rect 16254 0 16314 1395
rect 16987 644 17053 645
rect 16987 580 16988 644
rect 17052 580 17053 644
rect 16987 579 17053 580
rect 17723 644 17789 645
rect 17723 580 17724 644
rect 17788 580 17789 644
rect 17723 579 17789 580
rect 18459 644 18525 645
rect 18459 580 18460 644
rect 18524 580 18525 644
rect 18459 579 18525 580
rect 16990 0 17050 579
rect 17726 0 17786 579
rect 18462 0 18522 579
rect 19198 0 19258 2891
rect 19931 2820 19997 2821
rect 19931 2756 19932 2820
rect 19996 2756 19997 2820
rect 19931 2755 19997 2756
rect 22139 2820 22205 2821
rect 22139 2756 22140 2820
rect 22204 2756 22205 2820
rect 22139 2755 22205 2756
rect 19934 0 19994 2755
rect 21403 1732 21469 1733
rect 21403 1668 21404 1732
rect 21468 1668 21469 1732
rect 21403 1667 21469 1668
rect 20667 1460 20733 1461
rect 20667 1396 20668 1460
rect 20732 1396 20733 1460
rect 20667 1395 20733 1396
rect 20670 0 20730 1395
rect 21406 0 21466 1667
rect 22142 0 22202 2755
rect 22878 0 22938 2891
rect 23611 644 23677 645
rect 23611 580 23612 644
rect 23676 580 23677 644
rect 23611 579 23677 580
rect 23614 0 23674 579
rect 24350 0 24410 3299
rect 25083 2820 25149 2821
rect 25083 2756 25084 2820
rect 25148 2756 25149 2820
rect 25083 2755 25149 2756
rect 25086 0 25146 2755
rect 34742 2752 35062 3776
rect 68540 9824 68860 9840
rect 68540 9760 68548 9824
rect 68612 9760 68628 9824
rect 68692 9760 68708 9824
rect 68772 9760 68788 9824
rect 68852 9760 68860 9824
rect 68540 8736 68860 9760
rect 69062 9621 69122 10880
rect 69059 9620 69125 9621
rect 69059 9556 69060 9620
rect 69124 9556 69125 9620
rect 69059 9555 69125 9556
rect 69798 9077 69858 10880
rect 70534 9621 70594 10880
rect 71270 10573 71330 10880
rect 71267 10572 71333 10573
rect 71267 10508 71268 10572
rect 71332 10508 71333 10572
rect 71267 10507 71333 10508
rect 72006 10437 72066 10880
rect 72003 10436 72069 10437
rect 72003 10372 72004 10436
rect 72068 10372 72069 10436
rect 72003 10371 72069 10372
rect 72742 9621 72802 10880
rect 70531 9620 70597 9621
rect 70531 9556 70532 9620
rect 70596 9556 70597 9620
rect 70531 9555 70597 9556
rect 72739 9620 72805 9621
rect 72739 9556 72740 9620
rect 72804 9556 72805 9620
rect 72739 9555 72805 9556
rect 73478 9077 73538 10880
rect 74214 10573 74274 10880
rect 74211 10572 74277 10573
rect 74211 10508 74212 10572
rect 74276 10508 74277 10572
rect 74211 10507 74277 10508
rect 74950 9077 75010 10880
rect 75686 9621 75746 10880
rect 76422 9757 76482 10880
rect 77158 10437 77218 10880
rect 77155 10436 77221 10437
rect 77155 10372 77156 10436
rect 77220 10372 77221 10436
rect 77155 10371 77221 10372
rect 76419 9756 76485 9757
rect 76419 9692 76420 9756
rect 76484 9692 76485 9756
rect 76419 9691 76485 9692
rect 77894 9621 77954 10880
rect 75683 9620 75749 9621
rect 75683 9556 75684 9620
rect 75748 9556 75749 9620
rect 75683 9555 75749 9556
rect 77891 9620 77957 9621
rect 77891 9556 77892 9620
rect 77956 9556 77957 9620
rect 77891 9555 77957 9556
rect 78630 9077 78690 10880
rect 79366 9757 79426 10880
rect 79363 9756 79429 9757
rect 79363 9692 79364 9756
rect 79428 9692 79429 9756
rect 79363 9691 79429 9692
rect 80102 9077 80162 10880
rect 80838 9621 80898 10880
rect 81574 9757 81634 10880
rect 82310 10437 82370 10880
rect 82307 10436 82373 10437
rect 82307 10372 82308 10436
rect 82372 10372 82373 10436
rect 82307 10371 82373 10372
rect 81571 9756 81637 9757
rect 81571 9692 81572 9756
rect 81636 9692 81637 9756
rect 81571 9691 81637 9692
rect 83046 9621 83106 10880
rect 83782 10437 83842 10880
rect 84518 10573 84578 10880
rect 84515 10572 84581 10573
rect 84515 10508 84516 10572
rect 84580 10508 84581 10572
rect 84515 10507 84581 10508
rect 83779 10436 83845 10437
rect 83779 10372 83780 10436
rect 83844 10372 83845 10436
rect 83779 10371 83845 10372
rect 85254 9893 85314 10880
rect 85990 9893 86050 10880
rect 86726 10573 86786 10880
rect 86723 10572 86789 10573
rect 86723 10508 86724 10572
rect 86788 10508 86789 10572
rect 86723 10507 86789 10508
rect 85251 9892 85317 9893
rect 85251 9828 85252 9892
rect 85316 9828 85317 9892
rect 85251 9827 85317 9828
rect 85987 9892 86053 9893
rect 85987 9828 85988 9892
rect 86052 9828 86053 9892
rect 85987 9827 86053 9828
rect 80835 9620 80901 9621
rect 80835 9556 80836 9620
rect 80900 9556 80901 9620
rect 80835 9555 80901 9556
rect 83043 9620 83109 9621
rect 83043 9556 83044 9620
rect 83108 9556 83109 9620
rect 83043 9555 83109 9556
rect 69795 9076 69861 9077
rect 69795 9012 69796 9076
rect 69860 9012 69861 9076
rect 69795 9011 69861 9012
rect 73475 9076 73541 9077
rect 73475 9012 73476 9076
rect 73540 9012 73541 9076
rect 73475 9011 73541 9012
rect 74947 9076 75013 9077
rect 74947 9012 74948 9076
rect 75012 9012 75013 9076
rect 74947 9011 75013 9012
rect 78627 9076 78693 9077
rect 78627 9012 78628 9076
rect 78692 9012 78693 9076
rect 78627 9011 78693 9012
rect 80099 9076 80165 9077
rect 80099 9012 80100 9076
rect 80164 9012 80165 9076
rect 80099 9011 80165 9012
rect 68540 8672 68548 8736
rect 68612 8672 68628 8736
rect 68692 8672 68708 8736
rect 68772 8672 68788 8736
rect 68852 8672 68860 8736
rect 68540 7648 68860 8672
rect 87462 8669 87522 10880
rect 88198 9213 88258 10880
rect 88195 9212 88261 9213
rect 88195 9148 88196 9212
rect 88260 9148 88261 9212
rect 88195 9147 88261 9148
rect 87459 8668 87525 8669
rect 87459 8604 87460 8668
rect 87524 8604 87525 8668
rect 87459 8603 87525 8604
rect 88934 8125 88994 10880
rect 89670 10301 89730 10880
rect 89667 10300 89733 10301
rect 89667 10236 89668 10300
rect 89732 10236 89733 10300
rect 89667 10235 89733 10236
rect 90406 8669 90466 10880
rect 91142 8805 91202 10880
rect 91139 8804 91205 8805
rect 91139 8740 91140 8804
rect 91204 8740 91205 8804
rect 91139 8739 91205 8740
rect 91878 8669 91938 10880
rect 90403 8668 90469 8669
rect 90403 8604 90404 8668
rect 90468 8604 90469 8668
rect 90403 8603 90469 8604
rect 91875 8668 91941 8669
rect 91875 8604 91876 8668
rect 91940 8604 91941 8668
rect 91875 8603 91941 8604
rect 92614 8397 92674 10880
rect 93350 9757 93410 10880
rect 93347 9756 93413 9757
rect 93347 9692 93348 9756
rect 93412 9692 93413 9756
rect 93347 9691 93413 9692
rect 94086 8669 94146 10880
rect 94822 8669 94882 10880
rect 95558 9757 95618 10880
rect 96294 9757 96354 10880
rect 95555 9756 95621 9757
rect 95555 9692 95556 9756
rect 95620 9692 95621 9756
rect 95555 9691 95621 9692
rect 96291 9756 96357 9757
rect 96291 9692 96292 9756
rect 96356 9692 96357 9756
rect 96291 9691 96357 9692
rect 97030 8669 97090 10880
rect 97766 9757 97826 10880
rect 97763 9756 97829 9757
rect 97763 9692 97764 9756
rect 97828 9692 97829 9756
rect 97763 9691 97829 9692
rect 98502 8669 98562 10880
rect 94083 8668 94149 8669
rect 94083 8604 94084 8668
rect 94148 8604 94149 8668
rect 94083 8603 94149 8604
rect 94819 8668 94885 8669
rect 94819 8604 94820 8668
rect 94884 8604 94885 8668
rect 94819 8603 94885 8604
rect 97027 8668 97093 8669
rect 97027 8604 97028 8668
rect 97092 8604 97093 8668
rect 97027 8603 97093 8604
rect 98499 8668 98565 8669
rect 98499 8604 98500 8668
rect 98564 8604 98565 8668
rect 98499 8603 98565 8604
rect 92611 8396 92677 8397
rect 92611 8332 92612 8396
rect 92676 8332 92677 8396
rect 92611 8331 92677 8332
rect 99238 8261 99298 10880
rect 99974 8669 100034 10880
rect 100710 9757 100770 10880
rect 103194 10301 103254 10880
rect 103930 10301 103990 10880
rect 104666 10301 104726 10880
rect 105402 10301 105462 10880
rect 106138 10301 106198 10880
rect 106874 10301 106934 10880
rect 107610 10301 107670 10880
rect 108346 10301 108406 10880
rect 109082 10301 109142 10880
rect 109818 10301 109878 10880
rect 110554 10301 110614 10880
rect 111290 10301 111350 10880
rect 112026 10301 112086 10880
rect 112762 10301 112822 10880
rect 113498 10301 113558 10880
rect 114234 10301 114294 10880
rect 114970 10301 115030 10880
rect 115706 10301 115766 10880
rect 116442 10301 116502 10880
rect 117178 10301 117238 10880
rect 117914 10301 117974 10880
rect 118650 10301 118710 10880
rect 119386 10301 119446 10880
rect 120122 10301 120182 10880
rect 120858 10301 120918 10880
rect 121594 10301 121654 10880
rect 122330 10301 122390 10880
rect 123066 10301 123126 10880
rect 123802 10301 123862 10880
rect 124538 10301 124598 10880
rect 125274 10437 125334 10880
rect 125271 10436 125337 10437
rect 125271 10372 125272 10436
rect 125336 10372 125337 10436
rect 125271 10371 125337 10372
rect 126010 10301 126070 10880
rect 126746 10301 126806 10880
rect 127482 10301 127542 10880
rect 128218 10437 128278 10880
rect 128215 10436 128281 10437
rect 128215 10372 128216 10436
rect 128280 10372 128281 10436
rect 128215 10371 128281 10372
rect 128954 10301 129014 10880
rect 129690 10301 129750 10880
rect 130426 10301 130486 10880
rect 131162 10301 131222 10880
rect 131898 10301 131958 10880
rect 132634 10301 132694 10880
rect 133370 10301 133430 10880
rect 134106 10301 134166 10880
rect 134842 10301 134902 10880
rect 103191 10300 103257 10301
rect 103191 10236 103192 10300
rect 103256 10236 103257 10300
rect 103191 10235 103257 10236
rect 103927 10300 103993 10301
rect 103927 10236 103928 10300
rect 103992 10236 103993 10300
rect 103927 10235 103993 10236
rect 104663 10300 104729 10301
rect 104663 10236 104664 10300
rect 104728 10236 104729 10300
rect 104663 10235 104729 10236
rect 105399 10300 105465 10301
rect 105399 10236 105400 10300
rect 105464 10236 105465 10300
rect 105399 10235 105465 10236
rect 106135 10300 106201 10301
rect 106135 10236 106136 10300
rect 106200 10236 106201 10300
rect 106135 10235 106201 10236
rect 106871 10300 106937 10301
rect 106871 10236 106872 10300
rect 106936 10236 106937 10300
rect 106871 10235 106937 10236
rect 107607 10300 107673 10301
rect 107607 10236 107608 10300
rect 107672 10236 107673 10300
rect 107607 10235 107673 10236
rect 108343 10300 108409 10301
rect 108343 10236 108344 10300
rect 108408 10236 108409 10300
rect 108343 10235 108409 10236
rect 109079 10300 109145 10301
rect 109079 10236 109080 10300
rect 109144 10236 109145 10300
rect 109079 10235 109145 10236
rect 109815 10300 109881 10301
rect 109815 10236 109816 10300
rect 109880 10236 109881 10300
rect 109815 10235 109881 10236
rect 110551 10300 110617 10301
rect 110551 10236 110552 10300
rect 110616 10236 110617 10300
rect 110551 10235 110617 10236
rect 111287 10300 111353 10301
rect 111287 10236 111288 10300
rect 111352 10236 111353 10300
rect 111287 10235 111353 10236
rect 112023 10300 112089 10301
rect 112023 10236 112024 10300
rect 112088 10236 112089 10300
rect 112023 10235 112089 10236
rect 112759 10300 112825 10301
rect 112759 10236 112760 10300
rect 112824 10236 112825 10300
rect 112759 10235 112825 10236
rect 113495 10300 113561 10301
rect 113495 10236 113496 10300
rect 113560 10236 113561 10300
rect 113495 10235 113561 10236
rect 114231 10300 114297 10301
rect 114231 10236 114232 10300
rect 114296 10236 114297 10300
rect 114231 10235 114297 10236
rect 114967 10300 115033 10301
rect 114967 10236 114968 10300
rect 115032 10236 115033 10300
rect 114967 10235 115033 10236
rect 115703 10300 115769 10301
rect 115703 10236 115704 10300
rect 115768 10236 115769 10300
rect 115703 10235 115769 10236
rect 116439 10300 116505 10301
rect 116439 10236 116440 10300
rect 116504 10236 116505 10300
rect 116439 10235 116505 10236
rect 117175 10300 117241 10301
rect 117175 10236 117176 10300
rect 117240 10236 117241 10300
rect 117175 10235 117241 10236
rect 117911 10300 117977 10301
rect 117911 10236 117912 10300
rect 117976 10236 117977 10300
rect 117911 10235 117977 10236
rect 118647 10300 118713 10301
rect 118647 10236 118648 10300
rect 118712 10236 118713 10300
rect 118647 10235 118713 10236
rect 119383 10300 119449 10301
rect 119383 10236 119384 10300
rect 119448 10236 119449 10300
rect 119383 10235 119449 10236
rect 120119 10300 120185 10301
rect 120119 10236 120120 10300
rect 120184 10236 120185 10300
rect 120119 10235 120185 10236
rect 120855 10300 120921 10301
rect 120855 10236 120856 10300
rect 120920 10236 120921 10300
rect 120855 10235 120921 10236
rect 121591 10300 121657 10301
rect 121591 10236 121592 10300
rect 121656 10236 121657 10300
rect 121591 10235 121657 10236
rect 122327 10300 122393 10301
rect 122327 10236 122328 10300
rect 122392 10236 122393 10300
rect 122327 10235 122393 10236
rect 123063 10300 123129 10301
rect 123063 10236 123064 10300
rect 123128 10236 123129 10300
rect 123063 10235 123129 10236
rect 123799 10300 123865 10301
rect 123799 10236 123800 10300
rect 123864 10236 123865 10300
rect 123799 10235 123865 10236
rect 124535 10300 124601 10301
rect 124535 10236 124536 10300
rect 124600 10236 124601 10300
rect 124535 10235 124601 10236
rect 126007 10300 126073 10301
rect 126007 10236 126008 10300
rect 126072 10236 126073 10300
rect 126007 10235 126073 10236
rect 126743 10300 126809 10301
rect 126743 10236 126744 10300
rect 126808 10236 126809 10300
rect 126743 10235 126809 10236
rect 127479 10300 127545 10301
rect 127479 10236 127480 10300
rect 127544 10236 127545 10300
rect 127479 10235 127545 10236
rect 128951 10300 129017 10301
rect 128951 10236 128952 10300
rect 129016 10236 129017 10300
rect 128951 10235 129017 10236
rect 129687 10300 129753 10301
rect 129687 10236 129688 10300
rect 129752 10236 129753 10300
rect 129687 10235 129753 10236
rect 130423 10300 130489 10301
rect 130423 10236 130424 10300
rect 130488 10236 130489 10300
rect 130423 10235 130489 10236
rect 131159 10300 131225 10301
rect 131159 10236 131160 10300
rect 131224 10236 131225 10300
rect 131159 10235 131225 10236
rect 131895 10300 131961 10301
rect 131895 10236 131896 10300
rect 131960 10236 131961 10300
rect 131895 10235 131961 10236
rect 132631 10300 132697 10301
rect 132631 10236 132632 10300
rect 132696 10236 132697 10300
rect 132631 10235 132697 10236
rect 133367 10300 133433 10301
rect 133367 10236 133368 10300
rect 133432 10236 133433 10300
rect 133367 10235 133433 10236
rect 134103 10300 134169 10301
rect 134103 10236 134104 10300
rect 134168 10236 134169 10300
rect 134103 10235 134169 10236
rect 134839 10300 134905 10301
rect 134839 10236 134840 10300
rect 134904 10236 134905 10300
rect 134839 10235 134905 10236
rect 100707 9756 100773 9757
rect 100707 9692 100708 9756
rect 100772 9692 100773 9756
rect 100707 9691 100773 9692
rect 102339 9280 102659 9840
rect 102339 9216 102347 9280
rect 102411 9216 102427 9280
rect 102491 9216 102507 9280
rect 102571 9216 102587 9280
rect 102651 9216 102659 9280
rect 99971 8668 100037 8669
rect 99971 8604 99972 8668
rect 100036 8604 100037 8668
rect 99971 8603 100037 8604
rect 99235 8260 99301 8261
rect 99235 8196 99236 8260
rect 99300 8196 99301 8260
rect 99235 8195 99301 8196
rect 102339 8192 102659 9216
rect 102339 8128 102347 8192
rect 102411 8128 102427 8192
rect 102491 8128 102507 8192
rect 102571 8128 102587 8192
rect 102651 8128 102659 8192
rect 88931 8124 88997 8125
rect 88931 8060 88932 8124
rect 88996 8060 88997 8124
rect 88931 8059 88997 8060
rect 68540 7584 68548 7648
rect 68612 7584 68628 7648
rect 68692 7584 68708 7648
rect 68772 7584 68788 7648
rect 68852 7584 68860 7648
rect 68540 6560 68860 7584
rect 68540 6496 68548 6560
rect 68612 6496 68628 6560
rect 68692 6496 68708 6560
rect 68772 6496 68788 6560
rect 68852 6496 68860 6560
rect 68540 5472 68860 6496
rect 68540 5408 68548 5472
rect 68612 5408 68628 5472
rect 68692 5408 68708 5472
rect 68772 5408 68788 5472
rect 68852 5408 68860 5472
rect 68540 4384 68860 5408
rect 68540 4320 68548 4384
rect 68612 4320 68628 4384
rect 68692 4320 68708 4384
rect 68772 4320 68788 4384
rect 68852 4320 68860 4384
rect 68540 3296 68860 4320
rect 68540 3232 68548 3296
rect 68612 3232 68628 3296
rect 68692 3232 68708 3296
rect 68772 3232 68788 3296
rect 68852 3232 68860 3296
rect 60043 2820 60109 2821
rect 60043 2756 60044 2820
rect 60108 2756 60109 2820
rect 60043 2755 60109 2756
rect 34742 2688 34750 2752
rect 34814 2688 34830 2752
rect 34894 2688 34910 2752
rect 34974 2688 34990 2752
rect 35054 2688 35062 2752
rect 34742 1664 35062 2688
rect 34742 1600 34750 1664
rect 34814 1600 34830 1664
rect 34894 1600 34910 1664
rect 34974 1600 34990 1664
rect 35054 1600 35062 1664
rect 32443 1460 32509 1461
rect 32443 1396 32444 1460
rect 32508 1396 32509 1460
rect 32443 1395 32509 1396
rect 25819 1324 25885 1325
rect 25819 1260 25820 1324
rect 25884 1260 25885 1324
rect 25819 1259 25885 1260
rect 26555 1324 26621 1325
rect 26555 1260 26556 1324
rect 26620 1260 26621 1324
rect 26555 1259 26621 1260
rect 27291 1324 27357 1325
rect 27291 1260 27292 1324
rect 27356 1260 27357 1324
rect 27291 1259 27357 1260
rect 25822 0 25882 1259
rect 26558 0 26618 1259
rect 27294 0 27354 1259
rect 28763 644 28829 645
rect 28763 580 28764 644
rect 28828 580 28829 644
rect 28763 579 28829 580
rect 30235 644 30301 645
rect 30235 580 30236 644
rect 30300 580 30301 644
rect 30235 579 30301 580
rect 28027 508 28093 509
rect 28027 444 28028 508
rect 28092 444 28093 508
rect 28027 443 28093 444
rect 28030 0 28090 443
rect 28766 0 28826 579
rect 29499 508 29565 509
rect 29499 444 29500 508
rect 29564 444 29565 508
rect 29499 443 29565 444
rect 29502 0 29562 443
rect 30238 0 30298 579
rect 31707 508 31773 509
rect 31707 444 31708 508
rect 31772 444 31773 508
rect 31707 443 31773 444
rect 30971 372 31037 373
rect 30971 308 30972 372
rect 31036 308 31037 372
rect 30971 307 31037 308
rect 30974 0 31034 307
rect 31710 0 31770 443
rect 32446 0 32506 1395
rect 34742 1040 35062 1600
rect 59307 1596 59373 1597
rect 59307 1532 59308 1596
rect 59372 1532 59373 1596
rect 59307 1531 59373 1532
rect 53971 1460 54037 1461
rect 53971 1396 53972 1460
rect 54036 1396 54037 1460
rect 53971 1395 54037 1396
rect 35663 644 35729 645
rect 35663 580 35664 644
rect 35728 580 35729 644
rect 35663 579 35729 580
rect 36399 644 36465 645
rect 36399 580 36400 644
rect 36464 580 36465 644
rect 36399 579 36465 580
rect 37135 644 37201 645
rect 37135 580 37136 644
rect 37200 580 37201 644
rect 37135 579 37201 580
rect 37871 644 37937 645
rect 37871 580 37872 644
rect 37936 580 37937 644
rect 37871 579 37937 580
rect 38607 644 38673 645
rect 38607 580 38608 644
rect 38672 580 38673 644
rect 38607 579 38673 580
rect 40079 644 40145 645
rect 40079 580 40080 644
rect 40144 580 40145 644
rect 40079 579 40145 580
rect 40815 644 40881 645
rect 40815 580 40816 644
rect 40880 580 40881 644
rect 40815 579 40881 580
rect 41551 644 41617 645
rect 41551 580 41552 644
rect 41616 580 41617 644
rect 41551 579 41617 580
rect 42287 644 42353 645
rect 42287 580 42288 644
rect 42352 580 42353 644
rect 42287 579 42353 580
rect 43023 644 43089 645
rect 43023 580 43024 644
rect 43088 580 43089 644
rect 43023 579 43089 580
rect 43759 644 43825 645
rect 43759 580 43760 644
rect 43824 580 43825 644
rect 43759 579 43825 580
rect 44495 644 44561 645
rect 44495 580 44496 644
rect 44560 580 44561 644
rect 44495 579 44561 580
rect 45231 644 45297 645
rect 45231 580 45232 644
rect 45296 580 45297 644
rect 45231 579 45297 580
rect 45967 644 46033 645
rect 45967 580 45968 644
rect 46032 580 46033 644
rect 45967 579 46033 580
rect 46703 644 46769 645
rect 46703 580 46704 644
rect 46768 580 46769 644
rect 46703 579 46769 580
rect 47439 644 47505 645
rect 47439 580 47440 644
rect 47504 580 47505 644
rect 47439 579 47505 580
rect 48175 644 48241 645
rect 48175 580 48176 644
rect 48240 580 48241 644
rect 48175 579 48241 580
rect 48911 644 48977 645
rect 48911 580 48912 644
rect 48976 580 48977 644
rect 48911 579 48977 580
rect 49647 644 49713 645
rect 49647 580 49648 644
rect 49712 580 49713 644
rect 49647 579 49713 580
rect 50383 644 50449 645
rect 50383 580 50384 644
rect 50448 580 50449 644
rect 50383 579 50449 580
rect 51119 644 51185 645
rect 51119 580 51120 644
rect 51184 580 51185 644
rect 51119 579 51185 580
rect 51855 644 51921 645
rect 51855 580 51856 644
rect 51920 580 51921 644
rect 51855 579 51921 580
rect 52591 644 52657 645
rect 52591 580 52592 644
rect 52656 580 52657 644
rect 52591 579 52657 580
rect 53327 644 53393 645
rect 53327 580 53328 644
rect 53392 580 53393 644
rect 53327 579 53393 580
rect 34927 372 34993 373
rect 34927 308 34928 372
rect 34992 308 34993 372
rect 34927 307 34993 308
rect 34930 0 34990 307
rect 35666 0 35726 579
rect 36402 0 36462 579
rect 37138 0 37198 579
rect 37874 0 37934 579
rect 38610 0 38670 579
rect 39343 372 39409 373
rect 39343 308 39344 372
rect 39408 308 39409 372
rect 39343 307 39409 308
rect 39346 0 39406 307
rect 40082 0 40142 579
rect 40818 0 40878 579
rect 41554 0 41614 579
rect 42290 0 42350 579
rect 43026 0 43086 579
rect 43762 0 43822 579
rect 44498 0 44558 579
rect 45234 0 45294 579
rect 45970 0 46030 579
rect 46706 0 46766 579
rect 47442 0 47502 579
rect 48178 0 48238 579
rect 48914 0 48974 579
rect 49650 0 49710 579
rect 50386 0 50446 579
rect 51122 0 51182 579
rect 51858 0 51918 579
rect 52594 0 52654 579
rect 53330 0 53390 579
rect 53974 370 54034 1395
rect 54799 644 54865 645
rect 54799 580 54800 644
rect 54864 580 54865 644
rect 54799 579 54865 580
rect 55535 644 55601 645
rect 55535 580 55536 644
rect 55600 580 55601 644
rect 55535 579 55601 580
rect 56271 644 56337 645
rect 56271 580 56272 644
rect 56336 580 56337 644
rect 56271 579 56337 580
rect 57007 644 57073 645
rect 57007 580 57008 644
rect 57072 580 57073 644
rect 57007 579 57073 580
rect 57743 644 57809 645
rect 57743 580 57744 644
rect 57808 580 57809 644
rect 57743 579 57809 580
rect 58479 644 58545 645
rect 58479 580 58480 644
rect 58544 580 58545 644
rect 58479 579 58545 580
rect 53974 310 54126 370
rect 54066 0 54126 310
rect 54802 0 54862 579
rect 55538 0 55598 579
rect 56274 0 56334 579
rect 57010 0 57070 579
rect 57746 0 57806 579
rect 58482 0 58542 579
rect 59310 370 59370 1531
rect 60046 370 60106 2755
rect 68540 2208 68860 3232
rect 68540 2144 68548 2208
rect 68612 2144 68628 2208
rect 68692 2144 68708 2208
rect 68772 2144 68788 2208
rect 68852 2144 68860 2208
rect 68540 1120 68860 2144
rect 102339 7104 102659 8128
rect 102339 7040 102347 7104
rect 102411 7040 102427 7104
rect 102491 7040 102507 7104
rect 102571 7040 102587 7104
rect 102651 7040 102659 7104
rect 102339 6016 102659 7040
rect 102339 5952 102347 6016
rect 102411 5952 102427 6016
rect 102491 5952 102507 6016
rect 102571 5952 102587 6016
rect 102651 5952 102659 6016
rect 102339 4928 102659 5952
rect 102339 4864 102347 4928
rect 102411 4864 102427 4928
rect 102491 4864 102507 4928
rect 102571 4864 102587 4928
rect 102651 4864 102659 4928
rect 102339 3840 102659 4864
rect 102339 3776 102347 3840
rect 102411 3776 102427 3840
rect 102491 3776 102507 3840
rect 102571 3776 102587 3840
rect 102651 3776 102659 3840
rect 102339 2752 102659 3776
rect 102339 2688 102347 2752
rect 102411 2688 102427 2752
rect 102491 2688 102507 2752
rect 102571 2688 102587 2752
rect 102651 2688 102659 2752
rect 102339 1664 102659 2688
rect 102339 1600 102347 1664
rect 102411 1600 102427 1664
rect 102491 1600 102507 1664
rect 102571 1600 102587 1664
rect 102651 1600 102659 1664
rect 80099 1596 80165 1597
rect 80099 1532 80100 1596
rect 80164 1532 80165 1596
rect 80099 1531 80165 1532
rect 81571 1596 81637 1597
rect 81571 1532 81572 1596
rect 81636 1532 81637 1596
rect 81571 1531 81637 1532
rect 83043 1596 83109 1597
rect 83043 1532 83044 1596
rect 83108 1532 83109 1596
rect 83043 1531 83109 1532
rect 83779 1596 83845 1597
rect 83779 1532 83780 1596
rect 83844 1532 83845 1596
rect 83779 1531 83845 1532
rect 99235 1596 99301 1597
rect 99235 1532 99236 1596
rect 99300 1532 99301 1596
rect 99235 1531 99301 1532
rect 71267 1324 71333 1325
rect 71267 1260 71268 1324
rect 71332 1260 71333 1324
rect 71267 1259 71333 1260
rect 73475 1324 73541 1325
rect 73475 1260 73476 1324
rect 73540 1260 73541 1324
rect 73475 1259 73541 1260
rect 76419 1324 76485 1325
rect 76419 1260 76420 1324
rect 76484 1260 76485 1324
rect 76419 1259 76485 1260
rect 77891 1324 77957 1325
rect 77891 1260 77892 1324
rect 77956 1260 77957 1324
rect 77891 1259 77957 1260
rect 79363 1324 79429 1325
rect 79363 1260 79364 1324
rect 79428 1260 79429 1324
rect 79363 1259 79429 1260
rect 68540 1056 68548 1120
rect 68612 1056 68628 1120
rect 68692 1056 68708 1120
rect 68772 1056 68788 1120
rect 68852 1056 68860 1120
rect 68540 1040 68860 1056
rect 70531 1052 70597 1053
rect 70531 988 70532 1052
rect 70596 988 70597 1052
rect 70531 987 70597 988
rect 69059 780 69125 781
rect 69059 716 69060 780
rect 69124 716 69125 780
rect 69059 715 69125 716
rect 69795 780 69861 781
rect 69795 716 69796 780
rect 69860 716 69861 780
rect 69795 715 69861 716
rect 60687 644 60753 645
rect 60687 580 60688 644
rect 60752 580 60753 644
rect 60687 579 60753 580
rect 61423 644 61489 645
rect 61423 580 61424 644
rect 61488 580 61489 644
rect 61423 579 61489 580
rect 62159 644 62225 645
rect 62159 580 62160 644
rect 62224 580 62225 644
rect 62159 579 62225 580
rect 62895 644 62961 645
rect 62895 580 62896 644
rect 62960 580 62961 644
rect 62895 579 62961 580
rect 63631 644 63697 645
rect 63631 580 63632 644
rect 63696 580 63697 644
rect 63631 579 63697 580
rect 64367 644 64433 645
rect 64367 580 64368 644
rect 64432 580 64433 644
rect 64367 579 64433 580
rect 65103 644 65169 645
rect 65103 580 65104 644
rect 65168 580 65169 644
rect 65103 579 65169 580
rect 59218 310 59370 370
rect 59954 310 60106 370
rect 59218 0 59278 310
rect 59954 0 60014 310
rect 60690 0 60750 579
rect 61426 0 61486 579
rect 62162 0 62222 579
rect 62898 0 62958 579
rect 63634 0 63694 579
rect 64370 0 64430 579
rect 65106 0 65166 579
rect 65839 508 65905 509
rect 65839 444 65840 508
rect 65904 444 65905 508
rect 65839 443 65905 444
rect 66575 508 66641 509
rect 66575 444 66576 508
rect 66640 444 66641 508
rect 66575 443 66641 444
rect 65842 0 65902 443
rect 66578 0 66638 443
rect 69062 0 69122 715
rect 69798 0 69858 715
rect 70534 0 70594 987
rect 71270 0 71330 1259
rect 72003 1052 72069 1053
rect 72003 988 72004 1052
rect 72068 988 72069 1052
rect 72003 987 72069 988
rect 72006 0 72066 987
rect 72739 644 72805 645
rect 72739 580 72740 644
rect 72804 580 72805 644
rect 72739 579 72805 580
rect 72742 0 72802 579
rect 73478 0 73538 1259
rect 74211 1052 74277 1053
rect 74211 988 74212 1052
rect 74276 988 74277 1052
rect 74211 987 74277 988
rect 75683 1052 75749 1053
rect 75683 988 75684 1052
rect 75748 988 75749 1052
rect 75683 987 75749 988
rect 74214 0 74274 987
rect 74947 644 75013 645
rect 74947 580 74948 644
rect 75012 580 75013 644
rect 74947 579 75013 580
rect 74950 0 75010 579
rect 75686 0 75746 987
rect 76422 0 76482 1259
rect 77155 1052 77221 1053
rect 77155 988 77156 1052
rect 77220 988 77221 1052
rect 77155 987 77221 988
rect 77158 0 77218 987
rect 77894 0 77954 1259
rect 78627 780 78693 781
rect 78627 716 78628 780
rect 78692 716 78693 780
rect 78627 715 78693 716
rect 78630 0 78690 715
rect 79366 0 79426 1259
rect 80102 0 80162 1531
rect 80835 780 80901 781
rect 80835 716 80836 780
rect 80900 716 80901 780
rect 80835 715 80901 716
rect 80838 0 80898 715
rect 81574 0 81634 1531
rect 82307 1324 82373 1325
rect 82307 1260 82308 1324
rect 82372 1260 82373 1324
rect 82307 1259 82373 1260
rect 82310 0 82370 1259
rect 83046 0 83106 1531
rect 83782 0 83842 1531
rect 87459 1324 87525 1325
rect 87459 1260 87460 1324
rect 87524 1260 87525 1324
rect 87459 1259 87525 1260
rect 88931 1324 88997 1325
rect 88931 1260 88932 1324
rect 88996 1260 88997 1324
rect 88931 1259 88997 1260
rect 85987 1052 86053 1053
rect 85987 988 85988 1052
rect 86052 988 86053 1052
rect 85987 987 86053 988
rect 84515 780 84581 781
rect 84515 716 84516 780
rect 84580 716 84581 780
rect 84515 715 84581 716
rect 85251 780 85317 781
rect 85251 716 85252 780
rect 85316 716 85317 780
rect 85251 715 85317 716
rect 84518 0 84578 715
rect 85254 0 85314 715
rect 85990 0 86050 987
rect 86723 780 86789 781
rect 86723 716 86724 780
rect 86788 716 86789 780
rect 86723 715 86789 716
rect 86726 0 86786 715
rect 87462 0 87522 1259
rect 88195 1188 88261 1189
rect 88195 1124 88196 1188
rect 88260 1124 88261 1188
rect 88195 1123 88261 1124
rect 88198 0 88258 1123
rect 88934 0 88994 1259
rect 94083 1188 94149 1189
rect 94083 1124 94084 1188
rect 94148 1124 94149 1188
rect 94083 1123 94149 1124
rect 94819 1188 94885 1189
rect 94819 1124 94820 1188
rect 94884 1124 94885 1188
rect 94819 1123 94885 1124
rect 95555 1188 95621 1189
rect 95555 1124 95556 1188
rect 95620 1124 95621 1188
rect 95555 1123 95621 1124
rect 96291 1188 96357 1189
rect 96291 1124 96292 1188
rect 96356 1124 96357 1188
rect 96291 1123 96357 1124
rect 90403 780 90469 781
rect 90403 716 90404 780
rect 90468 716 90469 780
rect 90403 715 90469 716
rect 91875 780 91941 781
rect 91875 716 91876 780
rect 91940 716 91941 780
rect 91875 715 91941 716
rect 93347 780 93413 781
rect 93347 716 93348 780
rect 93412 716 93413 780
rect 93347 715 93413 716
rect 89667 372 89733 373
rect 89667 308 89668 372
rect 89732 308 89733 372
rect 89667 307 89733 308
rect 89670 0 89730 307
rect 90406 0 90466 715
rect 91139 372 91205 373
rect 91139 308 91140 372
rect 91204 308 91205 372
rect 91139 307 91205 308
rect 91142 0 91202 307
rect 91878 0 91938 715
rect 92611 372 92677 373
rect 92611 308 92612 372
rect 92676 308 92677 372
rect 92611 307 92677 308
rect 92614 0 92674 307
rect 93350 0 93410 715
rect 94086 0 94146 1123
rect 94822 0 94882 1123
rect 95558 0 95618 1123
rect 96294 0 96354 1123
rect 97763 780 97829 781
rect 97763 716 97764 780
rect 97828 716 97829 780
rect 97763 715 97829 716
rect 98499 780 98565 781
rect 98499 716 98500 780
rect 98564 716 98565 780
rect 98499 715 98565 716
rect 97027 508 97093 509
rect 97027 444 97028 508
rect 97092 444 97093 508
rect 97027 443 97093 444
rect 97030 0 97090 443
rect 97766 0 97826 715
rect 98502 0 98562 715
rect 99238 0 99298 1531
rect 102339 1040 102659 1600
rect 136137 9824 136457 9840
rect 136137 9760 136145 9824
rect 136209 9760 136225 9824
rect 136289 9760 136305 9824
rect 136369 9760 136385 9824
rect 136449 9760 136457 9824
rect 136137 8736 136457 9760
rect 137326 9621 137386 10880
rect 138062 10301 138122 10880
rect 138059 10300 138125 10301
rect 138059 10236 138060 10300
rect 138124 10236 138125 10300
rect 138059 10235 138125 10236
rect 138798 10165 138858 10880
rect 138795 10164 138861 10165
rect 138795 10100 138796 10164
rect 138860 10100 138861 10164
rect 138795 10099 138861 10100
rect 139534 9893 139594 10880
rect 140270 10165 140330 10880
rect 141006 10165 141066 10880
rect 141742 10165 141802 10880
rect 142478 10301 142538 10880
rect 142475 10300 142541 10301
rect 142475 10236 142476 10300
rect 142540 10236 142541 10300
rect 142475 10235 142541 10236
rect 143214 10165 143274 10880
rect 143950 10165 144010 10880
rect 140267 10164 140333 10165
rect 140267 10100 140268 10164
rect 140332 10100 140333 10164
rect 140267 10099 140333 10100
rect 141003 10164 141069 10165
rect 141003 10100 141004 10164
rect 141068 10100 141069 10164
rect 141003 10099 141069 10100
rect 141739 10164 141805 10165
rect 141739 10100 141740 10164
rect 141804 10100 141805 10164
rect 141739 10099 141805 10100
rect 143211 10164 143277 10165
rect 143211 10100 143212 10164
rect 143276 10100 143277 10164
rect 143211 10099 143277 10100
rect 143947 10164 144013 10165
rect 143947 10100 143948 10164
rect 144012 10100 144013 10164
rect 143947 10099 144013 10100
rect 144686 9893 144746 10880
rect 145422 10165 145482 10880
rect 146158 10165 146218 10880
rect 146894 10165 146954 10880
rect 147630 10437 147690 10880
rect 147627 10436 147693 10437
rect 147627 10372 147628 10436
rect 147692 10372 147693 10436
rect 147627 10371 147693 10372
rect 148366 10165 148426 10880
rect 149102 10165 149162 10880
rect 145419 10164 145485 10165
rect 145419 10100 145420 10164
rect 145484 10100 145485 10164
rect 145419 10099 145485 10100
rect 146155 10164 146221 10165
rect 146155 10100 146156 10164
rect 146220 10100 146221 10164
rect 146155 10099 146221 10100
rect 146891 10164 146957 10165
rect 146891 10100 146892 10164
rect 146956 10100 146957 10164
rect 146891 10099 146957 10100
rect 148363 10164 148429 10165
rect 148363 10100 148364 10164
rect 148428 10100 148429 10164
rect 148363 10099 148429 10100
rect 149099 10164 149165 10165
rect 149099 10100 149100 10164
rect 149164 10100 149165 10164
rect 149099 10099 149165 10100
rect 149838 9893 149898 10880
rect 150574 10165 150634 10880
rect 151310 10165 151370 10880
rect 152046 10165 152106 10880
rect 152782 10165 152842 10880
rect 153518 10301 153578 10880
rect 153515 10300 153581 10301
rect 153515 10236 153516 10300
rect 153580 10236 153581 10300
rect 153515 10235 153581 10236
rect 154254 10165 154314 10880
rect 150571 10164 150637 10165
rect 150571 10100 150572 10164
rect 150636 10100 150637 10164
rect 150571 10099 150637 10100
rect 151307 10164 151373 10165
rect 151307 10100 151308 10164
rect 151372 10100 151373 10164
rect 151307 10099 151373 10100
rect 152043 10164 152109 10165
rect 152043 10100 152044 10164
rect 152108 10100 152109 10164
rect 152043 10099 152109 10100
rect 152779 10164 152845 10165
rect 152779 10100 152780 10164
rect 152844 10100 152845 10164
rect 152779 10099 152845 10100
rect 154251 10164 154317 10165
rect 154251 10100 154252 10164
rect 154316 10100 154317 10164
rect 154251 10099 154317 10100
rect 154990 9893 155050 10880
rect 139531 9892 139597 9893
rect 139531 9828 139532 9892
rect 139596 9828 139597 9892
rect 139531 9827 139597 9828
rect 144683 9892 144749 9893
rect 144683 9828 144684 9892
rect 144748 9828 144749 9892
rect 144683 9827 144749 9828
rect 149835 9892 149901 9893
rect 149835 9828 149836 9892
rect 149900 9828 149901 9892
rect 149835 9827 149901 9828
rect 154987 9892 155053 9893
rect 154987 9828 154988 9892
rect 155052 9828 155053 9892
rect 154987 9827 155053 9828
rect 155726 9757 155786 10880
rect 156462 9757 156522 10880
rect 157198 10301 157258 10880
rect 157195 10300 157261 10301
rect 157195 10236 157196 10300
rect 157260 10236 157261 10300
rect 157195 10235 157261 10236
rect 157934 9757 157994 10880
rect 155723 9756 155789 9757
rect 155723 9692 155724 9756
rect 155788 9692 155789 9756
rect 155723 9691 155789 9692
rect 156459 9756 156525 9757
rect 156459 9692 156460 9756
rect 156524 9692 156525 9756
rect 156459 9691 156525 9692
rect 157931 9756 157997 9757
rect 157931 9692 157932 9756
rect 157996 9692 157997 9756
rect 157931 9691 157997 9692
rect 137323 9620 137389 9621
rect 137323 9556 137324 9620
rect 137388 9556 137389 9620
rect 137323 9555 137389 9556
rect 158670 9485 158730 10880
rect 159406 9757 159466 10880
rect 159403 9756 159469 9757
rect 159403 9692 159404 9756
rect 159468 9692 159469 9756
rect 159403 9691 159469 9692
rect 158667 9484 158733 9485
rect 158667 9420 158668 9484
rect 158732 9420 158733 9484
rect 158667 9419 158733 9420
rect 136137 8672 136145 8736
rect 136209 8672 136225 8736
rect 136289 8672 136305 8736
rect 136369 8672 136385 8736
rect 136449 8672 136457 8736
rect 136137 7648 136457 8672
rect 160142 8397 160202 10880
rect 160878 8397 160938 10880
rect 161614 8533 161674 10880
rect 161611 8532 161677 8533
rect 161611 8468 161612 8532
rect 161676 8468 161677 8532
rect 161611 8467 161677 8468
rect 162350 8397 162410 10880
rect 163086 8397 163146 10880
rect 163822 9757 163882 10880
rect 163819 9756 163885 9757
rect 163819 9692 163820 9756
rect 163884 9692 163885 9756
rect 163819 9691 163885 9692
rect 164558 8397 164618 10880
rect 165294 8397 165354 10880
rect 166030 8397 166090 10880
rect 160139 8396 160205 8397
rect 160139 8332 160140 8396
rect 160204 8332 160205 8396
rect 160139 8331 160205 8332
rect 160875 8396 160941 8397
rect 160875 8332 160876 8396
rect 160940 8332 160941 8396
rect 160875 8331 160941 8332
rect 162347 8396 162413 8397
rect 162347 8332 162348 8396
rect 162412 8332 162413 8396
rect 162347 8331 162413 8332
rect 163083 8396 163149 8397
rect 163083 8332 163084 8396
rect 163148 8332 163149 8396
rect 163083 8331 163149 8332
rect 164555 8396 164621 8397
rect 164555 8332 164556 8396
rect 164620 8332 164621 8396
rect 164555 8331 164621 8332
rect 165291 8396 165357 8397
rect 165291 8332 165292 8396
rect 165356 8332 165357 8396
rect 165291 8331 165357 8332
rect 166027 8396 166093 8397
rect 166027 8332 166028 8396
rect 166092 8332 166093 8396
rect 166027 8331 166093 8332
rect 166766 8261 166826 10880
rect 167502 8397 167562 10880
rect 167499 8396 167565 8397
rect 167499 8332 167500 8396
rect 167564 8332 167565 8396
rect 167499 8331 167565 8332
rect 166763 8260 166829 8261
rect 166763 8196 166764 8260
rect 166828 8196 166829 8260
rect 166763 8195 166829 8196
rect 168238 8125 168298 10880
rect 168974 9213 169034 10880
rect 171458 10301 171518 10880
rect 172194 10301 172254 10880
rect 172930 10301 172990 10880
rect 173666 10301 173726 10880
rect 174402 10301 174462 10880
rect 175138 10301 175198 10880
rect 175874 10301 175934 10880
rect 176610 10301 176670 10880
rect 177346 10301 177406 10880
rect 178082 10301 178142 10880
rect 178818 10301 178878 10880
rect 179554 10301 179614 10880
rect 180290 10301 180350 10880
rect 181026 10301 181086 10880
rect 181762 10437 181822 10880
rect 181759 10436 181825 10437
rect 181759 10372 181760 10436
rect 181824 10372 181825 10436
rect 181759 10371 181825 10372
rect 182498 10301 182558 10880
rect 183234 10301 183294 10880
rect 183970 10301 184030 10880
rect 184706 10301 184766 10880
rect 185442 10301 185502 10880
rect 186178 10301 186238 10880
rect 186914 10301 186974 10880
rect 187650 10301 187710 10880
rect 188386 10301 188446 10880
rect 189122 10301 189182 10880
rect 189858 10301 189918 10880
rect 190594 10437 190654 10880
rect 190591 10436 190657 10437
rect 190591 10372 190592 10436
rect 190656 10372 190657 10436
rect 190591 10371 190657 10372
rect 191330 10301 191390 10880
rect 192066 10301 192126 10880
rect 192802 10301 192862 10880
rect 193538 10437 193598 10880
rect 193535 10436 193601 10437
rect 193535 10372 193536 10436
rect 193600 10372 193601 10436
rect 193535 10371 193601 10372
rect 194274 10301 194334 10880
rect 195010 10301 195070 10880
rect 195746 10301 195806 10880
rect 196482 10301 196542 10880
rect 197218 10301 197278 10880
rect 197954 10301 198014 10880
rect 198690 10437 198750 10880
rect 198687 10436 198753 10437
rect 198687 10372 198688 10436
rect 198752 10372 198753 10436
rect 198687 10371 198753 10372
rect 199426 10301 199486 10880
rect 200162 10301 200222 10880
rect 200898 10437 200958 10880
rect 200895 10436 200961 10437
rect 200895 10372 200896 10436
rect 200960 10372 200961 10436
rect 200895 10371 200961 10372
rect 201634 10301 201694 10880
rect 202370 10437 202430 10880
rect 202367 10436 202433 10437
rect 202367 10372 202368 10436
rect 202432 10372 202433 10436
rect 202367 10371 202433 10372
rect 203106 10301 203166 10880
rect 171455 10300 171521 10301
rect 171455 10236 171456 10300
rect 171520 10236 171521 10300
rect 171455 10235 171521 10236
rect 172191 10300 172257 10301
rect 172191 10236 172192 10300
rect 172256 10236 172257 10300
rect 172191 10235 172257 10236
rect 172927 10300 172993 10301
rect 172927 10236 172928 10300
rect 172992 10236 172993 10300
rect 172927 10235 172993 10236
rect 173663 10300 173729 10301
rect 173663 10236 173664 10300
rect 173728 10236 173729 10300
rect 173663 10235 173729 10236
rect 174399 10300 174465 10301
rect 174399 10236 174400 10300
rect 174464 10236 174465 10300
rect 174399 10235 174465 10236
rect 175135 10300 175201 10301
rect 175135 10236 175136 10300
rect 175200 10236 175201 10300
rect 175135 10235 175201 10236
rect 175871 10300 175937 10301
rect 175871 10236 175872 10300
rect 175936 10236 175937 10300
rect 175871 10235 175937 10236
rect 176607 10300 176673 10301
rect 176607 10236 176608 10300
rect 176672 10236 176673 10300
rect 176607 10235 176673 10236
rect 177343 10300 177409 10301
rect 177343 10236 177344 10300
rect 177408 10236 177409 10300
rect 177343 10235 177409 10236
rect 178079 10300 178145 10301
rect 178079 10236 178080 10300
rect 178144 10236 178145 10300
rect 178079 10235 178145 10236
rect 178815 10300 178881 10301
rect 178815 10236 178816 10300
rect 178880 10236 178881 10300
rect 178815 10235 178881 10236
rect 179551 10300 179617 10301
rect 179551 10236 179552 10300
rect 179616 10236 179617 10300
rect 179551 10235 179617 10236
rect 180287 10300 180353 10301
rect 180287 10236 180288 10300
rect 180352 10236 180353 10300
rect 180287 10235 180353 10236
rect 181023 10300 181089 10301
rect 181023 10236 181024 10300
rect 181088 10236 181089 10300
rect 181023 10235 181089 10236
rect 182495 10300 182561 10301
rect 182495 10236 182496 10300
rect 182560 10236 182561 10300
rect 182495 10235 182561 10236
rect 183231 10300 183297 10301
rect 183231 10236 183232 10300
rect 183296 10236 183297 10300
rect 183231 10235 183297 10236
rect 183967 10300 184033 10301
rect 183967 10236 183968 10300
rect 184032 10236 184033 10300
rect 183967 10235 184033 10236
rect 184703 10300 184769 10301
rect 184703 10236 184704 10300
rect 184768 10236 184769 10300
rect 184703 10235 184769 10236
rect 185439 10300 185505 10301
rect 185439 10236 185440 10300
rect 185504 10236 185505 10300
rect 185439 10235 185505 10236
rect 186175 10300 186241 10301
rect 186175 10236 186176 10300
rect 186240 10236 186241 10300
rect 186175 10235 186241 10236
rect 186911 10300 186977 10301
rect 186911 10236 186912 10300
rect 186976 10236 186977 10300
rect 186911 10235 186977 10236
rect 187647 10300 187713 10301
rect 187647 10236 187648 10300
rect 187712 10236 187713 10300
rect 187647 10235 187713 10236
rect 188383 10300 188449 10301
rect 188383 10236 188384 10300
rect 188448 10236 188449 10300
rect 188383 10235 188449 10236
rect 189119 10300 189185 10301
rect 189119 10236 189120 10300
rect 189184 10236 189185 10300
rect 189119 10235 189185 10236
rect 189855 10300 189921 10301
rect 189855 10236 189856 10300
rect 189920 10236 189921 10300
rect 189855 10235 189921 10236
rect 191327 10300 191393 10301
rect 191327 10236 191328 10300
rect 191392 10236 191393 10300
rect 191327 10235 191393 10236
rect 192063 10300 192129 10301
rect 192063 10236 192064 10300
rect 192128 10236 192129 10300
rect 192063 10235 192129 10236
rect 192799 10300 192865 10301
rect 192799 10236 192800 10300
rect 192864 10236 192865 10300
rect 192799 10235 192865 10236
rect 194271 10300 194337 10301
rect 194271 10236 194272 10300
rect 194336 10236 194337 10300
rect 194271 10235 194337 10236
rect 195007 10300 195073 10301
rect 195007 10236 195008 10300
rect 195072 10236 195073 10300
rect 195007 10235 195073 10236
rect 195743 10300 195809 10301
rect 195743 10236 195744 10300
rect 195808 10236 195809 10300
rect 195743 10235 195809 10236
rect 196479 10300 196545 10301
rect 196479 10236 196480 10300
rect 196544 10236 196545 10300
rect 196479 10235 196545 10236
rect 197215 10300 197281 10301
rect 197215 10236 197216 10300
rect 197280 10236 197281 10300
rect 197215 10235 197281 10236
rect 197951 10300 198017 10301
rect 197951 10236 197952 10300
rect 198016 10236 198017 10300
rect 197951 10235 198017 10236
rect 199423 10300 199489 10301
rect 199423 10236 199424 10300
rect 199488 10236 199489 10300
rect 199423 10235 199489 10236
rect 200159 10300 200225 10301
rect 200159 10236 200160 10300
rect 200224 10236 200225 10300
rect 200159 10235 200225 10236
rect 201631 10300 201697 10301
rect 201631 10236 201632 10300
rect 201696 10236 201697 10300
rect 201631 10235 201697 10236
rect 203103 10300 203169 10301
rect 203103 10236 203104 10300
rect 203168 10236 203169 10300
rect 203103 10235 203169 10236
rect 169936 9280 170256 9840
rect 169936 9216 169944 9280
rect 170008 9216 170024 9280
rect 170088 9216 170104 9280
rect 170168 9216 170184 9280
rect 170248 9216 170256 9280
rect 168971 9212 169037 9213
rect 168971 9148 168972 9212
rect 169036 9148 169037 9212
rect 168971 9147 169037 9148
rect 169936 8192 170256 9216
rect 169936 8128 169944 8192
rect 170008 8128 170024 8192
rect 170088 8128 170104 8192
rect 170168 8128 170184 8192
rect 170248 8128 170256 8192
rect 168235 8124 168301 8125
rect 168235 8060 168236 8124
rect 168300 8060 168301 8124
rect 168235 8059 168301 8060
rect 136137 7584 136145 7648
rect 136209 7584 136225 7648
rect 136289 7584 136305 7648
rect 136369 7584 136385 7648
rect 136449 7584 136457 7648
rect 136137 6560 136457 7584
rect 136137 6496 136145 6560
rect 136209 6496 136225 6560
rect 136289 6496 136305 6560
rect 136369 6496 136385 6560
rect 136449 6496 136457 6560
rect 136137 5472 136457 6496
rect 136137 5408 136145 5472
rect 136209 5408 136225 5472
rect 136289 5408 136305 5472
rect 136369 5408 136385 5472
rect 136449 5408 136457 5472
rect 136137 4384 136457 5408
rect 136137 4320 136145 4384
rect 136209 4320 136225 4384
rect 136289 4320 136305 4384
rect 136369 4320 136385 4384
rect 136449 4320 136457 4384
rect 136137 3296 136457 4320
rect 136137 3232 136145 3296
rect 136209 3232 136225 3296
rect 136289 3232 136305 3296
rect 136369 3232 136385 3296
rect 136449 3232 136457 3296
rect 136137 2208 136457 3232
rect 169936 7104 170256 8128
rect 169936 7040 169944 7104
rect 170008 7040 170024 7104
rect 170088 7040 170104 7104
rect 170168 7040 170184 7104
rect 170248 7040 170256 7104
rect 169936 6016 170256 7040
rect 169936 5952 169944 6016
rect 170008 5952 170024 6016
rect 170088 5952 170104 6016
rect 170168 5952 170184 6016
rect 170248 5952 170256 6016
rect 169936 4928 170256 5952
rect 169936 4864 169944 4928
rect 170008 4864 170024 4928
rect 170088 4864 170104 4928
rect 170168 4864 170184 4928
rect 170248 4864 170256 4928
rect 169936 3840 170256 4864
rect 169936 3776 169944 3840
rect 170008 3776 170024 3840
rect 170088 3776 170104 3840
rect 170168 3776 170184 3840
rect 170248 3776 170256 3840
rect 157195 2820 157261 2821
rect 157195 2756 157196 2820
rect 157260 2756 157261 2820
rect 157195 2755 157261 2756
rect 159403 2820 159469 2821
rect 159403 2756 159404 2820
rect 159468 2756 159469 2820
rect 159403 2755 159469 2756
rect 136137 2144 136145 2208
rect 136209 2144 136225 2208
rect 136289 2144 136305 2208
rect 136369 2144 136385 2208
rect 136449 2144 136457 2208
rect 117267 1460 117333 1461
rect 117267 1396 117268 1460
rect 117332 1396 117333 1460
rect 117267 1395 117333 1396
rect 128307 1460 128373 1461
rect 128307 1396 128308 1460
rect 128372 1396 128373 1460
rect 128307 1395 128373 1396
rect 134931 1460 134997 1461
rect 134931 1396 134932 1460
rect 134996 1396 134997 1460
rect 134931 1395 134997 1396
rect 100707 916 100773 917
rect 100707 852 100708 916
rect 100772 852 100773 916
rect 100707 851 100773 852
rect 99971 508 100037 509
rect 99971 444 99972 508
rect 100036 444 100037 508
rect 99971 443 100037 444
rect 99974 0 100034 443
rect 100710 0 100770 851
rect 114231 644 114297 645
rect 114231 580 114232 644
rect 114296 580 114297 644
rect 114231 579 114297 580
rect 114967 644 115033 645
rect 114967 580 114968 644
rect 115032 580 115033 644
rect 114967 579 115033 580
rect 115703 644 115769 645
rect 115703 580 115704 644
rect 115768 580 115769 644
rect 115703 579 115769 580
rect 116439 644 116505 645
rect 116439 580 116440 644
rect 116504 580 116505 644
rect 116439 579 116505 580
rect 103191 508 103257 509
rect 103191 444 103192 508
rect 103256 444 103257 508
rect 103191 443 103257 444
rect 103927 508 103993 509
rect 103927 444 103928 508
rect 103992 444 103993 508
rect 103927 443 103993 444
rect 104663 508 104729 509
rect 104663 444 104664 508
rect 104728 444 104729 508
rect 104663 443 104729 444
rect 105399 508 105465 509
rect 105399 444 105400 508
rect 105464 444 105465 508
rect 105399 443 105465 444
rect 106135 508 106201 509
rect 106135 444 106136 508
rect 106200 444 106201 508
rect 106135 443 106201 444
rect 106871 508 106937 509
rect 106871 444 106872 508
rect 106936 444 106937 508
rect 106871 443 106937 444
rect 107607 508 107673 509
rect 107607 444 107608 508
rect 107672 444 107673 508
rect 107607 443 107673 444
rect 108343 508 108409 509
rect 108343 444 108344 508
rect 108408 444 108409 508
rect 108343 443 108409 444
rect 109079 508 109145 509
rect 109079 444 109080 508
rect 109144 444 109145 508
rect 109079 443 109145 444
rect 109815 508 109881 509
rect 109815 444 109816 508
rect 109880 444 109881 508
rect 109815 443 109881 444
rect 110551 508 110617 509
rect 110551 444 110552 508
rect 110616 444 110617 508
rect 110551 443 110617 444
rect 111287 508 111353 509
rect 111287 444 111288 508
rect 111352 444 111353 508
rect 111287 443 111353 444
rect 112023 508 112089 509
rect 112023 444 112024 508
rect 112088 444 112089 508
rect 112023 443 112089 444
rect 112759 508 112825 509
rect 112759 444 112760 508
rect 112824 444 112825 508
rect 112759 443 112825 444
rect 103194 0 103254 443
rect 103930 0 103990 443
rect 104666 0 104726 443
rect 105402 0 105462 443
rect 106138 0 106198 443
rect 106874 0 106934 443
rect 107610 0 107670 443
rect 108346 0 108406 443
rect 109082 0 109142 443
rect 109818 0 109878 443
rect 110554 0 110614 443
rect 111290 0 111350 443
rect 112026 0 112086 443
rect 112762 0 112822 443
rect 113495 372 113561 373
rect 113495 308 113496 372
rect 113560 308 113561 372
rect 113495 307 113561 308
rect 113498 0 113558 307
rect 114234 0 114294 579
rect 114970 0 115030 579
rect 115706 0 115766 579
rect 116442 0 116502 579
rect 117270 370 117330 1395
rect 117911 644 117977 645
rect 117911 580 117912 644
rect 117976 580 117977 644
rect 117911 579 117977 580
rect 118647 644 118713 645
rect 118647 580 118648 644
rect 118712 580 118713 644
rect 118647 579 118713 580
rect 119383 644 119449 645
rect 119383 580 119384 644
rect 119448 580 119449 644
rect 119383 579 119449 580
rect 120119 644 120185 645
rect 120119 580 120120 644
rect 120184 580 120185 644
rect 120119 579 120185 580
rect 120855 644 120921 645
rect 120855 580 120856 644
rect 120920 580 120921 644
rect 120855 579 120921 580
rect 121591 644 121657 645
rect 121591 580 121592 644
rect 121656 580 121657 644
rect 121591 579 121657 580
rect 122327 644 122393 645
rect 122327 580 122328 644
rect 122392 580 122393 644
rect 122327 579 122393 580
rect 123063 644 123129 645
rect 123063 580 123064 644
rect 123128 580 123129 644
rect 123063 579 123129 580
rect 123799 644 123865 645
rect 123799 580 123800 644
rect 123864 580 123865 644
rect 123799 579 123865 580
rect 124535 644 124601 645
rect 124535 580 124536 644
rect 124600 580 124601 644
rect 124535 579 124601 580
rect 125271 644 125337 645
rect 125271 580 125272 644
rect 125336 580 125337 644
rect 125271 579 125337 580
rect 126007 644 126073 645
rect 126007 580 126008 644
rect 126072 580 126073 644
rect 126007 579 126073 580
rect 126743 644 126809 645
rect 126743 580 126744 644
rect 126808 580 126809 644
rect 126743 579 126809 580
rect 127479 644 127545 645
rect 127479 580 127480 644
rect 127544 580 127545 644
rect 127479 579 127545 580
rect 117178 310 117330 370
rect 117178 0 117238 310
rect 117914 0 117974 579
rect 118650 0 118710 579
rect 119386 0 119446 579
rect 120122 0 120182 579
rect 120858 0 120918 579
rect 121594 0 121654 579
rect 122330 0 122390 579
rect 123066 0 123126 579
rect 123802 0 123862 579
rect 124538 0 124598 579
rect 125274 0 125334 579
rect 126010 0 126070 579
rect 126746 0 126806 579
rect 127482 0 127542 579
rect 128310 370 128370 1395
rect 128951 644 129017 645
rect 128951 580 128952 644
rect 129016 580 129017 644
rect 128951 579 129017 580
rect 129687 644 129753 645
rect 129687 580 129688 644
rect 129752 580 129753 644
rect 129687 579 129753 580
rect 131159 644 131225 645
rect 131159 580 131160 644
rect 131224 580 131225 644
rect 131159 579 131225 580
rect 131895 644 131961 645
rect 131895 580 131896 644
rect 131960 580 131961 644
rect 131895 579 131961 580
rect 132631 644 132697 645
rect 132631 580 132632 644
rect 132696 580 132697 644
rect 132631 579 132697 580
rect 133367 644 133433 645
rect 133367 580 133368 644
rect 133432 580 133433 644
rect 133367 579 133433 580
rect 134103 644 134169 645
rect 134103 580 134104 644
rect 134168 580 134169 644
rect 134103 579 134169 580
rect 128218 310 128370 370
rect 128218 0 128278 310
rect 128954 0 129014 579
rect 129690 0 129750 579
rect 130423 372 130489 373
rect 130423 308 130424 372
rect 130488 308 130489 372
rect 130423 307 130489 308
rect 130426 0 130486 307
rect 131162 0 131222 579
rect 131898 0 131958 579
rect 132634 0 132694 579
rect 133370 0 133430 579
rect 134106 0 134166 579
rect 134934 370 134994 1395
rect 136137 1120 136457 2144
rect 137323 1460 137389 1461
rect 137323 1396 137324 1460
rect 137388 1396 137389 1460
rect 137323 1395 137389 1396
rect 144683 1460 144749 1461
rect 144683 1396 144684 1460
rect 144748 1396 144749 1460
rect 144683 1395 144749 1396
rect 155723 1460 155789 1461
rect 155723 1396 155724 1460
rect 155788 1396 155789 1460
rect 155723 1395 155789 1396
rect 156459 1460 156525 1461
rect 156459 1396 156460 1460
rect 156524 1396 156525 1460
rect 156459 1395 156525 1396
rect 136137 1056 136145 1120
rect 136209 1056 136225 1120
rect 136289 1056 136305 1120
rect 136369 1056 136385 1120
rect 136449 1056 136457 1120
rect 136137 1040 136457 1056
rect 134842 310 134994 370
rect 134842 0 134902 310
rect 137326 0 137386 1395
rect 140267 1324 140333 1325
rect 140267 1260 140268 1324
rect 140332 1260 140333 1324
rect 140267 1259 140333 1260
rect 138795 780 138861 781
rect 138795 716 138796 780
rect 138860 716 138861 780
rect 138795 715 138861 716
rect 138059 644 138125 645
rect 138059 580 138060 644
rect 138124 580 138125 644
rect 138059 579 138125 580
rect 138062 0 138122 579
rect 138798 0 138858 715
rect 139531 508 139597 509
rect 139531 444 139532 508
rect 139596 444 139597 508
rect 139531 443 139597 444
rect 139534 0 139594 443
rect 140270 0 140330 1259
rect 142475 1052 142541 1053
rect 142475 988 142476 1052
rect 142540 988 142541 1052
rect 142475 987 142541 988
rect 141003 780 141069 781
rect 141003 716 141004 780
rect 141068 716 141069 780
rect 141003 715 141069 716
rect 141006 0 141066 715
rect 141739 644 141805 645
rect 141739 580 141740 644
rect 141804 580 141805 644
rect 141739 579 141805 580
rect 141742 0 141802 579
rect 142478 0 142538 987
rect 143211 780 143277 781
rect 143211 716 143212 780
rect 143276 716 143277 780
rect 143211 715 143277 716
rect 143947 780 144013 781
rect 143947 716 143948 780
rect 144012 716 144013 780
rect 143947 715 144013 716
rect 143214 0 143274 715
rect 143950 0 144010 715
rect 144686 0 144746 1395
rect 154987 1324 155053 1325
rect 154987 1260 154988 1324
rect 155052 1260 155053 1324
rect 154987 1259 155053 1260
rect 149835 1052 149901 1053
rect 149835 988 149836 1052
rect 149900 988 149901 1052
rect 149835 987 149901 988
rect 145419 780 145485 781
rect 145419 716 145420 780
rect 145484 716 145485 780
rect 145419 715 145485 716
rect 146155 780 146221 781
rect 146155 716 146156 780
rect 146220 716 146221 780
rect 146155 715 146221 716
rect 146891 780 146957 781
rect 146891 716 146892 780
rect 146956 716 146957 780
rect 146891 715 146957 716
rect 148363 780 148429 781
rect 148363 716 148364 780
rect 148428 716 148429 780
rect 148363 715 148429 716
rect 149099 780 149165 781
rect 149099 716 149100 780
rect 149164 716 149165 780
rect 149099 715 149165 716
rect 145422 0 145482 715
rect 146158 0 146218 715
rect 146894 0 146954 715
rect 147627 644 147693 645
rect 147627 580 147628 644
rect 147692 580 147693 644
rect 147627 579 147693 580
rect 147630 0 147690 579
rect 148366 0 148426 715
rect 149102 0 149162 715
rect 149838 0 149898 987
rect 150571 780 150637 781
rect 150571 716 150572 780
rect 150636 716 150637 780
rect 150571 715 150637 716
rect 151307 780 151373 781
rect 151307 716 151308 780
rect 151372 716 151373 780
rect 151307 715 151373 716
rect 152043 780 152109 781
rect 152043 716 152044 780
rect 152108 716 152109 780
rect 152043 715 152109 716
rect 152779 780 152845 781
rect 152779 716 152780 780
rect 152844 716 152845 780
rect 152779 715 152845 716
rect 154251 780 154317 781
rect 154251 716 154252 780
rect 154316 716 154317 780
rect 154251 715 154317 716
rect 150574 0 150634 715
rect 151310 0 151370 715
rect 152046 0 152106 715
rect 152782 0 152842 715
rect 153515 644 153581 645
rect 153515 580 153516 644
rect 153580 580 153581 644
rect 153515 579 153581 580
rect 153518 0 153578 579
rect 154254 0 154314 715
rect 154990 0 155050 1259
rect 155726 0 155786 1395
rect 156462 0 156522 1395
rect 157198 0 157258 2755
rect 157931 1460 157997 1461
rect 157931 1396 157932 1460
rect 157996 1396 157997 1460
rect 157931 1395 157997 1396
rect 157934 0 157994 1395
rect 158667 644 158733 645
rect 158667 580 158668 644
rect 158732 580 158733 644
rect 158667 579 158733 580
rect 158670 0 158730 579
rect 159406 0 159466 2755
rect 169936 2752 170256 3776
rect 203734 9824 204054 9840
rect 203734 9760 203742 9824
rect 203806 9760 203822 9824
rect 203886 9760 203902 9824
rect 203966 9760 203982 9824
rect 204046 9760 204054 9824
rect 203734 8736 204054 9760
rect 205590 9621 205650 10880
rect 206326 10165 206386 10880
rect 207062 10165 207122 10880
rect 207798 10573 207858 10880
rect 207795 10572 207861 10573
rect 207795 10508 207796 10572
rect 207860 10508 207861 10572
rect 207795 10507 207861 10508
rect 208534 10165 208594 10880
rect 209270 10165 209330 10880
rect 210006 10437 210066 10880
rect 210003 10436 210069 10437
rect 210003 10372 210004 10436
rect 210068 10372 210069 10436
rect 210003 10371 210069 10372
rect 210742 10165 210802 10880
rect 211478 10437 211538 10880
rect 211475 10436 211541 10437
rect 211475 10372 211476 10436
rect 211540 10372 211541 10436
rect 211475 10371 211541 10372
rect 206323 10164 206389 10165
rect 206323 10100 206324 10164
rect 206388 10100 206389 10164
rect 206323 10099 206389 10100
rect 207059 10164 207125 10165
rect 207059 10100 207060 10164
rect 207124 10100 207125 10164
rect 207059 10099 207125 10100
rect 208531 10164 208597 10165
rect 208531 10100 208532 10164
rect 208596 10100 208597 10164
rect 208531 10099 208597 10100
rect 209267 10164 209333 10165
rect 209267 10100 209268 10164
rect 209332 10100 209333 10164
rect 209267 10099 209333 10100
rect 210739 10164 210805 10165
rect 210739 10100 210740 10164
rect 210804 10100 210805 10164
rect 210739 10099 210805 10100
rect 205587 9620 205653 9621
rect 205587 9556 205588 9620
rect 205652 9556 205653 9620
rect 205587 9555 205653 9556
rect 203734 8672 203742 8736
rect 203806 8672 203822 8736
rect 203886 8672 203902 8736
rect 203966 8672 203982 8736
rect 204046 8672 204054 8736
rect 203734 7648 204054 8672
rect 203734 7584 203742 7648
rect 203806 7584 203822 7648
rect 203886 7584 203902 7648
rect 203966 7584 203982 7648
rect 204046 7584 204054 7648
rect 203734 6560 204054 7584
rect 212214 6901 212274 10880
rect 212950 10165 213010 10880
rect 213686 10165 213746 10880
rect 214422 10165 214482 10880
rect 215158 10301 215218 10880
rect 215155 10300 215221 10301
rect 215155 10236 215156 10300
rect 215220 10236 215221 10300
rect 215155 10235 215221 10236
rect 215894 10165 215954 10880
rect 212947 10164 213013 10165
rect 212947 10100 212948 10164
rect 213012 10100 213013 10164
rect 212947 10099 213013 10100
rect 213683 10164 213749 10165
rect 213683 10100 213684 10164
rect 213748 10100 213749 10164
rect 213683 10099 213749 10100
rect 214419 10164 214485 10165
rect 214419 10100 214420 10164
rect 214484 10100 214485 10164
rect 214419 10099 214485 10100
rect 215891 10164 215957 10165
rect 215891 10100 215892 10164
rect 215956 10100 215957 10164
rect 215891 10099 215957 10100
rect 216630 9893 216690 10880
rect 217366 10165 217426 10880
rect 218102 10573 218162 10880
rect 218099 10572 218165 10573
rect 218099 10508 218100 10572
rect 218164 10508 218165 10572
rect 218099 10507 218165 10508
rect 218838 10165 218898 10880
rect 219574 10165 219634 10880
rect 220310 10301 220370 10880
rect 221046 10437 221106 10880
rect 221043 10436 221109 10437
rect 221043 10372 221044 10436
rect 221108 10372 221109 10436
rect 221043 10371 221109 10372
rect 221782 10301 221842 10880
rect 222518 10301 222578 10880
rect 220307 10300 220373 10301
rect 220307 10236 220308 10300
rect 220372 10236 220373 10300
rect 220307 10235 220373 10236
rect 221779 10300 221845 10301
rect 221779 10236 221780 10300
rect 221844 10236 221845 10300
rect 221779 10235 221845 10236
rect 222515 10300 222581 10301
rect 222515 10236 222516 10300
rect 222580 10236 222581 10300
rect 222515 10235 222581 10236
rect 223254 10165 223314 10880
rect 217363 10164 217429 10165
rect 217363 10100 217364 10164
rect 217428 10100 217429 10164
rect 217363 10099 217429 10100
rect 218835 10164 218901 10165
rect 218835 10100 218836 10164
rect 218900 10100 218901 10164
rect 218835 10099 218901 10100
rect 219571 10164 219637 10165
rect 219571 10100 219572 10164
rect 219636 10100 219637 10164
rect 219571 10099 219637 10100
rect 223251 10164 223317 10165
rect 223251 10100 223252 10164
rect 223316 10100 223317 10164
rect 223251 10099 223317 10100
rect 216627 9892 216693 9893
rect 216627 9828 216628 9892
rect 216692 9828 216693 9892
rect 216627 9827 216693 9828
rect 223990 9213 224050 10880
rect 223987 9212 224053 9213
rect 223987 9148 223988 9212
rect 224052 9148 224053 9212
rect 223987 9147 224053 9148
rect 224726 8397 224786 10880
rect 225462 9757 225522 10880
rect 225459 9756 225525 9757
rect 225459 9692 225460 9756
rect 225524 9692 225525 9756
rect 225459 9691 225525 9692
rect 226198 8669 226258 10880
rect 226934 8669 226994 10880
rect 227670 8669 227730 10880
rect 228406 9485 228466 10880
rect 228403 9484 228469 9485
rect 228403 9420 228404 9484
rect 228468 9420 228469 9484
rect 228403 9419 228469 9420
rect 229142 8669 229202 10880
rect 229878 9757 229938 10880
rect 229875 9756 229941 9757
rect 229875 9692 229876 9756
rect 229940 9692 229941 9756
rect 229875 9691 229941 9692
rect 226195 8668 226261 8669
rect 226195 8604 226196 8668
rect 226260 8604 226261 8668
rect 226195 8603 226261 8604
rect 226931 8668 226997 8669
rect 226931 8604 226932 8668
rect 226996 8604 226997 8668
rect 226931 8603 226997 8604
rect 227667 8668 227733 8669
rect 227667 8604 227668 8668
rect 227732 8604 227733 8668
rect 227667 8603 227733 8604
rect 229139 8668 229205 8669
rect 229139 8604 229140 8668
rect 229204 8604 229205 8668
rect 229139 8603 229205 8604
rect 230614 8397 230674 10880
rect 231350 9757 231410 10880
rect 231347 9756 231413 9757
rect 231347 9692 231348 9756
rect 231412 9692 231413 9756
rect 231347 9691 231413 9692
rect 232086 8669 232146 10880
rect 232822 8669 232882 10880
rect 233558 9757 233618 10880
rect 234294 9757 234354 10880
rect 235030 9757 235090 10880
rect 233555 9756 233621 9757
rect 233555 9692 233556 9756
rect 233620 9692 233621 9756
rect 233555 9691 233621 9692
rect 234291 9756 234357 9757
rect 234291 9692 234292 9756
rect 234356 9692 234357 9756
rect 234291 9691 234357 9692
rect 235027 9756 235093 9757
rect 235027 9692 235028 9756
rect 235092 9692 235093 9756
rect 235027 9691 235093 9692
rect 235766 9213 235826 10880
rect 235763 9212 235829 9213
rect 235763 9148 235764 9212
rect 235828 9148 235829 9212
rect 235763 9147 235829 9148
rect 236502 8669 236562 10880
rect 237238 9213 237298 10880
rect 239722 10301 239782 10880
rect 240458 10301 240518 10880
rect 241194 10301 241254 10880
rect 241930 10301 241990 10880
rect 242666 10301 242726 10880
rect 243402 10301 243462 10880
rect 244138 10301 244198 10880
rect 244874 10301 244934 10880
rect 245610 10301 245670 10880
rect 246346 10301 246406 10880
rect 247082 10301 247142 10880
rect 247818 10301 247878 10880
rect 248554 10301 248614 10880
rect 249290 10301 249350 10880
rect 250026 10301 250086 10880
rect 250762 10301 250822 10880
rect 251498 10301 251558 10880
rect 252234 10301 252294 10880
rect 252970 10301 253030 10880
rect 253706 10301 253766 10880
rect 254442 10301 254502 10880
rect 255178 10301 255238 10880
rect 255914 10301 255974 10880
rect 256650 10301 256710 10880
rect 257386 10301 257446 10880
rect 258122 10301 258182 10880
rect 258858 10301 258918 10880
rect 259594 10301 259654 10880
rect 260330 10301 260390 10880
rect 261066 10437 261126 10880
rect 261063 10436 261129 10437
rect 261063 10372 261064 10436
rect 261128 10372 261129 10436
rect 261063 10371 261129 10372
rect 261802 10301 261862 10880
rect 262538 10301 262598 10880
rect 263274 10301 263334 10880
rect 264010 10301 264070 10880
rect 264746 10437 264806 10880
rect 264743 10436 264809 10437
rect 264743 10372 264744 10436
rect 264808 10372 264809 10436
rect 264743 10371 264809 10372
rect 265482 10301 265542 10880
rect 266218 10570 266278 10880
rect 266126 10510 266278 10570
rect 239719 10300 239785 10301
rect 239719 10236 239720 10300
rect 239784 10236 239785 10300
rect 239719 10235 239785 10236
rect 240455 10300 240521 10301
rect 240455 10236 240456 10300
rect 240520 10236 240521 10300
rect 240455 10235 240521 10236
rect 241191 10300 241257 10301
rect 241191 10236 241192 10300
rect 241256 10236 241257 10300
rect 241191 10235 241257 10236
rect 241927 10300 241993 10301
rect 241927 10236 241928 10300
rect 241992 10236 241993 10300
rect 241927 10235 241993 10236
rect 242663 10300 242729 10301
rect 242663 10236 242664 10300
rect 242728 10236 242729 10300
rect 242663 10235 242729 10236
rect 243399 10300 243465 10301
rect 243399 10236 243400 10300
rect 243464 10236 243465 10300
rect 243399 10235 243465 10236
rect 244135 10300 244201 10301
rect 244135 10236 244136 10300
rect 244200 10236 244201 10300
rect 244135 10235 244201 10236
rect 244871 10300 244937 10301
rect 244871 10236 244872 10300
rect 244936 10236 244937 10300
rect 244871 10235 244937 10236
rect 245607 10300 245673 10301
rect 245607 10236 245608 10300
rect 245672 10236 245673 10300
rect 245607 10235 245673 10236
rect 246343 10300 246409 10301
rect 246343 10236 246344 10300
rect 246408 10236 246409 10300
rect 246343 10235 246409 10236
rect 247079 10300 247145 10301
rect 247079 10236 247080 10300
rect 247144 10236 247145 10300
rect 247079 10235 247145 10236
rect 247815 10300 247881 10301
rect 247815 10236 247816 10300
rect 247880 10236 247881 10300
rect 247815 10235 247881 10236
rect 248551 10300 248617 10301
rect 248551 10236 248552 10300
rect 248616 10236 248617 10300
rect 248551 10235 248617 10236
rect 249287 10300 249353 10301
rect 249287 10236 249288 10300
rect 249352 10236 249353 10300
rect 249287 10235 249353 10236
rect 250023 10300 250089 10301
rect 250023 10236 250024 10300
rect 250088 10236 250089 10300
rect 250023 10235 250089 10236
rect 250759 10300 250825 10301
rect 250759 10236 250760 10300
rect 250824 10236 250825 10300
rect 250759 10235 250825 10236
rect 251495 10300 251561 10301
rect 251495 10236 251496 10300
rect 251560 10236 251561 10300
rect 251495 10235 251561 10236
rect 252231 10300 252297 10301
rect 252231 10236 252232 10300
rect 252296 10236 252297 10300
rect 252231 10235 252297 10236
rect 252967 10300 253033 10301
rect 252967 10236 252968 10300
rect 253032 10236 253033 10300
rect 252967 10235 253033 10236
rect 253703 10300 253769 10301
rect 253703 10236 253704 10300
rect 253768 10236 253769 10300
rect 253703 10235 253769 10236
rect 254439 10300 254505 10301
rect 254439 10236 254440 10300
rect 254504 10236 254505 10300
rect 254439 10235 254505 10236
rect 255175 10300 255241 10301
rect 255175 10236 255176 10300
rect 255240 10236 255241 10300
rect 255175 10235 255241 10236
rect 255911 10300 255977 10301
rect 255911 10236 255912 10300
rect 255976 10236 255977 10300
rect 255911 10235 255977 10236
rect 256647 10300 256713 10301
rect 256647 10236 256648 10300
rect 256712 10236 256713 10300
rect 256647 10235 256713 10236
rect 257383 10300 257449 10301
rect 257383 10236 257384 10300
rect 257448 10236 257449 10300
rect 257383 10235 257449 10236
rect 258119 10300 258185 10301
rect 258119 10236 258120 10300
rect 258184 10236 258185 10300
rect 258119 10235 258185 10236
rect 258855 10300 258921 10301
rect 258855 10236 258856 10300
rect 258920 10236 258921 10300
rect 258855 10235 258921 10236
rect 259591 10300 259657 10301
rect 259591 10236 259592 10300
rect 259656 10236 259657 10300
rect 259591 10235 259657 10236
rect 260327 10300 260393 10301
rect 260327 10236 260328 10300
rect 260392 10236 260393 10300
rect 260327 10235 260393 10236
rect 261799 10300 261865 10301
rect 261799 10236 261800 10300
rect 261864 10236 261865 10300
rect 261799 10235 261865 10236
rect 262535 10300 262601 10301
rect 262535 10236 262536 10300
rect 262600 10236 262601 10300
rect 262535 10235 262601 10236
rect 263271 10300 263337 10301
rect 263271 10236 263272 10300
rect 263336 10236 263337 10300
rect 263271 10235 263337 10236
rect 264007 10300 264073 10301
rect 264007 10236 264008 10300
rect 264072 10236 264073 10300
rect 264007 10235 264073 10236
rect 265479 10300 265545 10301
rect 265479 10236 265480 10300
rect 265544 10236 265545 10300
rect 265479 10235 265545 10236
rect 237533 9280 237853 9840
rect 237533 9216 237541 9280
rect 237605 9216 237621 9280
rect 237685 9216 237701 9280
rect 237765 9216 237781 9280
rect 237845 9216 237853 9280
rect 237235 9212 237301 9213
rect 237235 9148 237236 9212
rect 237300 9148 237301 9212
rect 237235 9147 237301 9148
rect 232083 8668 232149 8669
rect 232083 8604 232084 8668
rect 232148 8604 232149 8668
rect 232083 8603 232149 8604
rect 232819 8668 232885 8669
rect 232819 8604 232820 8668
rect 232884 8604 232885 8668
rect 232819 8603 232885 8604
rect 236499 8668 236565 8669
rect 236499 8604 236500 8668
rect 236564 8604 236565 8668
rect 236499 8603 236565 8604
rect 224723 8396 224789 8397
rect 224723 8332 224724 8396
rect 224788 8332 224789 8396
rect 224723 8331 224789 8332
rect 230611 8396 230677 8397
rect 230611 8332 230612 8396
rect 230676 8332 230677 8396
rect 230611 8331 230677 8332
rect 237533 8192 237853 9216
rect 262075 8804 262141 8805
rect 262075 8740 262076 8804
rect 262140 8740 262141 8804
rect 262075 8739 262141 8740
rect 237533 8128 237541 8192
rect 237605 8128 237621 8192
rect 237685 8128 237701 8192
rect 237765 8128 237781 8192
rect 237845 8128 237853 8192
rect 237533 7104 237853 8128
rect 237533 7040 237541 7104
rect 237605 7040 237621 7104
rect 237685 7040 237701 7104
rect 237765 7040 237781 7104
rect 237845 7040 237853 7104
rect 212211 6900 212277 6901
rect 212211 6836 212212 6900
rect 212276 6836 212277 6900
rect 212211 6835 212277 6836
rect 216627 6628 216693 6629
rect 216627 6564 216628 6628
rect 216692 6564 216693 6628
rect 216627 6563 216693 6564
rect 203734 6496 203742 6560
rect 203806 6496 203822 6560
rect 203886 6496 203902 6560
rect 203966 6496 203982 6560
rect 204046 6496 204054 6560
rect 203734 5472 204054 6496
rect 203734 5408 203742 5472
rect 203806 5408 203822 5472
rect 203886 5408 203902 5472
rect 203966 5408 203982 5472
rect 204046 5408 204054 5472
rect 203734 4384 204054 5408
rect 203734 4320 203742 4384
rect 203806 4320 203822 4384
rect 203886 4320 203902 4384
rect 203966 4320 203982 4384
rect 204046 4320 204054 4384
rect 203734 3296 204054 4320
rect 215339 3772 215405 3773
rect 215339 3708 215340 3772
rect 215404 3708 215405 3772
rect 215339 3707 215405 3708
rect 203734 3232 203742 3296
rect 203806 3232 203822 3296
rect 203886 3232 203902 3296
rect 203966 3232 203982 3296
rect 204046 3232 204054 3296
rect 189947 2820 190013 2821
rect 189947 2756 189948 2820
rect 190012 2756 190013 2820
rect 189947 2755 190013 2756
rect 191419 2820 191485 2821
rect 191419 2756 191420 2820
rect 191484 2756 191485 2820
rect 191419 2755 191485 2756
rect 202459 2820 202525 2821
rect 202459 2756 202460 2820
rect 202524 2756 202525 2820
rect 202459 2755 202525 2756
rect 169936 2688 169944 2752
rect 170008 2688 170024 2752
rect 170088 2688 170104 2752
rect 170168 2688 170184 2752
rect 170248 2688 170256 2752
rect 169936 1664 170256 2688
rect 169936 1600 169944 1664
rect 170008 1600 170024 1664
rect 170088 1600 170104 1664
rect 170168 1600 170184 1664
rect 170248 1600 170256 1664
rect 163819 1460 163885 1461
rect 163819 1396 163820 1460
rect 163884 1396 163885 1460
rect 163819 1395 163885 1396
rect 168235 1460 168301 1461
rect 168235 1396 168236 1460
rect 168300 1396 168301 1460
rect 168235 1395 168301 1396
rect 160139 1188 160205 1189
rect 160139 1124 160140 1188
rect 160204 1124 160205 1188
rect 160139 1123 160205 1124
rect 161611 1188 161677 1189
rect 161611 1124 161612 1188
rect 161676 1124 161677 1188
rect 161611 1123 161677 1124
rect 163083 1188 163149 1189
rect 163083 1124 163084 1188
rect 163148 1124 163149 1188
rect 163083 1123 163149 1124
rect 160142 0 160202 1123
rect 160875 644 160941 645
rect 160875 580 160876 644
rect 160940 580 160941 644
rect 160875 579 160941 580
rect 160878 0 160938 579
rect 161614 0 161674 1123
rect 162347 644 162413 645
rect 162347 580 162348 644
rect 162412 580 162413 644
rect 162347 579 162413 580
rect 162350 0 162410 579
rect 163086 0 163146 1123
rect 163822 0 163882 1395
rect 165291 1188 165357 1189
rect 165291 1124 165292 1188
rect 165356 1124 165357 1188
rect 165291 1123 165357 1124
rect 166027 1188 166093 1189
rect 166027 1124 166028 1188
rect 166092 1124 166093 1188
rect 166027 1123 166093 1124
rect 166763 1188 166829 1189
rect 166763 1124 166764 1188
rect 166828 1124 166829 1188
rect 166763 1123 166829 1124
rect 164555 644 164621 645
rect 164555 580 164556 644
rect 164620 580 164621 644
rect 164555 579 164621 580
rect 164558 0 164618 579
rect 165294 0 165354 1123
rect 166030 0 166090 1123
rect 166766 0 166826 1123
rect 167499 644 167565 645
rect 167499 580 167500 644
rect 167564 580 167565 644
rect 167499 579 167565 580
rect 167502 0 167562 579
rect 168238 0 168298 1395
rect 169936 1040 170256 1600
rect 186267 1460 186333 1461
rect 186267 1396 186268 1460
rect 186332 1396 186333 1460
rect 186267 1395 186333 1396
rect 176699 1324 176765 1325
rect 176699 1260 176700 1324
rect 176764 1260 176765 1324
rect 176699 1259 176765 1260
rect 179643 1324 179709 1325
rect 179643 1260 179644 1324
rect 179708 1260 179709 1324
rect 179643 1259 179709 1260
rect 181851 1324 181917 1325
rect 181851 1260 181852 1324
rect 181916 1260 181917 1324
rect 181851 1259 181917 1260
rect 171547 916 171613 917
rect 171547 852 171548 916
rect 171612 852 171613 916
rect 171547 851 171613 852
rect 172283 916 172349 917
rect 172283 852 172284 916
rect 172348 852 172349 916
rect 172283 851 172349 852
rect 173019 916 173085 917
rect 173019 852 173020 916
rect 173084 852 173085 916
rect 173019 851 173085 852
rect 173755 916 173821 917
rect 173755 852 173756 916
rect 173820 852 173821 916
rect 173755 851 173821 852
rect 174491 916 174557 917
rect 174491 852 174492 916
rect 174556 852 174557 916
rect 174491 851 174557 852
rect 175227 916 175293 917
rect 175227 852 175228 916
rect 175292 852 175293 916
rect 175227 851 175293 852
rect 175963 916 176029 917
rect 175963 852 175964 916
rect 176028 852 176029 916
rect 175963 851 176029 852
rect 168971 644 169037 645
rect 168971 580 168972 644
rect 169036 580 169037 644
rect 168971 579 169037 580
rect 168974 0 169034 579
rect 171550 370 171610 851
rect 172286 370 172346 851
rect 173022 370 173082 851
rect 173758 370 173818 851
rect 174494 370 174554 851
rect 175230 370 175290 851
rect 175966 370 176026 851
rect 176702 370 176762 1259
rect 177435 916 177501 917
rect 177435 852 177436 916
rect 177500 852 177501 916
rect 177435 851 177501 852
rect 178171 916 178237 917
rect 178171 852 178172 916
rect 178236 852 178237 916
rect 178171 851 178237 852
rect 178907 916 178973 917
rect 178907 852 178908 916
rect 178972 852 178973 916
rect 178907 851 178973 852
rect 177438 370 177498 851
rect 178174 370 178234 851
rect 178910 370 178970 851
rect 179646 370 179706 1259
rect 180379 916 180445 917
rect 180379 852 180380 916
rect 180444 852 180445 916
rect 180379 851 180445 852
rect 181115 916 181181 917
rect 181115 852 181116 916
rect 181180 852 181181 916
rect 181115 851 181181 852
rect 180382 370 180442 851
rect 181118 370 181178 851
rect 181854 370 181914 1259
rect 183323 1052 183389 1053
rect 183323 988 183324 1052
rect 183388 988 183389 1052
rect 183323 987 183389 988
rect 184795 1052 184861 1053
rect 184795 988 184796 1052
rect 184860 988 184861 1052
rect 184795 987 184861 988
rect 182587 916 182653 917
rect 182587 852 182588 916
rect 182652 852 182653 916
rect 182587 851 182653 852
rect 182590 370 182650 851
rect 183326 370 183386 987
rect 184059 916 184125 917
rect 184059 852 184060 916
rect 184124 852 184125 916
rect 184059 851 184125 852
rect 184062 370 184122 851
rect 184798 370 184858 987
rect 185531 916 185597 917
rect 185531 852 185532 916
rect 185596 852 185597 916
rect 185531 851 185597 852
rect 185534 370 185594 851
rect 186270 370 186330 1395
rect 187003 1324 187069 1325
rect 187003 1260 187004 1324
rect 187068 1260 187069 1324
rect 187003 1259 187069 1260
rect 187006 370 187066 1259
rect 187739 1052 187805 1053
rect 187739 988 187740 1052
rect 187804 988 187805 1052
rect 187739 987 187805 988
rect 189211 1052 189277 1053
rect 189211 988 189212 1052
rect 189276 988 189277 1052
rect 189211 987 189277 988
rect 187742 370 187802 987
rect 188475 916 188541 917
rect 188475 852 188476 916
rect 188540 852 188541 916
rect 188475 851 188541 852
rect 188478 370 188538 851
rect 189214 370 189274 987
rect 189950 370 190010 2755
rect 190683 1188 190749 1189
rect 190683 1124 190684 1188
rect 190748 1124 190749 1188
rect 190683 1123 190749 1124
rect 190686 370 190746 1123
rect 191422 370 191482 2755
rect 201723 1596 201789 1597
rect 201723 1532 201724 1596
rect 201788 1532 201789 1596
rect 201723 1531 201789 1532
rect 194363 1460 194429 1461
rect 194363 1396 194364 1460
rect 194428 1396 194429 1460
rect 194363 1395 194429 1396
rect 195835 1460 195901 1461
rect 195835 1396 195836 1460
rect 195900 1396 195901 1460
rect 195835 1395 195901 1396
rect 192155 916 192221 917
rect 192155 852 192156 916
rect 192220 852 192221 916
rect 192155 851 192221 852
rect 192891 916 192957 917
rect 192891 852 192892 916
rect 192956 852 192957 916
rect 192891 851 192957 852
rect 193627 916 193693 917
rect 193627 852 193628 916
rect 193692 852 193693 916
rect 193627 851 193693 852
rect 192158 370 192218 851
rect 192894 370 192954 851
rect 193630 370 193690 851
rect 194366 370 194426 1395
rect 195099 916 195165 917
rect 195099 852 195100 916
rect 195164 852 195165 916
rect 195099 851 195165 852
rect 195102 370 195162 851
rect 195838 370 195898 1395
rect 199515 1324 199581 1325
rect 199515 1260 199516 1324
rect 199580 1260 199581 1324
rect 199515 1259 199581 1260
rect 198043 1188 198109 1189
rect 198043 1124 198044 1188
rect 198108 1124 198109 1188
rect 198043 1123 198109 1124
rect 196571 916 196637 917
rect 196571 852 196572 916
rect 196636 852 196637 916
rect 196571 851 196637 852
rect 197307 916 197373 917
rect 197307 852 197308 916
rect 197372 852 197373 916
rect 197307 851 197373 852
rect 196574 370 196634 851
rect 197310 370 197370 851
rect 198046 370 198106 1123
rect 198779 916 198845 917
rect 198779 852 198780 916
rect 198844 852 198845 916
rect 198779 851 198845 852
rect 198782 370 198842 851
rect 199518 370 199578 1259
rect 200987 1188 201053 1189
rect 200987 1124 200988 1188
rect 201052 1124 201053 1188
rect 200987 1123 201053 1124
rect 200251 916 200317 917
rect 200251 852 200252 916
rect 200316 852 200317 916
rect 200251 851 200317 852
rect 200254 370 200314 851
rect 200990 370 201050 1123
rect 201726 370 201786 1531
rect 202462 370 202522 2755
rect 203734 2208 204054 3232
rect 203734 2144 203742 2208
rect 203806 2144 203822 2208
rect 203886 2144 203902 2208
rect 203966 2144 203982 2208
rect 204046 2144 204054 2208
rect 203734 1120 204054 2144
rect 215342 1733 215402 3707
rect 216630 2413 216690 6563
rect 237533 6016 237853 7040
rect 262078 6221 262138 8739
rect 263179 8396 263245 8397
rect 263179 8332 263180 8396
rect 263244 8332 263245 8396
rect 263179 8331 263245 8332
rect 262075 6220 262141 6221
rect 262075 6156 262076 6220
rect 262140 6156 262141 6220
rect 262075 6155 262141 6156
rect 237533 5952 237541 6016
rect 237605 5952 237621 6016
rect 237685 5952 237701 6016
rect 237765 5952 237781 6016
rect 237845 5952 237853 6016
rect 230611 5540 230677 5541
rect 230611 5476 230612 5540
rect 230676 5476 230677 5540
rect 230611 5475 230677 5476
rect 230614 5133 230674 5475
rect 230611 5132 230677 5133
rect 230611 5068 230612 5132
rect 230676 5068 230677 5132
rect 230611 5067 230677 5068
rect 237533 4928 237853 5952
rect 263182 5269 263242 8331
rect 266126 6765 266186 10510
rect 266954 10298 267014 10880
rect 266862 10238 267014 10298
rect 267690 10298 267750 10880
rect 268426 10298 268486 10880
rect 267690 10238 267842 10298
rect 266491 8396 266557 8397
rect 266491 8332 266492 8396
rect 266556 8332 266557 8396
rect 266491 8331 266557 8332
rect 266123 6764 266189 6765
rect 266123 6700 266124 6764
rect 266188 6700 266189 6764
rect 266123 6699 266189 6700
rect 263179 5268 263245 5269
rect 263179 5204 263180 5268
rect 263244 5204 263245 5268
rect 263179 5203 263245 5204
rect 237533 4864 237541 4928
rect 237605 4864 237621 4928
rect 237685 4864 237701 4928
rect 237765 4864 237781 4928
rect 237845 4864 237853 4928
rect 237533 3840 237853 4864
rect 237533 3776 237541 3840
rect 237605 3776 237621 3840
rect 237685 3776 237701 3840
rect 237765 3776 237781 3840
rect 237845 3776 237853 3840
rect 223251 2820 223317 2821
rect 223251 2756 223252 2820
rect 223316 2756 223317 2820
rect 223251 2755 223317 2756
rect 224723 2820 224789 2821
rect 224723 2756 224724 2820
rect 224788 2756 224789 2820
rect 224723 2755 224789 2756
rect 226195 2820 226261 2821
rect 226195 2756 226196 2820
rect 226260 2756 226261 2820
rect 226195 2755 226261 2756
rect 235763 2820 235829 2821
rect 235763 2756 235764 2820
rect 235828 2756 235829 2820
rect 235763 2755 235829 2756
rect 216627 2412 216693 2413
rect 216627 2348 216628 2412
rect 216692 2348 216693 2412
rect 216627 2347 216693 2348
rect 215339 1732 215405 1733
rect 215339 1668 215340 1732
rect 215404 1668 215405 1732
rect 215339 1667 215405 1668
rect 216627 1460 216693 1461
rect 216627 1396 216628 1460
rect 216692 1396 216693 1460
rect 216627 1395 216693 1396
rect 220307 1460 220373 1461
rect 220307 1396 220308 1460
rect 220372 1396 220373 1460
rect 220307 1395 220373 1396
rect 210739 1324 210805 1325
rect 210739 1260 210740 1324
rect 210804 1260 210805 1324
rect 210739 1259 210805 1260
rect 203734 1056 203742 1120
rect 203806 1056 203822 1120
rect 203886 1056 203902 1120
rect 203966 1056 203982 1120
rect 204046 1056 204054 1120
rect 203734 1040 204054 1056
rect 210003 1052 210069 1053
rect 210003 988 210004 1052
rect 210068 988 210069 1052
rect 210003 987 210069 988
rect 203195 916 203261 917
rect 203195 852 203196 916
rect 203260 852 203261 916
rect 203195 851 203261 852
rect 205771 916 205837 917
rect 205771 852 205772 916
rect 205836 852 205837 916
rect 205771 851 205837 852
rect 206323 916 206389 917
rect 206323 852 206324 916
rect 206388 852 206389 916
rect 206323 851 206389 852
rect 207059 916 207125 917
rect 207059 852 207060 916
rect 207124 852 207125 916
rect 207059 851 207125 852
rect 207795 916 207861 917
rect 207795 852 207796 916
rect 207860 852 207861 916
rect 207795 851 207861 852
rect 208531 916 208597 917
rect 208531 852 208532 916
rect 208596 852 208597 916
rect 208531 851 208597 852
rect 209267 916 209333 917
rect 209267 852 209268 916
rect 209332 852 209333 916
rect 209267 851 209333 852
rect 203198 370 203258 851
rect 205774 370 205834 851
rect 171458 310 171610 370
rect 172194 310 172346 370
rect 172930 310 173082 370
rect 173666 310 173818 370
rect 174402 310 174554 370
rect 175138 310 175290 370
rect 175874 310 176026 370
rect 176610 310 176762 370
rect 177346 310 177498 370
rect 178082 310 178234 370
rect 178818 310 178970 370
rect 179554 310 179706 370
rect 180290 310 180442 370
rect 181026 310 181178 370
rect 181762 310 181914 370
rect 182498 310 182650 370
rect 183234 310 183386 370
rect 183970 310 184122 370
rect 184706 310 184858 370
rect 185442 310 185594 370
rect 186178 310 186330 370
rect 186914 310 187066 370
rect 187650 310 187802 370
rect 188386 310 188538 370
rect 189122 310 189274 370
rect 189858 310 190010 370
rect 190594 310 190746 370
rect 191330 310 191482 370
rect 192066 310 192218 370
rect 192802 310 192954 370
rect 193538 310 193690 370
rect 194274 310 194426 370
rect 195010 310 195162 370
rect 195746 310 195898 370
rect 196482 310 196634 370
rect 197218 310 197370 370
rect 197954 310 198106 370
rect 198690 310 198842 370
rect 199426 310 199578 370
rect 200162 310 200314 370
rect 200898 310 201050 370
rect 201634 310 201786 370
rect 202370 310 202522 370
rect 203106 310 203258 370
rect 205590 310 205834 370
rect 171458 0 171518 310
rect 172194 0 172254 310
rect 172930 0 172990 310
rect 173666 0 173726 310
rect 174402 0 174462 310
rect 175138 0 175198 310
rect 175874 0 175934 310
rect 176610 0 176670 310
rect 177346 0 177406 310
rect 178082 0 178142 310
rect 178818 0 178878 310
rect 179554 0 179614 310
rect 180290 0 180350 310
rect 181026 0 181086 310
rect 181762 0 181822 310
rect 182498 0 182558 310
rect 183234 0 183294 310
rect 183970 0 184030 310
rect 184706 0 184766 310
rect 185442 0 185502 310
rect 186178 0 186238 310
rect 186914 0 186974 310
rect 187650 0 187710 310
rect 188386 0 188446 310
rect 189122 0 189182 310
rect 189858 0 189918 310
rect 190594 0 190654 310
rect 191330 0 191390 310
rect 192066 0 192126 310
rect 192802 0 192862 310
rect 193538 0 193598 310
rect 194274 0 194334 310
rect 195010 0 195070 310
rect 195746 0 195806 310
rect 196482 0 196542 310
rect 197218 0 197278 310
rect 197954 0 198014 310
rect 198690 0 198750 310
rect 199426 0 199486 310
rect 200162 0 200222 310
rect 200898 0 200958 310
rect 201634 0 201694 310
rect 202370 0 202430 310
rect 203106 0 203166 310
rect 205590 0 205650 310
rect 206326 0 206386 851
rect 207062 0 207122 851
rect 207798 0 207858 851
rect 208534 0 208594 851
rect 209270 0 209330 851
rect 210006 0 210066 987
rect 210742 0 210802 1259
rect 211475 1052 211541 1053
rect 211475 988 211476 1052
rect 211540 988 211541 1052
rect 211475 987 211541 988
rect 211478 0 211538 987
rect 212211 916 212277 917
rect 212211 852 212212 916
rect 212276 852 212277 916
rect 212211 851 212277 852
rect 212947 916 213013 917
rect 212947 852 212948 916
rect 213012 852 213013 916
rect 212947 851 213013 852
rect 213683 916 213749 917
rect 213683 852 213684 916
rect 213748 852 213749 916
rect 213683 851 213749 852
rect 214419 916 214485 917
rect 214419 852 214420 916
rect 214484 852 214485 916
rect 214419 851 214485 852
rect 215155 916 215221 917
rect 215155 852 215156 916
rect 215220 852 215221 916
rect 215155 851 215221 852
rect 215891 916 215957 917
rect 215891 852 215892 916
rect 215956 852 215957 916
rect 215891 851 215957 852
rect 212214 0 212274 851
rect 212950 0 213010 851
rect 213686 0 213746 851
rect 214422 0 214482 851
rect 215158 0 215218 851
rect 215894 0 215954 851
rect 216630 0 216690 1395
rect 217363 916 217429 917
rect 217363 852 217364 916
rect 217428 852 217429 916
rect 217363 851 217429 852
rect 218099 916 218165 917
rect 218099 852 218100 916
rect 218164 852 218165 916
rect 218099 851 218165 852
rect 217366 0 217426 851
rect 218102 0 218162 851
rect 218835 372 218901 373
rect 218835 308 218836 372
rect 218900 308 218901 372
rect 218835 307 218901 308
rect 219571 372 219637 373
rect 219571 308 219572 372
rect 219636 308 219637 372
rect 219571 307 219637 308
rect 218838 0 218898 307
rect 219574 0 219634 307
rect 220310 0 220370 1395
rect 222515 1324 222581 1325
rect 222515 1260 222516 1324
rect 222580 1260 222581 1324
rect 222515 1259 222581 1260
rect 221043 916 221109 917
rect 221043 852 221044 916
rect 221108 852 221109 916
rect 221043 851 221109 852
rect 221046 0 221106 851
rect 221779 372 221845 373
rect 221779 308 221780 372
rect 221844 308 221845 372
rect 221779 307 221845 308
rect 221782 0 221842 307
rect 222518 0 222578 1259
rect 223254 0 223314 2755
rect 223619 2548 223685 2549
rect 223619 2484 223620 2548
rect 223684 2484 223685 2548
rect 223619 2483 223685 2484
rect 223622 2410 223682 2483
rect 223622 2350 224234 2410
rect 224174 2277 224234 2350
rect 224171 2276 224237 2277
rect 224171 2212 224172 2276
rect 224236 2212 224237 2276
rect 224171 2211 224237 2212
rect 223987 1460 224053 1461
rect 223987 1396 223988 1460
rect 224052 1396 224053 1460
rect 223987 1395 224053 1396
rect 223990 0 224050 1395
rect 224726 0 224786 2755
rect 225459 1460 225525 1461
rect 225459 1396 225460 1460
rect 225524 1396 225525 1460
rect 225459 1395 225525 1396
rect 225462 0 225522 1395
rect 226198 0 226258 2755
rect 226931 1324 226997 1325
rect 226931 1260 226932 1324
rect 226996 1260 226997 1324
rect 226931 1259 226997 1260
rect 227667 1324 227733 1325
rect 227667 1260 227668 1324
rect 227732 1260 227733 1324
rect 227667 1259 227733 1260
rect 226934 0 226994 1259
rect 227670 0 227730 1259
rect 228403 1188 228469 1189
rect 228403 1124 228404 1188
rect 228468 1124 228469 1188
rect 228403 1123 228469 1124
rect 231347 1188 231413 1189
rect 231347 1124 231348 1188
rect 231412 1124 231413 1188
rect 231347 1123 231413 1124
rect 232083 1188 232149 1189
rect 232083 1124 232084 1188
rect 232148 1124 232149 1188
rect 232083 1123 232149 1124
rect 232819 1188 232885 1189
rect 232819 1124 232820 1188
rect 232884 1124 232885 1188
rect 232819 1123 232885 1124
rect 228406 0 228466 1123
rect 229139 372 229205 373
rect 229139 308 229140 372
rect 229204 308 229205 372
rect 229139 307 229205 308
rect 229875 372 229941 373
rect 229875 308 229876 372
rect 229940 308 229941 372
rect 229875 307 229941 308
rect 230611 372 230677 373
rect 230611 308 230612 372
rect 230676 308 230677 372
rect 230611 307 230677 308
rect 229142 0 229202 307
rect 229878 0 229938 307
rect 230614 0 230674 307
rect 231350 0 231410 1123
rect 232086 0 232146 1123
rect 232822 0 232882 1123
rect 235027 508 235093 509
rect 235027 444 235028 508
rect 235092 444 235093 508
rect 235027 443 235093 444
rect 233555 372 233621 373
rect 233555 308 233556 372
rect 233620 308 233621 372
rect 233555 307 233621 308
rect 234291 372 234357 373
rect 234291 308 234292 372
rect 234356 308 234357 372
rect 234291 307 234357 308
rect 233558 0 233618 307
rect 234294 0 234354 307
rect 235030 0 235090 443
rect 235766 0 235826 2755
rect 237533 2752 237853 3776
rect 258027 2820 258093 2821
rect 258027 2756 258028 2820
rect 258092 2756 258093 2820
rect 258027 2755 258093 2756
rect 237533 2688 237541 2752
rect 237605 2688 237621 2752
rect 237685 2688 237701 2752
rect 237765 2688 237781 2752
rect 237845 2688 237853 2752
rect 237533 1664 237853 2688
rect 237533 1600 237541 1664
rect 237605 1600 237621 1664
rect 237685 1600 237701 1664
rect 237765 1600 237781 1664
rect 237845 1600 237853 1664
rect 237235 1460 237301 1461
rect 237235 1396 237236 1460
rect 237300 1396 237301 1460
rect 237235 1395 237301 1396
rect 236499 1188 236565 1189
rect 236499 1124 236500 1188
rect 236564 1124 236565 1188
rect 236499 1123 236565 1124
rect 236502 0 236562 1123
rect 237238 0 237298 1395
rect 237533 1040 237853 1600
rect 242755 1460 242821 1461
rect 242755 1396 242756 1460
rect 242820 1396 242821 1460
rect 242755 1395 242821 1396
rect 244043 1460 244109 1461
rect 244043 1396 244044 1460
rect 244108 1396 244109 1460
rect 244043 1395 244109 1396
rect 247907 1460 247973 1461
rect 247907 1396 247908 1460
rect 247972 1396 247973 1460
rect 247907 1395 247973 1396
rect 249379 1460 249445 1461
rect 249379 1396 249380 1460
rect 249444 1396 249445 1460
rect 249379 1395 249445 1396
rect 250851 1460 250917 1461
rect 250851 1396 250852 1460
rect 250916 1396 250917 1460
rect 250851 1395 250917 1396
rect 241191 508 241257 509
rect 241191 444 241192 508
rect 241256 444 241257 508
rect 241191 443 241257 444
rect 241927 508 241993 509
rect 241927 444 241928 508
rect 241992 444 241993 508
rect 241927 443 241993 444
rect 239719 372 239785 373
rect 239719 308 239720 372
rect 239784 308 239785 372
rect 239719 307 239785 308
rect 240455 372 240521 373
rect 240455 308 240456 372
rect 240520 308 240521 372
rect 240455 307 240521 308
rect 239722 0 239782 307
rect 240458 0 240518 307
rect 241194 0 241254 443
rect 241930 0 241990 443
rect 242758 370 242818 1395
rect 243399 508 243465 509
rect 243399 444 243400 508
rect 243464 444 243465 508
rect 243399 443 243465 444
rect 242666 310 242818 370
rect 242666 0 242726 310
rect 243402 0 243462 443
rect 244046 370 244106 1395
rect 247171 1188 247237 1189
rect 247171 1124 247172 1188
rect 247236 1124 247237 1188
rect 247171 1123 247237 1124
rect 244871 508 244937 509
rect 244871 444 244872 508
rect 244936 444 244937 508
rect 244871 443 244937 444
rect 245607 508 245673 509
rect 245607 444 245608 508
rect 245672 444 245673 508
rect 245607 443 245673 444
rect 246343 508 246409 509
rect 246343 444 246344 508
rect 246408 444 246409 508
rect 246343 443 246409 444
rect 244046 310 244198 370
rect 244138 0 244198 310
rect 244874 0 244934 443
rect 245610 0 245670 443
rect 246346 0 246406 443
rect 247174 370 247234 1123
rect 247910 370 247970 1395
rect 248551 508 248617 509
rect 248551 444 248552 508
rect 248616 444 248617 508
rect 248551 443 248617 444
rect 247082 310 247234 370
rect 247818 310 247970 370
rect 247082 0 247142 310
rect 247818 0 247878 310
rect 248554 0 248614 443
rect 249382 370 249442 1395
rect 250023 644 250089 645
rect 250023 580 250024 644
rect 250088 580 250089 644
rect 250023 579 250089 580
rect 249290 310 249442 370
rect 249290 0 249350 310
rect 250026 0 250086 579
rect 250854 370 250914 1395
rect 251495 644 251561 645
rect 251495 580 251496 644
rect 251560 580 251561 644
rect 251495 579 251561 580
rect 252231 644 252297 645
rect 252231 580 252232 644
rect 252296 580 252297 644
rect 252231 579 252297 580
rect 252967 644 253033 645
rect 252967 580 252968 644
rect 253032 580 253033 644
rect 252967 579 253033 580
rect 253703 644 253769 645
rect 253703 580 253704 644
rect 253768 580 253769 644
rect 253703 579 253769 580
rect 255175 644 255241 645
rect 255175 580 255176 644
rect 255240 580 255241 644
rect 255175 579 255241 580
rect 255911 644 255977 645
rect 255911 580 255912 644
rect 255976 580 255977 644
rect 255911 579 255977 580
rect 256647 644 256713 645
rect 256647 580 256648 644
rect 256712 580 256713 644
rect 256647 579 256713 580
rect 257383 644 257449 645
rect 257383 580 257384 644
rect 257448 580 257449 644
rect 258030 642 258090 2755
rect 266494 2685 266554 8331
rect 266862 5677 266922 10238
rect 267411 7716 267477 7717
rect 267411 7652 267412 7716
rect 267476 7652 267477 7716
rect 267411 7651 267477 7652
rect 266859 5676 266925 5677
rect 266859 5612 266860 5676
rect 266924 5612 266925 5676
rect 266859 5611 266925 5612
rect 266491 2684 266557 2685
rect 266491 2620 266492 2684
rect 266556 2620 266557 2684
rect 266491 2619 266557 2620
rect 267414 1733 267474 7651
rect 267595 6764 267661 6765
rect 267595 6700 267596 6764
rect 267660 6700 267661 6764
rect 267595 6699 267661 6700
rect 267598 3773 267658 6699
rect 267782 5677 267842 10238
rect 268334 10238 268486 10298
rect 269162 10298 269222 10880
rect 269898 10298 269958 10880
rect 270634 10298 270694 10880
rect 271370 10298 271430 10880
rect 269162 10238 269314 10298
rect 267963 7580 268029 7581
rect 267963 7516 267964 7580
rect 268028 7516 268029 7580
rect 267963 7515 268029 7516
rect 267779 5676 267845 5677
rect 267779 5612 267780 5676
rect 267844 5612 267845 5676
rect 267779 5611 267845 5612
rect 267595 3772 267661 3773
rect 267595 3708 267596 3772
rect 267660 3708 267661 3772
rect 267595 3707 267661 3708
rect 267966 3229 268026 7515
rect 268147 6220 268213 6221
rect 268147 6156 268148 6220
rect 268212 6156 268213 6220
rect 268147 6155 268213 6156
rect 267963 3228 268029 3229
rect 267963 3164 267964 3228
rect 268028 3164 268029 3228
rect 267963 3163 268029 3164
rect 268150 2790 268210 6155
rect 268334 5677 268394 10238
rect 269254 5677 269314 10238
rect 269806 10238 269958 10298
rect 270542 10238 270694 10298
rect 271094 10238 271430 10298
rect 269806 5677 269866 10238
rect 270542 5677 270602 10238
rect 271094 5813 271154 10238
rect 271331 9824 271651 9840
rect 271331 9760 271339 9824
rect 271403 9760 271419 9824
rect 271483 9760 271499 9824
rect 271563 9760 271579 9824
rect 271643 9760 271651 9824
rect 271331 8736 271651 9760
rect 271331 8672 271339 8736
rect 271403 8672 271419 8736
rect 271483 8672 271499 8736
rect 271563 8672 271579 8736
rect 271643 8672 271651 8736
rect 271331 7648 271651 8672
rect 271331 7584 271339 7648
rect 271403 7584 271419 7648
rect 271483 7584 271499 7648
rect 271563 7584 271579 7648
rect 271643 7584 271651 7648
rect 271331 6560 271651 7584
rect 271331 6496 271339 6560
rect 271403 6496 271419 6560
rect 271483 6496 271499 6560
rect 271563 6496 271579 6560
rect 271643 6496 271651 6560
rect 271091 5812 271157 5813
rect 271091 5748 271092 5812
rect 271156 5748 271157 5812
rect 271091 5747 271157 5748
rect 268331 5676 268397 5677
rect 268331 5612 268332 5676
rect 268396 5612 268397 5676
rect 268331 5611 268397 5612
rect 269251 5676 269317 5677
rect 269251 5612 269252 5676
rect 269316 5612 269317 5676
rect 269251 5611 269317 5612
rect 269803 5676 269869 5677
rect 269803 5612 269804 5676
rect 269868 5612 269869 5676
rect 269803 5611 269869 5612
rect 270539 5676 270605 5677
rect 270539 5612 270540 5676
rect 270604 5612 270605 5676
rect 270539 5611 270605 5612
rect 271331 5472 271651 6496
rect 271331 5408 271339 5472
rect 271403 5408 271419 5472
rect 271483 5408 271499 5472
rect 271563 5408 271579 5472
rect 271643 5408 271651 5472
rect 271331 4384 271651 5408
rect 271331 4320 271339 4384
rect 271403 4320 271419 4384
rect 271483 4320 271499 4384
rect 271563 4320 271579 4384
rect 271643 4320 271651 4384
rect 271331 3296 271651 4320
rect 271331 3232 271339 3296
rect 271403 3232 271419 3296
rect 271483 3232 271499 3296
rect 271563 3232 271579 3296
rect 271643 3232 271651 3296
rect 267966 2730 268210 2790
rect 270539 2820 270605 2821
rect 270539 2756 270540 2820
rect 270604 2756 270605 2820
rect 270539 2755 270605 2756
rect 267966 2549 268026 2730
rect 267963 2548 268029 2549
rect 267963 2484 267964 2548
rect 268028 2484 268029 2548
rect 267963 2483 268029 2484
rect 267411 1732 267477 1733
rect 267411 1668 267412 1732
rect 267476 1668 267477 1732
rect 267411 1667 267477 1668
rect 264835 1460 264901 1461
rect 264835 1396 264836 1460
rect 264900 1396 264901 1460
rect 264835 1395 264901 1396
rect 258855 644 258921 645
rect 258030 582 258182 642
rect 257383 579 257449 580
rect 250762 310 250914 370
rect 250762 0 250822 310
rect 251498 0 251558 579
rect 252234 0 252294 579
rect 252970 0 253030 579
rect 253706 0 253766 579
rect 254439 372 254505 373
rect 254439 308 254440 372
rect 254504 308 254505 372
rect 254439 307 254505 308
rect 254442 0 254502 307
rect 255178 0 255238 579
rect 255914 0 255974 579
rect 256650 0 256710 579
rect 257386 0 257446 579
rect 258122 0 258182 582
rect 258855 580 258856 644
rect 258920 580 258921 644
rect 258855 579 258921 580
rect 259591 644 259657 645
rect 259591 580 259592 644
rect 259656 580 259657 644
rect 259591 579 259657 580
rect 260327 644 260393 645
rect 260327 580 260328 644
rect 260392 580 260393 644
rect 260327 579 260393 580
rect 261063 644 261129 645
rect 261063 580 261064 644
rect 261128 580 261129 644
rect 261063 579 261129 580
rect 262535 644 262601 645
rect 262535 580 262536 644
rect 262600 580 262601 644
rect 262535 579 262601 580
rect 263271 644 263337 645
rect 263271 580 263272 644
rect 263336 580 263337 644
rect 263271 579 263337 580
rect 264007 644 264073 645
rect 264007 580 264008 644
rect 264072 580 264073 644
rect 264007 579 264073 580
rect 258858 0 258918 579
rect 259594 0 259654 579
rect 260330 0 260390 579
rect 261066 0 261126 579
rect 261799 508 261865 509
rect 261799 444 261800 508
rect 261864 444 261865 508
rect 261799 443 261865 444
rect 261802 0 261862 443
rect 262538 0 262598 579
rect 263274 0 263334 579
rect 264010 0 264070 579
rect 264838 370 264898 1395
rect 265479 644 265545 645
rect 265479 580 265480 644
rect 265544 580 265545 644
rect 265479 579 265545 580
rect 266215 644 266281 645
rect 266215 580 266216 644
rect 266280 580 266281 644
rect 266215 579 266281 580
rect 266951 644 267017 645
rect 266951 580 266952 644
rect 267016 580 267017 644
rect 266951 579 267017 580
rect 267687 644 267753 645
rect 267687 580 267688 644
rect 267752 580 267753 644
rect 267687 579 267753 580
rect 268423 644 268489 645
rect 268423 580 268424 644
rect 268488 580 268489 644
rect 268423 579 268489 580
rect 269895 644 269961 645
rect 269895 580 269896 644
rect 269960 580 269961 644
rect 269895 579 269961 580
rect 264746 310 264898 370
rect 264746 0 264806 310
rect 265482 0 265542 579
rect 266218 0 266278 579
rect 266954 0 267014 579
rect 267690 0 267750 579
rect 268426 0 268486 579
rect 269159 508 269225 509
rect 269159 444 269160 508
rect 269224 444 269225 508
rect 269159 443 269225 444
rect 269162 0 269222 443
rect 269898 0 269958 579
rect 270542 370 270602 2755
rect 271331 2208 271651 3232
rect 271331 2144 271339 2208
rect 271403 2144 271419 2208
rect 271483 2144 271499 2208
rect 271563 2144 271579 2208
rect 271643 2144 271651 2208
rect 271331 1120 271651 2144
rect 271331 1056 271339 1120
rect 271403 1056 271419 1120
rect 271483 1056 271499 1120
rect 271563 1056 271579 1120
rect 271643 1056 271651 1120
rect 271331 1040 271651 1056
rect 271367 372 271433 373
rect 270542 310 270694 370
rect 270634 0 270694 310
rect 271367 308 271368 372
rect 271432 308 271433 372
rect 271367 307 271433 308
rect 271370 0 271430 307
use sky130_fd_sc_hd__nor3_4  _048_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 181700 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3b_4  _049_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 181608 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__nor3b_2  _050_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 181700 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_1  _051_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 228068 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _052_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 229080 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _053_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 267812 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _054_
timestamp 1676037725
transform 1 0 268088 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _055_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 267444 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _056_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 270756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _057_
timestamp 1676037725
transform 1 0 270572 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _058_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 267168 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _059_
timestamp 1676037725
transform 1 0 269100 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _060_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 268180 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _061_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 270112 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _062_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 264224 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_2  _063_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 80132 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _064_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40112 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  _065_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 125028 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _066_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 81236 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _067_
timestamp 1676037725
transform 1 0 129812 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _068_
timestamp 1676037725
transform 1 0 79028 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1676037725
transform 1 0 42596 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _070_
timestamp 1676037725
transform 1 0 78936 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _071_
timestamp 1676037725
transform 1 0 66976 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _072_
timestamp 1676037725
transform 1 0 79028 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1676037725
transform 1 0 67344 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _074_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 99360 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _075_
timestamp 1676037725
transform 1 0 99360 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _076_
timestamp 1676037725
transform 1 0 100648 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _077_
timestamp 1676037725
transform 1 0 99728 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1676037725
transform 1 0 100004 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _079_
timestamp 1676037725
transform 1 0 120704 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _080_
timestamp 1676037725
transform 1 0 122452 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _081_
timestamp 1676037725
transform 1 0 119876 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1676037725
transform 1 0 121164 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _083_
timestamp 1676037725
transform 1 0 162472 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _084_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 162932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _085_
timestamp 1676037725
transform 1 0 180596 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _086_
timestamp 1676037725
transform 1 0 169188 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1676037725
transform 1 0 169096 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _088_
timestamp 1676037725
transform 1 0 188784 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _089_
timestamp 1676037725
transform 1 0 189888 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _090_
timestamp 1676037725
transform 1 0 188968 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1676037725
transform 1 0 189980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _092_
timestamp 1676037725
transform 1 0 230644 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1676037725
transform 1 0 230644 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _094_
timestamp 1676037725
transform 1 0 231472 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _095_
timestamp 1676037725
transform 1 0 229540 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1676037725
transform 1 0 229540 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _097_
timestamp 1676037725
transform 1 0 230920 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _098_
timestamp 1676037725
transform 1 0 235520 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _099_
timestamp 1676037725
transform 1 0 230644 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _100_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 232300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _137_
timestamp 1676037725
transform 1 0 244996 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _138_
timestamp 1676037725
transform 1 0 243800 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _139_
timestamp 1676037725
transform 1 0 242144 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _140_
timestamp 1676037725
transform 1 0 240304 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _141_
timestamp 1676037725
transform 1 0 260360 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _142_
timestamp 1676037725
transform 1 0 259808 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _143_
timestamp 1676037725
transform 1 0 260084 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _144_
timestamp 1676037725
transform 1 0 257968 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _145_
timestamp 1676037725
transform 1 0 259532 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _146_
timestamp 1676037725
transform 1 0 251988 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _147_
timestamp 1676037725
transform 1 0 260820 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _148_
timestamp 1676037725
transform 1 0 258888 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _149_
timestamp 1676037725
transform 1 0 259716 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _150_ openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 222916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _151_
timestamp 1676037725
transform 1 0 218868 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _152_
timestamp 1676037725
transform 1 0 216384 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _153_
timestamp 1676037725
transform 1 0 217764 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _154_
timestamp 1676037725
transform 1 0 218684 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _155_
timestamp 1676037725
transform 1 0 219788 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _156_
timestamp 1676037725
transform 1 0 220708 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _157_
timestamp 1676037725
transform 1 0 227884 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _158_
timestamp 1676037725
transform 1 0 222916 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _159_
timestamp 1676037725
transform 1 0 223836 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _160_
timestamp 1676037725
transform 1 0 223744 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _161_
timestamp 1676037725
transform 1 0 33120 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _162_
timestamp 1676037725
transform 1 0 32384 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _163_
timestamp 1676037725
transform 1 0 67344 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _164_
timestamp 1676037725
transform 1 0 66700 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _165_
timestamp 1676037725
transform 1 0 101108 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _166_
timestamp 1676037725
transform 1 0 100464 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _167_
timestamp 1676037725
transform 1 0 135332 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _168_
timestamp 1676037725
transform 1 0 134688 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _169_
timestamp 1676037725
transform 1 0 168820 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _170_
timestamp 1676037725
transform 1 0 170292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _171_
timestamp 1676037725
transform 1 0 203136 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _172_
timestamp 1676037725
transform 1 0 203872 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _173_
timestamp 1676037725
transform 1 0 237360 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _174_
timestamp 1676037725
transform 1 0 237360 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _175_
timestamp 1676037725
transform 1 0 270572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _176_
timestamp 1676037725
transform 1 0 269836 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _177_
timestamp 1676037725
transform 1 0 32292 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _178_
timestamp 1676037725
transform 1 0 31372 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _179_
timestamp 1676037725
transform 1 0 30544 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _180_
timestamp 1676037725
transform 1 0 29716 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _181_
timestamp 1676037725
transform 1 0 28888 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _182_
timestamp 1676037725
transform 1 0 28520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _183_
timestamp 1676037725
transform 1 0 27232 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _184_
timestamp 1676037725
transform 1 0 26496 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _185_
timestamp 1676037725
transform 1 0 25760 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _186_
timestamp 1676037725
transform 1 0 27968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _187_
timestamp 1676037725
transform 1 0 25760 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _188_
timestamp 1676037725
transform 1 0 23736 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _189_
timestamp 1676037725
transform 1 0 24288 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _190_
timestamp 1676037725
transform 1 0 23736 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _191_
timestamp 1676037725
transform 1 0 25116 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _192_
timestamp 1676037725
transform 1 0 25760 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _193_
timestamp 1676037725
transform 1 0 26128 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _194_
timestamp 1676037725
transform 1 0 27140 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _195_
timestamp 1676037725
transform 1 0 33396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _196_
timestamp 1676037725
transform 1 0 31096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _197_
timestamp 1676037725
transform 1 0 30268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _198_
timestamp 1676037725
transform 1 0 29440 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _199_
timestamp 1676037725
transform 1 0 28612 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _200_
timestamp 1676037725
transform 1 0 28152 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _201_
timestamp 1676037725
transform 1 0 28888 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _202_
timestamp 1676037725
transform 1 0 26496 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _203_
timestamp 1676037725
transform 1 0 29716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _204_
timestamp 1676037725
transform 1 0 27784 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _205_
timestamp 1676037725
transform 1 0 23276 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _206_
timestamp 1676037725
transform 1 0 25576 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _207_
timestamp 1676037725
transform 1 0 24472 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _208_
timestamp 1676037725
transform 1 0 25024 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _209_
timestamp 1676037725
transform 1 0 25024 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _210_
timestamp 1676037725
transform 1 0 25668 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _211_
timestamp 1676037725
transform 1 0 25944 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _212_
timestamp 1676037725
transform 1 0 27140 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _213_
timestamp 1676037725
transform 1 0 65964 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _214_
timestamp 1676037725
transform 1 0 65780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _215_
timestamp 1676037725
transform 1 0 64308 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _216_
timestamp 1676037725
transform 1 0 63572 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _217_
timestamp 1676037725
transform 1 0 62744 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _218_
timestamp 1676037725
transform 1 0 62100 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _219_
timestamp 1676037725
transform 1 0 61364 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _220_
timestamp 1676037725
transform 1 0 60628 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _221_
timestamp 1676037725
transform 1 0 60628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _222_
timestamp 1676037725
transform 1 0 59156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _223_
timestamp 1676037725
transform 1 0 58420 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _224_
timestamp 1676037725
transform 1 0 57592 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _225_
timestamp 1676037725
transform 1 0 56856 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _226_
timestamp 1676037725
transform 1 0 56028 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _227_
timestamp 1676037725
transform 1 0 55476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _228_
timestamp 1676037725
transform 1 0 54648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _229_
timestamp 1676037725
transform 1 0 52900 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _230_
timestamp 1676037725
transform 1 0 53176 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _231_
timestamp 1676037725
transform 1 0 65964 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _232_
timestamp 1676037725
transform 1 0 65228 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _233_
timestamp 1676037725
transform 1 0 64400 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _234_
timestamp 1676037725
transform 1 0 63572 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _235_
timestamp 1676037725
transform 1 0 63204 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _236_
timestamp 1676037725
transform 1 0 62100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _237_
timestamp 1676037725
transform 1 0 61364 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _238_
timestamp 1676037725
transform 1 0 60628 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _239_
timestamp 1676037725
transform 1 0 59800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _240_
timestamp 1676037725
transform 1 0 59064 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _241_
timestamp 1676037725
transform 1 0 58420 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _242_
timestamp 1676037725
transform 1 0 58052 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _243_
timestamp 1676037725
transform 1 0 56856 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _244_
timestamp 1676037725
transform 1 0 56028 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _245_
timestamp 1676037725
transform 1 0 55292 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _246_
timestamp 1676037725
transform 1 0 54556 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _247_
timestamp 1676037725
transform 1 0 54464 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _248_
timestamp 1676037725
transform 1 0 52992 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _249_
timestamp 1676037725
transform 1 0 100740 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _250_
timestamp 1676037725
transform 1 0 101844 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _251_
timestamp 1676037725
transform 1 0 97612 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _252_
timestamp 1676037725
transform 1 0 96876 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _253_
timestamp 1676037725
transform 1 0 95864 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _254_
timestamp 1676037725
transform 1 0 95864 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _255_
timestamp 1676037725
transform 1 0 95128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _256_
timestamp 1676037725
transform 1 0 94392 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _257_
timestamp 1676037725
transform 1 0 93656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _258_
timestamp 1676037725
transform 1 0 93288 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _259_
timestamp 1676037725
transform 1 0 92828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _260_
timestamp 1676037725
transform 1 0 92000 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _261_
timestamp 1676037725
transform 1 0 91540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _262_
timestamp 1676037725
transform 1 0 90436 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _263_
timestamp 1676037725
transform 1 0 90620 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _264_
timestamp 1676037725
transform 1 0 89148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _265_
timestamp 1676037725
transform 1 0 87400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _266_
timestamp 1676037725
transform 1 0 87952 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _267_
timestamp 1676037725
transform 1 0 100648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _268_
timestamp 1676037725
transform 1 0 99360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _269_
timestamp 1676037725
transform 1 0 98440 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _270_
timestamp 1676037725
transform 1 0 97980 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _271_
timestamp 1676037725
transform 1 0 97244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _272_
timestamp 1676037725
transform 1 0 96692 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _273_
timestamp 1676037725
transform 1 0 95772 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _274_
timestamp 1676037725
transform 1 0 95128 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _275_
timestamp 1676037725
transform 1 0 94392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _276_
timestamp 1676037725
transform 1 0 93288 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _277_
timestamp 1676037725
transform 1 0 93104 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _278_
timestamp 1676037725
transform 1 0 92368 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _279_
timestamp 1676037725
transform 1 0 91632 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _280_
timestamp 1676037725
transform 1 0 90896 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _281_
timestamp 1676037725
transform 1 0 90160 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _282_
timestamp 1676037725
transform 1 0 89516 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _283_
timestamp 1676037725
transform 1 0 88228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _284_
timestamp 1676037725
transform 1 0 88780 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _285_
timestamp 1676037725
transform 1 0 134228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _286_
timestamp 1676037725
transform 1 0 133492 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _287_
timestamp 1676037725
transform 1 0 132756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _288_
timestamp 1676037725
transform 1 0 131928 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _289_
timestamp 1676037725
transform 1 0 131376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _290_
timestamp 1676037725
transform 1 0 130640 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _291_
timestamp 1676037725
transform 1 0 129812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _292_
timestamp 1676037725
transform 1 0 129076 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _293_
timestamp 1676037725
transform 1 0 128340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _294_
timestamp 1676037725
transform 1 0 127604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _295_
timestamp 1676037725
transform 1 0 126776 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _296_
timestamp 1676037725
transform 1 0 126132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _297_
timestamp 1676037725
transform 1 0 125396 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _298_
timestamp 1676037725
transform 1 0 124568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _299_
timestamp 1676037725
transform 1 0 123740 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _300_
timestamp 1676037725
transform 1 0 122912 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _301_
timestamp 1676037725
transform 1 0 122452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _302_
timestamp 1676037725
transform 1 0 121624 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _303_
timestamp 1676037725
transform 1 0 134044 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _304_
timestamp 1676037725
transform 1 0 133308 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _305_
timestamp 1676037725
transform 1 0 132848 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _306_
timestamp 1676037725
transform 1 0 132112 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _307_
timestamp 1676037725
transform 1 0 131284 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _308_
timestamp 1676037725
transform 1 0 131376 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _309_
timestamp 1676037725
transform 1 0 129352 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _310_
timestamp 1676037725
transform 1 0 128616 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _311_
timestamp 1676037725
transform 1 0 127604 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _312_
timestamp 1676037725
transform 1 0 127696 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _313_
timestamp 1676037725
transform 1 0 126868 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _314_
timestamp 1676037725
transform 1 0 126132 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _315_
timestamp 1676037725
transform 1 0 125396 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _316_
timestamp 1676037725
transform 1 0 125028 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _317_
timestamp 1676037725
transform 1 0 123740 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _318_
timestamp 1676037725
transform 1 0 123004 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _319_
timestamp 1676037725
transform 1 0 122452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _320_
timestamp 1676037725
transform 1 0 120796 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _321_
timestamp 1676037725
transform 1 0 168728 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _322_
timestamp 1676037725
transform 1 0 167808 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _323_
timestamp 1676037725
transform 1 0 166612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _324_
timestamp 1676037725
transform 1 0 165876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _325_
timestamp 1676037725
transform 1 0 165140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _326_
timestamp 1676037725
transform 1 0 164496 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _327_
timestamp 1676037725
transform 1 0 164404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _328_
timestamp 1676037725
transform 1 0 163668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _329_
timestamp 1676037725
transform 1 0 162288 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _330_
timestamp 1676037725
transform 1 0 161552 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _331_
timestamp 1676037725
transform 1 0 161092 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _332_
timestamp 1676037725
transform 1 0 160724 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _333_
timestamp 1676037725
transform 1 0 160356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _334_
timestamp 1676037725
transform 1 0 160172 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _335_
timestamp 1676037725
transform 1 0 155112 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _336_
timestamp 1676037725
transform 1 0 157688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _337_
timestamp 1676037725
transform 1 0 157320 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _338_
timestamp 1676037725
transform 1 0 155940 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _339_
timestamp 1676037725
transform 1 0 168820 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _340_
timestamp 1676037725
transform 1 0 167624 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _341_
timestamp 1676037725
transform 1 0 166888 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _342_
timestamp 1676037725
transform 1 0 166152 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _343_
timestamp 1676037725
transform 1 0 165324 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _344_
timestamp 1676037725
transform 1 0 164588 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _345_
timestamp 1676037725
transform 1 0 165416 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _346_
timestamp 1676037725
transform 1 0 163852 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _347_
timestamp 1676037725
transform 1 0 162380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _348_
timestamp 1676037725
transform 1 0 162196 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _349_
timestamp 1676037725
transform 1 0 161092 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _350_
timestamp 1676037725
transform 1 0 160080 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _351_
timestamp 1676037725
transform 1 0 159988 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _352_
timestamp 1676037725
transform 1 0 159252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _353_
timestamp 1676037725
transform 1 0 158516 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _354_
timestamp 1676037725
transform 1 0 157412 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _355_
timestamp 1676037725
transform 1 0 156676 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _356_
timestamp 1676037725
transform 1 0 155940 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _357_
timestamp 1676037725
transform 1 0 202768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _358_
timestamp 1676037725
transform 1 0 203136 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _359_
timestamp 1676037725
transform 1 0 201204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _360_
timestamp 1676037725
transform 1 0 200468 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _361_
timestamp 1676037725
transform 1 0 199732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _362_
timestamp 1676037725
transform 1 0 199732 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _363_
timestamp 1676037725
transform 1 0 198352 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _364_
timestamp 1676037725
transform 1 0 197892 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _365_
timestamp 1676037725
transform 1 0 197156 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _366_
timestamp 1676037725
transform 1 0 196236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _367_
timestamp 1676037725
transform 1 0 195592 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _368_
timestamp 1676037725
transform 1 0 194856 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _369_
timestamp 1676037725
transform 1 0 194580 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _370_
timestamp 1676037725
transform 1 0 193292 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _371_
timestamp 1676037725
transform 1 0 192464 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _372_
timestamp 1676037725
transform 1 0 191820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _373_
timestamp 1676037725
transform 1 0 191084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _374_
timestamp 1676037725
transform 1 0 190348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _375_
timestamp 1676037725
transform 1 0 203044 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _376_
timestamp 1676037725
transform 1 0 202308 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _377_
timestamp 1676037725
transform 1 0 201388 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _378_
timestamp 1676037725
transform 1 0 200652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _379_
timestamp 1676037725
transform 1 0 199824 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _380_
timestamp 1676037725
transform 1 0 199272 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _381_
timestamp 1676037725
transform 1 0 198628 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _382_
timestamp 1676037725
transform 1 0 197892 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _383_
timestamp 1676037725
transform 1 0 197156 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _384_
timestamp 1676037725
transform 1 0 196144 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _385_
timestamp 1676037725
transform 1 0 195408 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _386_
timestamp 1676037725
transform 1 0 194672 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _387_
timestamp 1676037725
transform 1 0 194028 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _388_
timestamp 1676037725
transform 1 0 193200 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _389_
timestamp 1676037725
transform 1 0 192372 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _390_
timestamp 1676037725
transform 1 0 192004 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _391_
timestamp 1676037725
transform 1 0 191084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _392_
timestamp 1676037725
transform 1 0 190348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _393_
timestamp 1676037725
transform 1 0 236532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _394_
timestamp 1676037725
transform 1 0 235796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _395_
timestamp 1676037725
transform 1 0 234692 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _396_
timestamp 1676037725
transform 1 0 233956 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _397_
timestamp 1676037725
transform 1 0 233220 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _398_
timestamp 1676037725
transform 1 0 232576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _399_
timestamp 1676037725
transform 1 0 231840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _400_
timestamp 1676037725
transform 1 0 231104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _401_
timestamp 1676037725
transform 1 0 230644 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _402_
timestamp 1676037725
transform 1 0 229632 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _403_
timestamp 1676037725
transform 1 0 228896 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _404_
timestamp 1676037725
transform 1 0 228804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _405_
timestamp 1676037725
transform 1 0 228068 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _406_
timestamp 1676037725
transform 1 0 227056 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _407_
timestamp 1676037725
transform 1 0 226964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _408_
timestamp 1676037725
transform 1 0 226228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _409_
timestamp 1676037725
transform 1 0 225676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _410_
timestamp 1676037725
transform 1 0 225308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _411_
timestamp 1676037725
transform 1 0 236440 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _412_
timestamp 1676037725
transform 1 0 236624 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _413_
timestamp 1676037725
transform 1 0 234876 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _414_
timestamp 1676037725
transform 1 0 234140 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _415_
timestamp 1676037725
transform 1 0 233312 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _416_
timestamp 1676037725
transform 1 0 233220 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _417_
timestamp 1676037725
transform 1 0 231748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _418_
timestamp 1676037725
transform 1 0 231380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _419_
timestamp 1676037725
transform 1 0 230644 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _420_
timestamp 1676037725
transform 1 0 229632 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _421_
timestamp 1676037725
transform 1 0 228896 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _422_
timestamp 1676037725
transform 1 0 228160 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _423_
timestamp 1676037725
transform 1 0 228068 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _424_
timestamp 1676037725
transform 1 0 226504 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _425_
timestamp 1676037725
transform 1 0 225768 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _426_
timestamp 1676037725
transform 1 0 225492 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _427_
timestamp 1676037725
transform 1 0 225032 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _428_
timestamp 1676037725
transform 1 0 223192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _429_
timestamp 1676037725
transform 1 0 269836 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _430_
timestamp 1676037725
transform 1 0 270112 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _431_
timestamp 1676037725
transform 1 0 269836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _432_
timestamp 1676037725
transform 1 0 268180 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _433_
timestamp 1676037725
transform 1 0 267444 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _434_
timestamp 1676037725
transform 1 0 266708 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _435_
timestamp 1676037725
transform 1 0 265880 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _436_
timestamp 1676037725
transform 1 0 265144 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _437_
timestamp 1676037725
transform 1 0 264776 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _438_
timestamp 1676037725
transform 1 0 264132 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _439_
timestamp 1676037725
transform 1 0 263028 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _440_
timestamp 1676037725
transform 1 0 262292 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _441_
timestamp 1676037725
transform 1 0 261556 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _442_
timestamp 1676037725
transform 1 0 261556 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _443_
timestamp 1676037725
transform 1 0 260268 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _444_
timestamp 1676037725
transform 1 0 259716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _445_
timestamp 1676037725
transform 1 0 258980 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _446_
timestamp 1676037725
transform 1 0 257600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _447_
timestamp 1676037725
transform 1 0 270020 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _448_
timestamp 1676037725
transform 1 0 269100 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _449_
timestamp 1676037725
transform 1 0 269284 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _450_
timestamp 1676037725
transform 1 0 267628 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _451_
timestamp 1676037725
transform 1 0 267536 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _452_
timestamp 1676037725
transform 1 0 266708 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _453_
timestamp 1676037725
transform 1 0 263304 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _454_
timestamp 1676037725
transform 1 0 265512 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _455_
timestamp 1676037725
transform 1 0 264040 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _456_
timestamp 1676037725
transform 1 0 264132 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _457_
timestamp 1676037725
transform 1 0 263028 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _458_
timestamp 1676037725
transform 1 0 262292 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _459_
timestamp 1676037725
transform 1 0 261556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _460_
timestamp 1676037725
transform 1 0 262200 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _461_
timestamp 1676037725
transform 1 0 260268 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _462_
timestamp 1676037725
transform 1 0 259808 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _463_
timestamp 1676037725
transform 1 0 258796 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _464_
timestamp 1676037725
transform 1 0 258060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40848 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 43056 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 84364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 86848 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 124568 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 121808 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 161092 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 163116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 230184 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 227424 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 243524 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1676037725
transform 1 0 244812 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1676037725
transform 1 0 94116 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1676037725
transform 1 0 94484 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1676037725
transform 1 0 94852 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1676037725
transform 1 0 108652 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1676037725
transform 1 0 111136 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1676037725
transform 1 0 108284 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1676037725
transform 1 0 150328 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1676037725
transform 1 0 147568 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1676037725
transform 1 0 150696 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1676037725
transform 1 0 212428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1676037725
transform 1 0 215188 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1676037725
transform 1 0 212060 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1676037725
transform 1 0 259624 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1676037725
transform 1 0 258704 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1676037725
transform 1 0 256404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1676037725
transform 1 0 259072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1676037725
transform 1 0 88964 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1676037725
transform 1 0 88964 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1676037725
transform 1 0 103960 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1676037725
transform 1 0 104420 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1676037725
transform 1 0 141404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1676037725
transform 1 0 143888 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1676037725
transform 1 0 209300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1676037725
transform 1 0 210036 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1676037725
transform 1 0 218684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1676037725
transform 1 0 219512 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1676037725
transform 1 0 81052 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1676037725
transform 1 0 121348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1676037725
transform 1 0 160448 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_42
timestamp 1676037725
transform 1 0 226136 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_43
timestamp 1676037725
transform 1 0 242236 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_44
timestamp 1676037725
transform 1 0 83904 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_45
timestamp 1676037725
transform 1 0 83168 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_46
timestamp 1676037725
transform 1 0 99084 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_47
timestamp 1676037725
transform 1 0 98716 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_48
timestamp 1676037725
transform 1 0 142600 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_49
timestamp 1676037725
transform 1 0 139840 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_50
timestamp 1676037725
transform 1 0 207000 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_51
timestamp 1676037725
transform 1 0 204240 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_52
timestamp 1676037725
transform 1 0 220432 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_53
timestamp 1676037725
transform 1 0 222824 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_54
timestamp 1676037725
transform 1 0 83168 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_55
timestamp 1676037725
transform 1 0 85652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_56
timestamp 1676037725
transform 1 0 101476 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_57
timestamp 1676037725
transform 1 0 98624 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_58
timestamp 1676037725
transform 1 0 138552 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_59
timestamp 1676037725
transform 1 0 141036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_60
timestamp 1676037725
transform 1 0 204240 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_61
timestamp 1676037725
transform 1 0 203872 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_62
timestamp 1676037725
transform 1 0 224112 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_63
timestamp 1676037725
transform 1 0 224480 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_64
timestamp 1676037725
transform 1 0 85928 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_65
timestamp 1676037725
transform 1 0 98992 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_66
timestamp 1676037725
transform 1 0 138552 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_67
timestamp 1676037725
transform 1 0 203780 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_68
timestamp 1676037725
transform 1 0 224848 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_69
timestamp 1676037725
transform 1 0 81328 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_70
timestamp 1676037725
transform 1 0 80592 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_71
timestamp 1676037725
transform 1 0 80224 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_72
timestamp 1676037725
transform 1 0 117116 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_73
timestamp 1676037725
transform 1 0 119876 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_74
timestamp 1676037725
transform 1 0 116748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_75
timestamp 1676037725
transform 1 0 160356 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_76
timestamp 1676037725
transform 1 0 161460 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_77
timestamp 1676037725
transform 1 0 161552 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_78
timestamp 1676037725
transform 1 0 223284 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_79
timestamp 1676037725
transform 1 0 225768 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_80
timestamp 1676037725
transform 1 0 222916 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_81
timestamp 1676037725
transform 1 0 251528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_82
timestamp 1676037725
transform 1 0 252908 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_83
timestamp 1676037725
transform 1 0 251160 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_84
timestamp 1676037725
transform 1 0 250792 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_85
timestamp 1676037725
transform 1 0 83812 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_86
timestamp 1676037725
transform 1 0 84180 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_87
timestamp 1676037725
transform 1 0 84548 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_88
timestamp 1676037725
transform 1 0 116104 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_89
timestamp 1676037725
transform 1 0 118588 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_90
timestamp 1676037725
transform 1 0 115736 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_91
timestamp 1676037725
transform 1 0 155296 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_92
timestamp 1676037725
transform 1 0 160080 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_93
timestamp 1676037725
transform 1 0 160448 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_94
timestamp 1676037725
transform 1 0 225032 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_95
timestamp 1676037725
transform 1 0 222272 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_96
timestamp 1676037725
transform 1 0 224664 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_97
timestamp 1676037725
transform 1 0 254840 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_98
timestamp 1676037725
transform 1 0 255208 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_99
timestamp 1676037725
transform 1 0 256036 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_100
timestamp 1676037725
transform 1 0 86388 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_101
timestamp 1676037725
transform 1 0 86756 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_102
timestamp 1676037725
transform 1 0 87124 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_103
timestamp 1676037725
transform 1 0 87492 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_104
timestamp 1676037725
transform 1 0 114724 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_105
timestamp 1676037725
transform 1 0 114080 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_106
timestamp 1676037725
transform 1 0 119232 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_107
timestamp 1676037725
transform 1 0 118956 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_108
timestamp 1676037725
transform 1 0 157780 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_109
timestamp 1676037725
transform 1 0 158516 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_110
timestamp 1676037725
transform 1 0 158884 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_111
timestamp 1676037725
transform 1 0 159252 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_112
timestamp 1676037725
transform 1 0 221444 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_113
timestamp 1676037725
transform 1 0 223928 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_114
timestamp 1676037725
transform 1 0 221076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_115
timestamp 1676037725
transform 1 0 224296 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_116
timestamp 1676037725
transform 1 0 253920 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_117
timestamp 1676037725
transform 1 0 255300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_118
timestamp 1676037725
transform 1 0 253552 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_119
timestamp 1676037725
transform 1 0 255668 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_120
timestamp 1676037725
transform 1 0 89976 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_121
timestamp 1676037725
transform 1 0 90344 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_122
timestamp 1676037725
transform 1 0 90712 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_123
timestamp 1676037725
transform 1 0 113712 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_124
timestamp 1676037725
transform 1 0 116196 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_125
timestamp 1676037725
transform 1 0 113344 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_126
timestamp 1676037725
transform 1 0 152720 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_127
timestamp 1676037725
transform 1 0 152352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_128
timestamp 1676037725
transform 1 0 151984 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_129
timestamp 1676037725
transform 1 0 222732 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_130
timestamp 1676037725
transform 1 0 223100 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_131
timestamp 1676037725
transform 1 0 219696 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_132
timestamp 1676037725
transform 1 0 260544 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_133
timestamp 1676037725
transform 1 0 258520 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_134
timestamp 1676037725
transform 1 0 259072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_135
timestamp 1676037725
transform 1 0 89056 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_136
timestamp 1676037725
transform 1 0 88320 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_137
timestamp 1676037725
transform 1 0 112792 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_138
timestamp 1676037725
transform 1 0 115276 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_139
timestamp 1676037725
transform 1 0 158056 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_140
timestamp 1676037725
transform 1 0 158056 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_141
timestamp 1676037725
transform 1 0 218868 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_142
timestamp 1676037725
transform 1 0 221352 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_143
timestamp 1676037725
transform 1 0 256680 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_144
timestamp 1676037725
transform 1 0 259808 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_145
timestamp 1676037725
transform 1 0 162104 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_146
timestamp 1676037725
transform 1 0 267720 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_147
timestamp 1676037725
transform 1 0 163852 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_148
timestamp 1676037725
transform 1 0 266708 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_149
timestamp 1676037725
transform 1 0 163208 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_150
timestamp 1676037725
transform 1 0 263488 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_151
timestamp 1676037725
transform 1 0 164680 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_152
timestamp 1676037725
transform 1 0 264776 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_153
timestamp 1676037725
transform 1 0 161828 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_154
timestamp 1676037725
transform 1 0 263120 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_155
timestamp 1676037725
transform 1 0 161736 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_156
timestamp 1676037725
transform 1 0 262752 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_157
timestamp 1676037725
transform 1 0 81880 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_158
timestamp 1676037725
transform 1 0 100280 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_159
timestamp 1676037725
transform 1 0 180228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_160
timestamp 1676037725
transform 1 0 239016 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_161
timestamp 1676037725
transform 1 0 236624 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_162
timestamp 1676037725
transform 1 0 111688 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_163
timestamp 1676037725
transform 1 0 107732 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_164
timestamp 1676037725
transform 1 0 104144 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_165
timestamp 1676037725
transform 1 0 42688 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_166
timestamp 1676037725
transform 1 0 105708 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_167
timestamp 1676037725
transform 1 0 98992 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_168
timestamp 1676037725
transform 1 0 96508 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_169
timestamp 1676037725
transform 1 0 119876 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_170
timestamp 1676037725
transform 1 0 111412 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_171
timestamp 1676037725
transform 1 0 109388 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_172
timestamp 1676037725
transform 1 0 108928 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_173
timestamp 1676037725
transform 1 0 44436 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_174
timestamp 1676037725
transform 1 0 110216 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_175
timestamp 1676037725
transform 1 0 106076 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_176
timestamp 1676037725
transform 1 0 103776 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_177
timestamp 1676037725
transform 1 0 108192 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_178
timestamp 1676037725
transform 1 0 45172 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_179
timestamp 1676037725
transform 1 0 98624 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_180
timestamp 1676037725
transform 1 0 40388 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_181
timestamp 1676037725
transform 1 0 161276 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_182
timestamp 1676037725
transform 1 0 155296 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_183
timestamp 1676037725
transform 1 0 140300 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_184
timestamp 1676037725
transform 1 0 155296 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_185
timestamp 1676037725
transform 1 0 150144 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_186
timestamp 1676037725
transform 1 0 147752 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_187
timestamp 1676037725
transform 1 0 227608 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_188
timestamp 1676037725
transform 1 0 227608 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_189
timestamp 1676037725
transform 1 0 217304 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_190
timestamp 1676037725
transform 1 0 42596 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_191
timestamp 1676037725
transform 1 0 223928 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_192
timestamp 1676037725
transform 1 0 224848 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_193
timestamp 1676037725
transform 1 0 225032 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_194
timestamp 1676037725
transform 1 0 222272 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_195
timestamp 1676037725
transform 1 0 220248 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_196
timestamp 1676037725
transform 1 0 219880 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_197
timestamp 1676037725
transform 1 0 217120 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_198
timestamp 1676037725
transform 1 0 214084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_199
timestamp 1676037725
transform 1 0 217304 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_200
timestamp 1676037725
transform 1 0 214544 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_201
timestamp 1676037725
transform 1 0 214728 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_202
timestamp 1676037725
transform 1 0 40020 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_203
timestamp 1676037725
transform 1 0 40020 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_204
timestamp 1676037725
transform 1 0 35880 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_205
timestamp 1676037725
transform 1 0 46092 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_206
timestamp 1676037725
transform 1 0 46644 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_207
timestamp 1676037725
transform 1 0 79764 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_208
timestamp 1676037725
transform 1 0 53636 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_209
timestamp 1676037725
transform 1 0 120336 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_210
timestamp 1676037725
transform 1 0 27324 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_211
timestamp 1676037725
transform 1 0 58512 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_212
timestamp 1676037725
transform 1 0 24656 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_213
timestamp 1676037725
transform 1 0 59248 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_214
timestamp 1676037725
transform 1 0 197800 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_215
timestamp 1676037725
transform 1 0 26128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_216
timestamp 1676037725
transform 1 0 202952 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_217
timestamp 1676037725
transform 1 0 236440 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_218
timestamp 1676037725
transform 1 0 24472 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_219
timestamp 1676037725
transform 1 0 53268 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_220
timestamp 1676037725
transform 1 0 89700 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_221
timestamp 1676037725
transform 1 0 121164 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_222
timestamp 1676037725
transform 1 0 155388 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_223
timestamp 1676037725
transform 1 0 27140 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_224
timestamp 1676037725
transform 1 0 191176 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_225
timestamp 1676037725
transform 1 0 223836 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_226
timestamp 1676037725
transform 1 0 89332 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_227
timestamp 1676037725
transform 1 0 123188 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_228
timestamp 1676037725
transform 1 0 24564 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_229
timestamp 1676037725
transform 1 0 53452 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_230
timestamp 1676037725
transform 1 0 87676 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_231
timestamp 1676037725
transform 1 0 24840 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_232
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_233
timestamp 1676037725
transform 1 0 202676 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_234
timestamp 1676037725
transform 1 0 236440 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_235
timestamp 1676037725
transform 1 0 188416 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_236
timestamp 1676037725
transform 1 0 259256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_237
timestamp 1676037725
transform 1 0 89700 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_238
timestamp 1676037725
transform 1 0 92184 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_239
timestamp 1676037725
transform 1 0 104236 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_240
timestamp 1676037725
transform 1 0 106996 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_241
timestamp 1676037725
transform 1 0 147752 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_242
timestamp 1676037725
transform 1 0 144992 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_243
timestamp 1676037725
transform 1 0 211876 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_244
timestamp 1676037725
transform 1 0 212612 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_245
timestamp 1676037725
transform 1 0 216936 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_246
timestamp 1676037725
transform 1 0 218224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_247
timestamp 1676037725
transform 1 0 87952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_248
timestamp 1676037725
transform 1 0 90436 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_249
timestamp 1676037725
transform 1 0 106536 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_250
timestamp 1676037725
transform 1 0 103776 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_251
timestamp 1676037725
transform 1 0 145176 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_252
timestamp 1676037725
transform 1 0 142416 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_253
timestamp 1676037725
transform 1 0 206816 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_254
timestamp 1676037725
transform 1 0 206448 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_255
timestamp 1676037725
transform 1 0 218684 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_256
timestamp 1676037725
transform 1 0 217120 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_257
timestamp 1676037725
transform 1 0 83076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_258
timestamp 1676037725
transform 1 0 85560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_259
timestamp 1676037725
transform 1 0 82708 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_260
timestamp 1676037725
transform 1 0 120980 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_261
timestamp 1676037725
transform 1 0 123464 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_262
timestamp 1676037725
transform 1 0 120612 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_263
timestamp 1676037725
transform 1 0 163208 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_264
timestamp 1676037725
transform 1 0 160448 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_265
timestamp 1676037725
transform 1 0 163576 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_266
timestamp 1676037725
transform 1 0 225308 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_267
timestamp 1676037725
transform 1 0 228068 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_268
timestamp 1676037725
transform 1 0 224940 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_269
timestamp 1676037725
transform 1 0 241868 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_270
timestamp 1676037725
transform 1 0 240304 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_271
timestamp 1676037725
transform 1 0 242604 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_272
timestamp 1676037725
transform 1 0 82984 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_273
timestamp 1676037725
transform 1 0 85468 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_274
timestamp 1676037725
transform 1 0 82616 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_275
timestamp 1676037725
transform 1 0 119692 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_276
timestamp 1676037725
transform 1 0 122452 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_277
timestamp 1676037725
transform 1 0 119324 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_278
timestamp 1676037725
transform 1 0 160448 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_279
timestamp 1676037725
transform 1 0 158056 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_280
timestamp 1676037725
transform 1 0 160816 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_281
timestamp 1676037725
transform 1 0 227608 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_282
timestamp 1676037725
transform 1 0 224848 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_283
timestamp 1676037725
transform 1 0 227976 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_284
timestamp 1676037725
transform 1 0 238648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_285
timestamp 1676037725
transform 1 0 239936 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_286
timestamp 1676037725
transform 1 0 238280 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_287
timestamp 1676037725
transform 1 0 91172 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_288
timestamp 1676037725
transform 1 0 90804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_289
timestamp 1676037725
transform 1 0 114540 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_290
timestamp 1676037725
transform 1 0 114908 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_291
timestamp 1676037725
transform 1 0 150788 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_292
timestamp 1676037725
transform 1 0 153272 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_293
timestamp 1676037725
transform 1 0 215280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_294
timestamp 1676037725
transform 1 0 217764 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_295
timestamp 1676037725
transform 1 0 252172 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_296
timestamp 1676037725
transform 1 0 250608 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_297
timestamp 1676037725
transform 1 0 170108 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_298
timestamp 1676037725
transform 1 0 219880 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_299
timestamp 1676037725
transform 1 0 46920 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_300
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_301
timestamp 1676037725
transform 1 0 58512 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_302
timestamp 1676037725
transform 1 0 83812 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_303
timestamp 1676037725
transform 1 0 123832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_304
timestamp 1676037725
transform 1 0 160448 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_305
timestamp 1676037725
transform 1 0 228620 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_306
timestamp 1676037725
transform 1 0 242236 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_307
timestamp 1676037725
transform 1 0 80684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_308
timestamp 1676037725
transform 1 0 120980 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_309
timestamp 1676037725
transform 1 0 160080 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_310
timestamp 1676037725
transform 1 0 225768 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_311
timestamp 1676037725
transform 1 0 241868 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_312
timestamp 1676037725
transform 1 0 91540 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_313
timestamp 1676037725
transform 1 0 112424 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_314
timestamp 1676037725
transform 1 0 152720 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_315
timestamp 1676037725
transform 1 0 218500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_316
timestamp 1676037725
transform 1 0 257968 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_317
timestamp 1676037725
transform 1 0 87952 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_318
timestamp 1676037725
transform 1 0 87584 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_319
timestamp 1676037725
transform 1 0 111504 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_320
timestamp 1676037725
transform 1 0 115644 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_321
timestamp 1676037725
transform 1 0 157688 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_322
timestamp 1676037725
transform 1 0 157688 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_323
timestamp 1676037725
transform 1 0 218132 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_324
timestamp 1676037725
transform 1 0 221720 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_325
timestamp 1676037725
transform 1 0 255760 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_326
timestamp 1676037725
transform 1 0 259440 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_327
timestamp 1676037725
transform 1 0 162104 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_328
timestamp 1676037725
transform 1 0 42688 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_329
timestamp 1676037725
transform 1 0 44436 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[0\].cell0_I openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 51888 0 1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[1\].cell0_I
timestamp 1676037725
transform 1 0 50784 0 -1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[2\].cell0_I
timestamp 1676037725
transform 1 0 50416 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[3\].cell0_I
timestamp 1676037725
transform 1 0 50324 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[4\].cell0_I
timestamp 1676037725
transform 1 0 48760 0 -1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[5\].cell0_I
timestamp 1676037725
transform 1 0 47288 0 1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[6\].cell0_I
timestamp 1676037725
transform 1 0 46460 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[7\].cell0_I
timestamp 1676037725
transform 1 0 46368 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[8\].cell0_I
timestamp 1676037725
transform 1 0 45632 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[9\].cell0_I
timestamp 1676037725
transform 1 0 44804 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[10\].cell0_I
timestamp 1676037725
transform 1 0 43056 0 1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[11\].cell0_I
timestamp 1676037725
transform 1 0 43148 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[12\].cell0_I
timestamp 1676037725
transform 1 0 42596 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[13\].cell0_I
timestamp 1676037725
transform 1 0 42780 0 1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[14\].cell0_I
timestamp 1676037725
transform 1 0 40756 0 1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[15\].cell0_I
timestamp 1676037725
transform 1 0 41032 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[16\].cell0_I
timestamp 1676037725
transform 1 0 40388 0 -1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[17\].cell0_I
timestamp 1676037725
transform 1 0 39652 0 -1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[18\].cell0_I
timestamp 1676037725
transform 1 0 38824 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[19\].cell0_I
timestamp 1676037725
transform 1 0 37628 0 -1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[20\].cell0_I
timestamp 1676037725
transform 1 0 37444 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[21\].cell0_I
timestamp 1676037725
transform 1 0 36708 0 1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[22\].cell0_I
timestamp 1676037725
transform 1 0 36248 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  col\[0\].genblk1.mux4_I\[23\].cell0_I
timestamp 1676037725
transform 1 0 35328 0 -1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__inv_2  col\[0\].genblk1.tbuf_row_ena_I.cell0_I
timestamp 1676037725
transform 1 0 94392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[0\].cell0_I openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 84732 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[1\].cell0_I
timestamp 1676037725
transform 1 0 81420 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[2\].cell0_I
timestamp 1676037725
transform 1 0 83444 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[3\].cell0_I
timestamp 1676037725
transform 1 0 83352 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[4\].cell0_I
timestamp 1676037725
transform 1 0 81696 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[5\].cell0_I
timestamp 1676037725
transform 1 0 81420 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[6\].cell0_I
timestamp 1676037725
transform 1 0 83996 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[7\].cell0_I
timestamp 1676037725
transform 1 0 87860 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[8\].cell0_I
timestamp 1676037725
transform 1 0 89424 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[9\].cell0_I
timestamp 1676037725
transform 1 0 91540 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[10\].cell0_I
timestamp 1676037725
transform 1 0 92460 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[11\].cell0_I
timestamp 1676037725
transform 1 0 91724 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[12\].cell0_I
timestamp 1676037725
transform 1 0 92644 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[13\].cell0_I
timestamp 1676037725
transform 1 0 94208 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[14\].cell0_I
timestamp 1676037725
transform 1 0 94300 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[15\].cell0_I
timestamp 1676037725
transform 1 0 94024 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[16\].cell0_I
timestamp 1676037725
transform 1 0 91724 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[17\].cell0_I
timestamp 1676037725
transform 1 0 90068 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[18\].cell0_I
timestamp 1676037725
transform 1 0 88320 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[19\].cell0_I
timestamp 1676037725
transform 1 0 86572 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[20\].cell0_I
timestamp 1676037725
transform 1 0 84732 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[21\].cell0_I
timestamp 1676037725
transform 1 0 84272 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[22\].cell0_I
timestamp 1676037725
transform 1 0 83536 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[0\].genblk1.tbuf_spine_ow_I\[23\].cell0_I
timestamp 1676037725
transform 1 0 83812 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  col\[0\].zbuf_bot_ena_I.genblk1.cell0_I_536 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 32292 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 32200 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 31372 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 30360 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 29440 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 28612 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 27968 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 27140 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 26680 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 25852 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 27692 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 24840 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 24288 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 23460 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 24932 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 25208 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 24932 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 26036 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_bot_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 27324 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[0\].zbuf_top_ena_I.genblk1.cell0_I_537
timestamp 1676037725
transform 1 0 33120 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 32292 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 31832 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 31004 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 29992 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 28796 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 28336 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 27784 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 26220 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 26496 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 26220 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 27324 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 24840 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 23828 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 23644 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 22816 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 25208 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 23644 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 26036 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[0\].zbuf_top_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 24840 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[1\].zbuf_bot_ena_I.genblk1.cell0_I_538
timestamp 1676037725
transform 1 0 66608 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 66516 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 65688 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 64860 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 64032 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 63204 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 62284 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 61456 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 60628 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 59800 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 59616 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 58880 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 57868 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 57132 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 56304 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 55476 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 54648 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 53820 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 53912 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_bot_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 53728 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[1\].zbuf_top_ena_I.genblk1.cell0_I_539
timestamp 1676037725
transform 1 0 67436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 66608 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 65964 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 64860 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 64032 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 63204 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 62376 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 61548 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 60720 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 60352 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 59616 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 58788 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 57960 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 57132 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 56304 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 55476 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 54556 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 53728 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 53728 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[1\].zbuf_top_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 53636 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[0\].cell0_I openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 120060 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[1\].cell0_I
timestamp 1676037725
transform 1 0 119140 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[2\].cell0_I
timestamp 1676037725
transform 1 0 118220 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[3\].cell0_I
timestamp 1676037725
transform 1 0 117392 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[4\].cell0_I
timestamp 1676037725
transform 1 0 114908 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[5\].cell0_I
timestamp 1676037725
transform 1 0 114632 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[6\].cell0_I
timestamp 1676037725
transform 1 0 112332 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[7\].cell0_I
timestamp 1676037725
transform 1 0 111780 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[8\].cell0_I
timestamp 1676037725
transform 1 0 109756 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[9\].cell0_I
timestamp 1676037725
transform 1 0 109572 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[10\].cell0_I
timestamp 1676037725
transform 1 0 108100 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[11\].cell0_I
timestamp 1676037725
transform 1 0 106444 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[12\].cell0_I
timestamp 1676037725
transform 1 0 104512 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[13\].cell0_I
timestamp 1676037725
transform 1 0 107180 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[14\].cell0_I
timestamp 1676037725
transform 1 0 106996 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[15\].cell0_I
timestamp 1676037725
transform 1 0 106076 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[16\].cell0_I
timestamp 1676037725
transform 1 0 104880 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[17\].cell0_I
timestamp 1676037725
transform 1 0 103408 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[18\].cell0_I
timestamp 1676037725
transform 1 0 101660 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[19\].cell0_I
timestamp 1676037725
transform 1 0 99636 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[20\].cell0_I
timestamp 1676037725
transform 1 0 99360 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[21\].cell0_I
timestamp 1676037725
transform 1 0 96876 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[22\].cell0_I
timestamp 1676037725
transform 1 0 96692 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[2\].genblk1.mux4_I\[23\].cell0_I
timestamp 1676037725
transform 1 0 96600 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  col\[2\].genblk1.tbuf_row_ena_I.cell0_I
timestamp 1676037725
transform 1 0 101016 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[0\].cell0_I
timestamp 1676037725
transform 1 0 122452 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[1\].cell0_I
timestamp 1676037725
transform 1 0 121716 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[2\].cell0_I
timestamp 1676037725
transform 1 0 121348 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[3\].cell0_I
timestamp 1676037725
transform 1 0 120060 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[4\].cell0_I
timestamp 1676037725
transform 1 0 117484 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[5\].cell0_I
timestamp 1676037725
transform 1 0 116472 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[6\].cell0_I
timestamp 1676037725
transform 1 0 115092 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[7\].cell0_I
timestamp 1676037725
transform 1 0 114080 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[8\].cell0_I
timestamp 1676037725
transform 1 0 113160 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[9\].cell0_I
timestamp 1676037725
transform 1 0 112424 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[10\].cell0_I
timestamp 1676037725
transform 1 0 110860 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[11\].cell0_I
timestamp 1676037725
transform 1 0 109020 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[12\].cell0_I
timestamp 1676037725
transform 1 0 106904 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[13\].cell0_I
timestamp 1676037725
transform 1 0 110216 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[14\].cell0_I
timestamp 1676037725
transform 1 0 109112 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[15\].cell0_I
timestamp 1676037725
transform 1 0 108468 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[16\].cell0_I
timestamp 1676037725
transform 1 0 107088 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[17\].cell0_I
timestamp 1676037725
transform 1 0 104604 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[18\].cell0_I
timestamp 1676037725
transform 1 0 104420 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[19\].cell0_I
timestamp 1676037725
transform 1 0 101936 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[20\].cell0_I
timestamp 1676037725
transform 1 0 101752 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[21\].cell0_I
timestamp 1676037725
transform 1 0 99452 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[22\].cell0_I
timestamp 1676037725
transform 1 0 99360 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[2\].genblk1.tbuf_spine_ow_I\[23\].cell0_I
timestamp 1676037725
transform 1 0 99360 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 100280 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[2\].zbuf_bot_ena_I.genblk1.cell0_I_540
timestamp 1676037725
transform 1 0 99268 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 99912 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 98348 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 98348 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 97520 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 96692 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 95864 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 95036 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 94760 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 94116 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 93196 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 92368 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 91540 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 90712 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 89884 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 89056 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 88044 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 88964 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_bot_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 88044 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 99820 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[2\].zbuf_top_ena_I.genblk1.cell0_I_541
timestamp 1676037725
transform 1 0 100096 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 99268 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 99268 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 98440 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 97612 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 96784 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 96416 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 95772 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 94944 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 94116 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 93288 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 93104 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 92460 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 91632 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 90620 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 89792 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 89700 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 88964 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[2\].zbuf_top_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 89056 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[3\].zbuf_bot_ena_I.genblk1.cell0_I_542
timestamp 1676037725
transform 1 0 134964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 134044 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 133952 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 133216 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 132940 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 132204 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 131284 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 130456 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 129260 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 128432 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 128248 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 127512 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 126684 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 125856 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 125028 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 124108 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 123280 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 122452 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 121624 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_bot_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 120796 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[3\].zbuf_top_ena_I.genblk1.cell0_I_543
timestamp 1676037725
transform 1 0 135424 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 134136 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 133860 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 133032 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 132940 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 131836 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 131008 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 130548 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 130180 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 129076 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 128340 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 127604 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 126684 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 125856 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 125028 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 124200 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 123372 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 122544 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 121532 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[3\].zbuf_top_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 121532 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[0\].cell0_I
timestamp 1676037725
transform 1 0 158332 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[1\].cell0_I
timestamp 1676037725
transform 1 0 157872 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[2\].cell0_I
timestamp 1676037725
transform 1 0 158240 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[3\].cell0_I
timestamp 1676037725
transform 1 0 155940 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[4\].cell0_I
timestamp 1676037725
transform 1 0 155664 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[5\].cell0_I
timestamp 1676037725
transform 1 0 153180 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[6\].cell0_I
timestamp 1676037725
transform 1 0 151708 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[7\].cell0_I
timestamp 1676037725
transform 1 0 150604 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[8\].cell0_I
timestamp 1676037725
transform 1 0 150512 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[9\].cell0_I
timestamp 1676037725
transform 1 0 150512 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[10\].cell0_I
timestamp 1676037725
transform 1 0 148212 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[11\].cell0_I
timestamp 1676037725
transform 1 0 145820 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[12\].cell0_I
timestamp 1676037725
transform 1 0 145636 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[13\].cell0_I
timestamp 1676037725
transform 1 0 148212 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[14\].cell0_I
timestamp 1676037725
transform 1 0 147936 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[15\].cell0_I
timestamp 1676037725
transform 1 0 145636 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[16\].cell0_I
timestamp 1676037725
transform 1 0 145360 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[17\].cell0_I
timestamp 1676037725
transform 1 0 143060 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[18\].cell0_I
timestamp 1676037725
transform 1 0 143060 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[19\].cell0_I
timestamp 1676037725
transform 1 0 142784 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[20\].cell0_I
timestamp 1676037725
transform 1 0 140668 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[21\].cell0_I
timestamp 1676037725
transform 1 0 140484 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[22\].cell0_I
timestamp 1676037725
transform 1 0 138092 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[4\].genblk1.mux4_I\[23\].cell0_I
timestamp 1676037725
transform 1 0 137724 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  col\[4\].genblk1.tbuf_row_ena_I.cell0_I
timestamp 1676037725
transform 1 0 161092 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[0\].cell0_I
timestamp 1676037725
transform 1 0 161000 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[1\].cell0_I
timestamp 1676037725
transform 1 0 160816 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[2\].cell0_I
timestamp 1676037725
transform 1 0 161092 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[3\].cell0_I
timestamp 1676037725
transform 1 0 158332 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[4\].cell0_I
timestamp 1676037725
transform 1 0 158240 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[5\].cell0_I
timestamp 1676037725
transform 1 0 155940 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[6\].cell0_I
timestamp 1676037725
transform 1 0 155664 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[7\].cell0_I
timestamp 1676037725
transform 1 0 153364 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[8\].cell0_I
timestamp 1676037725
transform 1 0 153088 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[9\].cell0_I
timestamp 1676037725
transform 1 0 151156 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[10\].cell0_I
timestamp 1676037725
transform 1 0 150788 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[11\].cell0_I
timestamp 1676037725
transform 1 0 148212 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[12\].cell0_I
timestamp 1676037725
transform 1 0 146464 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[13\].cell0_I
timestamp 1676037725
transform 1 0 150512 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[14\].cell0_I
timestamp 1676037725
transform 1 0 150788 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[15\].cell0_I
timestamp 1676037725
transform 1 0 148212 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[16\].cell0_I
timestamp 1676037725
transform 1 0 147936 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[17\].cell0_I
timestamp 1676037725
transform 1 0 145636 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[18\].cell0_I
timestamp 1676037725
transform 1 0 143060 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[19\].cell0_I
timestamp 1676037725
transform 1 0 141772 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[20\].cell0_I
timestamp 1676037725
transform 1 0 143060 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[21\].cell0_I
timestamp 1676037725
transform 1 0 140484 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[22\].cell0_I
timestamp 1676037725
transform 1 0 138920 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[4\].genblk1.tbuf_spine_ow_I\[23\].cell0_I
timestamp 1676037725
transform 1 0 138920 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  col\[4\].zbuf_bot_ena_I.genblk1.cell0_I_544
timestamp 1676037725
transform 1 0 167716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 167624 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 167900 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 166980 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 167072 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 166244 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 165232 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 164404 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 163668 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 163576 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 162748 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 161920 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 161092 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 159896 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 159344 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 159896 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 159068 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 158516 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 157228 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_bot_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 156400 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 169556 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[4\].zbuf_top_ena_I.genblk1.cell0_I_545
timestamp 1676037725
transform 1 0 169556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 167900 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 167900 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 167072 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 166244 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 165324 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 164496 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 164772 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 163668 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 162288 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 161368 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 161092 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 159804 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 158976 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 157964 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 157412 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 156492 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 156584 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[4\].zbuf_top_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 155756 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[5\].zbuf_bot_ena_I.genblk1.cell0_I_546
timestamp 1676037725
transform 1 0 202308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 202308 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 201940 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 202308 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 201204 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 201296 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 200468 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 199640 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 198812 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 197984 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 197064 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 197156 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 196144 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 195316 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 194488 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 193660 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 192832 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 192004 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 190992 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_bot_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 190716 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 203136 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[5\].zbuf_top_ena_I.genblk1.cell0_I_547
timestamp 1676037725
transform 1 0 202768 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 203044 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 202308 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 202032 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 201388 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 200560 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 199732 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 198444 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 198536 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 197156 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 196236 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 196236 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 195408 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 194580 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 193200 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 193200 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 192372 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 191544 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[5\].zbuf_top_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 190532 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[0\].cell0_I
timestamp 1676037725
transform 1 0 225492 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[1\].cell0_I
timestamp 1676037725
transform 1 0 224296 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[2\].cell0_I
timestamp 1676037725
transform 1 0 225492 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[3\].cell0_I
timestamp 1676037725
transform 1 0 222916 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[4\].cell0_I
timestamp 1676037725
transform 1 0 222640 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[5\].cell0_I
timestamp 1676037725
transform 1 0 220524 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[6\].cell0_I
timestamp 1676037725
transform 1 0 220156 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[7\].cell0_I
timestamp 1676037725
transform 1 0 220248 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[8\].cell0_I
timestamp 1676037725
transform 1 0 217764 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[9\].cell0_I
timestamp 1676037725
transform 1 0 217764 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[10\].cell0_I
timestamp 1676037725
transform 1 0 217948 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[11\].cell0_I
timestamp 1676037725
transform 1 0 215372 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[12\].cell0_I
timestamp 1676037725
transform 1 0 214452 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[13\].cell0_I
timestamp 1676037725
transform 1 0 215372 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[14\].cell0_I
timestamp 1676037725
transform 1 0 215188 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[15\].cell0_I
timestamp 1676037725
transform 1 0 214912 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[16\].cell0_I
timestamp 1676037725
transform 1 0 215188 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[17\].cell0_I
timestamp 1676037725
transform 1 0 212796 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[18\].cell0_I
timestamp 1676037725
transform 1 0 212428 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[19\].cell0_I
timestamp 1676037725
transform 1 0 212612 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[20\].cell0_I
timestamp 1676037725
transform 1 0 210220 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[21\].cell0_I
timestamp 1676037725
transform 1 0 210036 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[22\].cell0_I
timestamp 1676037725
transform 1 0 210036 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  col\[6\].genblk1.mux4_I\[23\].cell0_I
timestamp 1676037725
transform 1 0 207736 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__clkinv_4  col\[6\].genblk1.tbuf_row_ena_I.cell0_I openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 229908 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[0\].cell0_I
timestamp 1676037725
transform 1 0 228068 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[1\].cell0_I
timestamp 1676037725
transform 1 0 226504 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[2\].cell0_I
timestamp 1676037725
transform 1 0 225676 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[3\].cell0_I
timestamp 1676037725
transform 1 0 225492 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[4\].cell0_I
timestamp 1676037725
transform 1 0 223652 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[5\].cell0_I
timestamp 1676037725
transform 1 0 222824 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[6\].cell0_I
timestamp 1676037725
transform 1 0 221812 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[7\].cell0_I
timestamp 1676037725
transform 1 0 220616 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[8\].cell0_I
timestamp 1676037725
transform 1 0 219236 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[9\].cell0_I
timestamp 1676037725
transform 1 0 215648 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[10\].cell0_I
timestamp 1676037725
transform 1 0 214176 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[11\].cell0_I
timestamp 1676037725
transform 1 0 212796 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[12\].cell0_I
timestamp 1676037725
transform 1 0 212520 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[13\].cell0_I
timestamp 1676037725
transform 1 0 217488 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[14\].cell0_I
timestamp 1676037725
transform 1 0 213992 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[15\].cell0_I
timestamp 1676037725
transform 1 0 212336 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[16\].cell0_I
timestamp 1676037725
transform 1 0 210496 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[17\].cell0_I
timestamp 1676037725
transform 1 0 209760 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[18\].cell0_I
timestamp 1676037725
transform 1 0 207460 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[19\].cell0_I
timestamp 1676037725
transform 1 0 207184 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[20\].cell0_I
timestamp 1676037725
transform 1 0 207552 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[21\].cell0_I
timestamp 1676037725
transform 1 0 204884 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[22\].cell0_I
timestamp 1676037725
transform 1 0 204884 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  col\[6\].genblk1.tbuf_spine_ow_I\[23\].cell0_I
timestamp 1676037725
transform 1 0 204148 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  col\[6\].zbuf_bot_ena_I.genblk1.cell0_I_548
timestamp 1676037725
transform 1 0 235796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 236532 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 235796 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 235704 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 234876 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 234048 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 233220 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 232116 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 232208 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 231380 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 230552 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 229724 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 228896 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 228068 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 228068 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 226504 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 226596 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 225492 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 225768 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_bot_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 224940 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 235612 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[6\].zbuf_top_ena_I.genblk1.cell0_I_549
timestamp 1676037725
transform 1 0 235796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 235796 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 235796 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 234508 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 234508 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 233680 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 232852 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 232024 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 230644 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 229816 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 229632 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 228804 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 227976 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 227148 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 226320 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 225492 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 224572 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 224204 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[6\].zbuf_top_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 223928 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[7\].zbuf_bot_ena_I.genblk1.cell0_I_550
timestamp 1676037725
transform 1 0 265972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 270112 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 269284 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 269008 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 269284 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 268272 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 267444 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 266616 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 265788 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 264960 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 263948 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 264132 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 263120 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 262292 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 261464 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 260636 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 259808 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 258888 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 258980 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_bot_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 257692 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 269284 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  col\[7\].zbuf_top_ena_I.genblk1.cell0_I_551
timestamp 1676037725
transform 1 0 265972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 265512 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 264868 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 269284 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 267168 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 266340 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 265696 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 265788 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 264960 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 264132 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 263396 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 262568 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 261740 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 261556 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 260636 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 259992 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 258980 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 258980 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  col\[7\].zbuf_top_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 257784 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  fanout419
timestamp 1676037725
transform 1 0 258060 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout420
timestamp 1676037725
transform 1 0 263672 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout421
timestamp 1676037725
transform 1 0 230644 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout422
timestamp 1676037725
transform 1 0 230736 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout423
timestamp 1676037725
transform 1 0 190716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout424
timestamp 1676037725
transform 1 0 197248 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout425
timestamp 1676037725
transform 1 0 163116 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout426
timestamp 1676037725
transform 1 0 169096 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout427
timestamp 1676037725
transform 1 0 121624 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout428
timestamp 1676037725
transform 1 0 129260 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout429
timestamp 1676037725
transform 1 0 94668 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout430
timestamp 1676037725
transform 1 0 100096 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout431
timestamp 1676037725
transform 1 0 59616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout432
timestamp 1676037725
transform 1 0 66792 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout433
timestamp 1676037725
transform 1 0 26864 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout434
timestamp 1676037725
transform 1 0 32660 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  fanout435 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 215832 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  fanout436
timestamp 1676037725
transform 1 0 228252 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_8  fanout437 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 228804 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_12  fanout438
timestamp 1676037725
transform 1 0 148764 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  fanout439
timestamp 1676037725
transform 1 0 161092 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  fanout440
timestamp 1676037725
transform 1 0 161644 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  fanout441
timestamp 1676037725
transform 1 0 101936 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  fanout442
timestamp 1676037725
transform 1 0 111872 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  fanout443
timestamp 1676037725
transform 1 0 102120 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  fanout444
timestamp 1676037725
transform 1 0 86664 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  fanout445
timestamp 1676037725
transform 1 0 92736 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  fanout446
timestamp 1676037725
transform 1 0 94760 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout447
timestamp 1676037725
transform 1 0 41952 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout448
timestamp 1676037725
transform 1 0 47932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout449
timestamp 1676037725
transform 1 0 52900 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout450
timestamp 1676037725
transform 1 0 108376 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout451
timestamp 1676037725
transform 1 0 107640 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout452
timestamp 1676037725
transform 1 0 122176 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout453
timestamp 1676037725
transform 1 0 124936 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout454
timestamp 1676037725
transform 1 0 155204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout455
timestamp 1676037725
transform 1 0 155940 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout456
timestamp 1676037725
transform 1 0 162656 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout457
timestamp 1676037725
transform 1 0 217672 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout458
timestamp 1676037725
transform 1 0 219328 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout459
timestamp 1676037725
transform 1 0 230368 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout460
timestamp 1676037725
transform 1 0 232300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout461
timestamp 1676037725
transform 1 0 41584 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout462
timestamp 1676037725
transform 1 0 47840 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout463
timestamp 1676037725
transform 1 0 52900 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout464
timestamp 1676037725
transform 1 0 108836 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout465
timestamp 1676037725
transform 1 0 109756 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout466
timestamp 1676037725
transform 1 0 120704 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout467
timestamp 1676037725
transform 1 0 130180 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout468
timestamp 1676037725
transform 1 0 154560 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout469
timestamp 1676037725
transform 1 0 156860 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout470
timestamp 1676037725
transform 1 0 170200 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout471
timestamp 1676037725
transform 1 0 216384 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout472
timestamp 1676037725
transform 1 0 218592 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout473
timestamp 1676037725
transform 1 0 230092 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout474
timestamp 1676037725
transform 1 0 230184 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout475
timestamp 1676037725
transform 1 0 162104 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout476
timestamp 1676037725
transform 1 0 263120 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout477
timestamp 1676037725
transform 1 0 162196 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout478
timestamp 1676037725
transform 1 0 264132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout479
timestamp 1676037725
transform 1 0 163668 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout480
timestamp 1676037725
transform 1 0 265144 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout481
timestamp 1676037725
transform 1 0 163576 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout482
timestamp 1676037725
transform 1 0 265052 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout483
timestamp 1676037725
transform 1 0 164220 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout484
timestamp 1676037725
transform 1 0 265972 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout485 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 164956 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  fanout486
timestamp 1676037725
transform 1 0 266708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout487
timestamp 1676037725
transform 1 0 166428 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  fanout488
timestamp 1676037725
transform 1 0 266984 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout489
timestamp 1676037725
transform 1 0 166612 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  fanout490
timestamp 1676037725
transform 1 0 268088 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout491
timestamp 1676037725
transform 1 0 168084 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  fanout492
timestamp 1676037725
transform 1 0 268272 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout493
timestamp 1676037725
transform 1 0 156492 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout494
timestamp 1676037725
transform 1 0 257968 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout495
timestamp 1676037725
transform 1 0 156676 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout496
timestamp 1676037725
transform 1 0 257784 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout497
timestamp 1676037725
transform 1 0 157872 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout498
timestamp 1676037725
transform 1 0 258980 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout499
timestamp 1676037725
transform 1 0 158516 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout500
timestamp 1676037725
transform 1 0 259992 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout501
timestamp 1676037725
transform 1 0 158516 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout502
timestamp 1676037725
transform 1 0 261556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout503
timestamp 1676037725
transform 1 0 159712 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout504
timestamp 1676037725
transform 1 0 261188 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout505
timestamp 1676037725
transform 1 0 160724 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout506
timestamp 1676037725
transform 1 0 262476 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout507
timestamp 1676037725
transform 1 0 161092 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout508
timestamp 1676037725
transform 1 0 262384 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout509
timestamp 1676037725
transform 1 0 168820 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  fanout510
timestamp 1676037725
transform 1 0 267168 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout511
timestamp 1676037725
transform 1 0 226596 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout512
timestamp 1676037725
transform 1 0 239292 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout513
timestamp 1676037725
transform 1 0 240212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout514
timestamp 1676037725
transform 1 0 269192 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  fanout515
timestamp 1676037725
transform 1 0 264868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout516
timestamp 1676037725
transform 1 0 264776 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_3 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_8 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1840 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26
timestamp 1676037725
transform 1 0 3496 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29
timestamp 1676037725
transform 1 0 3772 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_35
timestamp 1676037725
transform 1 0 4324 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_43 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5060 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54
timestamp 1676037725
transform 1 0 6072 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1676037725
transform 1 0 6348 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_69
timestamp 1676037725
transform 1 0 7452 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_85 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8924 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_89
timestamp 1676037725
transform 1 0 9292 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_94
timestamp 1676037725
transform 1 0 9752 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_102
timestamp 1676037725
transform 1 0 10488 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_110
timestamp 1676037725
transform 1 0 11224 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_113
timestamp 1676037725
transform 1 0 11500 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_121
timestamp 1676037725
transform 1 0 12236 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_129
timestamp 1676037725
transform 1 0 12972 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1676037725
transform 1 0 13708 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_141
timestamp 1676037725
transform 1 0 14076 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_159
timestamp 1676037725
transform 1 0 15732 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1676037725
transform 1 0 16468 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_169
timestamp 1676037725
transform 1 0 16652 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_177
timestamp 1676037725
transform 1 0 17388 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_185
timestamp 1676037725
transform 1 0 18124 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1676037725
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19228 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1676037725
transform 1 0 20332 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1676037725
transform 1 0 21436 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1676037725
transform 1 0 21804 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_237
timestamp 1676037725
transform 1 0 22908 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_245
timestamp 1676037725
transform 1 0 23644 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_250
timestamp 1676037725
transform 1 0 24104 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_253
timestamp 1676037725
transform 1 0 24380 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_257
timestamp 1676037725
transform 1 0 24748 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_264
timestamp 1676037725
transform 1 0 25392 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_274 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26312 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_281
timestamp 1676037725
transform 1 0 26956 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_288
timestamp 1676037725
transform 1 0 27600 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_297
timestamp 1676037725
transform 1 0 28428 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_301
timestamp 1676037725
transform 1 0 28796 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_306
timestamp 1676037725
transform 1 0 29256 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_309
timestamp 1676037725
transform 1 0 29532 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_315
timestamp 1676037725
transform 1 0 30084 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_319
timestamp 1676037725
transform 1 0 30452 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_324
timestamp 1676037725
transform 1 0 30912 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_328
timestamp 1676037725
transform 1 0 31280 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1676037725
transform 1 0 31740 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_337
timestamp 1676037725
transform 1 0 32108 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_343
timestamp 1676037725
transform 1 0 32660 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_355
timestamp 1676037725
transform 1 0 33764 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_362
timestamp 1676037725
transform 1 0 34408 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_365
timestamp 1676037725
transform 1 0 34684 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_376
timestamp 1676037725
transform 1 0 35696 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_383
timestamp 1676037725
transform 1 0 36340 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_390
timestamp 1676037725
transform 1 0 36984 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_393
timestamp 1676037725
transform 1 0 37260 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_404
timestamp 1676037725
transform 1 0 38272 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_411
timestamp 1676037725
transform 1 0 38916 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_418
timestamp 1676037725
transform 1 0 39560 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_421
timestamp 1676037725
transform 1 0 39836 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_432
timestamp 1676037725
transform 1 0 40848 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_439
timestamp 1676037725
transform 1 0 41492 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_446
timestamp 1676037725
transform 1 0 42136 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_449
timestamp 1676037725
transform 1 0 42412 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_455
timestamp 1676037725
transform 1 0 42964 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_459
timestamp 1676037725
transform 1 0 43332 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_463
timestamp 1676037725
transform 1 0 43700 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_467
timestamp 1676037725
transform 1 0 44068 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_474
timestamp 1676037725
transform 1 0 44712 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_477
timestamp 1676037725
transform 1 0 44988 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_488
timestamp 1676037725
transform 1 0 46000 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_495
timestamp 1676037725
transform 1 0 46644 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_502
timestamp 1676037725
transform 1 0 47288 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_505
timestamp 1676037725
transform 1 0 47564 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_511
timestamp 1676037725
transform 1 0 48116 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_515
timestamp 1676037725
transform 1 0 48484 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_519
timestamp 1676037725
transform 1 0 48852 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_523
timestamp 1676037725
transform 1 0 49220 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_530
timestamp 1676037725
transform 1 0 49864 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_533
timestamp 1676037725
transform 1 0 50140 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_544
timestamp 1676037725
transform 1 0 51152 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_551
timestamp 1676037725
transform 1 0 51796 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_558
timestamp 1676037725
transform 1 0 52440 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_561
timestamp 1676037725
transform 1 0 52716 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_565
timestamp 1676037725
transform 1 0 53084 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_570
timestamp 1676037725
transform 1 0 53544 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_579
timestamp 1676037725
transform 1 0 54372 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_587
timestamp 1676037725
transform 1 0 55108 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_589
timestamp 1676037725
transform 1 0 55292 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_601
timestamp 1676037725
transform 1 0 56396 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_605
timestamp 1676037725
transform 1 0 56764 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_610
timestamp 1676037725
transform 1 0 57224 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_617
timestamp 1676037725
transform 1 0 57868 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_627
timestamp 1676037725
transform 1 0 58788 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_631
timestamp 1676037725
transform 1 0 59156 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_634
timestamp 1676037725
transform 1 0 59432 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_641
timestamp 1676037725
transform 1 0 60076 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_645
timestamp 1676037725
transform 1 0 60444 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_651
timestamp 1676037725
transform 1 0 60996 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_659
timestamp 1676037725
transform 1 0 61732 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_667
timestamp 1676037725
transform 1 0 62468 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_671
timestamp 1676037725
transform 1 0 62836 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_673
timestamp 1676037725
transform 1 0 63020 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_683
timestamp 1676037725
transform 1 0 63940 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_691
timestamp 1676037725
transform 1 0 64676 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_699
timestamp 1676037725
transform 1 0 65412 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_701
timestamp 1676037725
transform 1 0 65596 0 1 1088
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_709
timestamp 1676037725
transform 1 0 66332 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_721
timestamp 1676037725
transform 1 0 67436 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_727
timestamp 1676037725
transform 1 0 67988 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_729
timestamp 1676037725
transform 1 0 68172 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_740
timestamp 1676037725
transform 1 0 69184 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_754
timestamp 1676037725
transform 1 0 70472 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_757
timestamp 1676037725
transform 1 0 70748 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_769
timestamp 1676037725
transform 1 0 71852 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_782
timestamp 1676037725
transform 1 0 73048 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_785
timestamp 1676037725
transform 1 0 73324 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_797
timestamp 1676037725
transform 1 0 74428 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_810
timestamp 1676037725
transform 1 0 75624 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_813
timestamp 1676037725
transform 1 0 75900 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_825
timestamp 1676037725
transform 1 0 77004 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_838
timestamp 1676037725
transform 1 0 78200 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_841
timestamp 1676037725
transform 1 0 78476 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_853
timestamp 1676037725
transform 1 0 79580 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_866
timestamp 1676037725
transform 1 0 80776 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_869
timestamp 1676037725
transform 1 0 81052 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_881
timestamp 1676037725
transform 1 0 82156 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_894
timestamp 1676037725
transform 1 0 83352 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_897
timestamp 1676037725
transform 1 0 83628 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_909
timestamp 1676037725
transform 1 0 84732 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_922
timestamp 1676037725
transform 1 0 85928 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_925
timestamp 1676037725
transform 1 0 86204 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_941
timestamp 1676037725
transform 1 0 87676 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_950
timestamp 1676037725
transform 1 0 88504 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_953
timestamp 1676037725
transform 1 0 88780 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_960
timestamp 1676037725
transform 1 0 89424 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_968
timestamp 1676037725
transform 1 0 90160 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_975
timestamp 1676037725
transform 1 0 90804 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_979
timestamp 1676037725
transform 1 0 91172 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_981
timestamp 1676037725
transform 1 0 91356 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_987
timestamp 1676037725
transform 1 0 91908 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_992
timestamp 1676037725
transform 1 0 92368 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1000
timestamp 1676037725
transform 1 0 93104 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1006
timestamp 1676037725
transform 1 0 93656 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1009
timestamp 1676037725
transform 1 0 93932 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1017
timestamp 1676037725
transform 1 0 94668 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1023
timestamp 1676037725
transform 1 0 95220 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1029
timestamp 1676037725
transform 1 0 95772 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1034
timestamp 1676037725
transform 1 0 96232 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1037
timestamp 1676037725
transform 1 0 96508 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1045
timestamp 1676037725
transform 1 0 97244 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1053
timestamp 1676037725
transform 1 0 97980 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1062
timestamp 1676037725
transform 1 0 98808 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1065
timestamp 1676037725
transform 1 0 99084 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1070
timestamp 1676037725
transform 1 0 99544 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1079
timestamp 1676037725
transform 1 0 100372 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1087
timestamp 1676037725
transform 1 0 101108 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1091
timestamp 1676037725
transform 1 0 101476 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1093
timestamp 1676037725
transform 1 0 101660 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1105
timestamp 1676037725
transform 1 0 102764 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1111
timestamp 1676037725
transform 1 0 103316 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1118
timestamp 1676037725
transform 1 0 103960 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1121
timestamp 1676037725
transform 1 0 104236 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1125
timestamp 1676037725
transform 1 0 104604 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1129
timestamp 1676037725
transform 1 0 104972 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1133
timestamp 1676037725
transform 1 0 105340 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1137
timestamp 1676037725
transform 1 0 105708 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1141
timestamp 1676037725
transform 1 0 106076 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1145
timestamp 1676037725
transform 1 0 106444 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1149
timestamp 1676037725
transform 1 0 106812 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1160
timestamp 1676037725
transform 1 0 107824 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1167
timestamp 1676037725
transform 1 0 108468 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1174
timestamp 1676037725
transform 1 0 109112 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1177
timestamp 1676037725
transform 1 0 109388 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1181
timestamp 1676037725
transform 1 0 109756 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1185
timestamp 1676037725
transform 1 0 110124 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1189
timestamp 1676037725
transform 1 0 110492 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1193
timestamp 1676037725
transform 1 0 110860 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1197
timestamp 1676037725
transform 1 0 111228 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1201
timestamp 1676037725
transform 1 0 111596 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1205
timestamp 1676037725
transform 1 0 111964 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1216
timestamp 1676037725
transform 1 0 112976 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1223
timestamp 1676037725
transform 1 0 113620 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1230
timestamp 1676037725
transform 1 0 114264 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1233
timestamp 1676037725
transform 1 0 114540 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1237
timestamp 1676037725
transform 1 0 114908 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1241
timestamp 1676037725
transform 1 0 115276 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1245
timestamp 1676037725
transform 1 0 115644 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1249
timestamp 1676037725
transform 1 0 116012 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1253
timestamp 1676037725
transform 1 0 116380 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1257
timestamp 1676037725
transform 1 0 116748 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1261
timestamp 1676037725
transform 1 0 117116 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1272
timestamp 1676037725
transform 1 0 118128 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1279
timestamp 1676037725
transform 1 0 118772 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1286
timestamp 1676037725
transform 1 0 119416 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1289
timestamp 1676037725
transform 1 0 119692 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1293
timestamp 1676037725
transform 1 0 120060 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1297
timestamp 1676037725
transform 1 0 120428 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1301
timestamp 1676037725
transform 1 0 120796 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1305
timestamp 1676037725
transform 1 0 121164 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1309
timestamp 1676037725
transform 1 0 121532 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1314
timestamp 1676037725
transform 1 0 121992 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1317
timestamp 1676037725
transform 1 0 122268 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1323
timestamp 1676037725
transform 1 0 122820 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1328
timestamp 1676037725
transform 1 0 123280 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1332
timestamp 1676037725
transform 1 0 123648 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1337
timestamp 1676037725
transform 1 0 124108 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1343
timestamp 1676037725
transform 1 0 124660 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1345
timestamp 1676037725
transform 1 0 124844 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1355
timestamp 1676037725
transform 1 0 125764 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1363
timestamp 1676037725
transform 1 0 126500 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1370
timestamp 1676037725
transform 1 0 127144 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1373
timestamp 1676037725
transform 1 0 127420 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1381
timestamp 1676037725
transform 1 0 128156 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1387
timestamp 1676037725
transform 1 0 128708 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1395
timestamp 1676037725
transform 1 0 129444 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1399
timestamp 1676037725
transform 1 0 129812 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1401
timestamp 1676037725
transform 1 0 129996 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1407
timestamp 1676037725
transform 1 0 130548 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1412
timestamp 1676037725
transform 1 0 131008 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1420
timestamp 1676037725
transform 1 0 131744 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1426
timestamp 1676037725
transform 1 0 132296 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1429
timestamp 1676037725
transform 1 0 132572 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1438
timestamp 1676037725
transform 1 0 133400 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1449
timestamp 1676037725
transform 1 0 134412 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1455
timestamp 1676037725
transform 1 0 134964 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1457
timestamp 1676037725
transform 1 0 135148 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1469
timestamp 1676037725
transform 1 0 136252 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1481
timestamp 1676037725
transform 1 0 137356 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1485
timestamp 1676037725
transform 1 0 137724 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1490
timestamp 1676037725
transform 1 0 138184 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1497
timestamp 1676037725
transform 1 0 138828 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1504
timestamp 1676037725
transform 1 0 139472 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1513
timestamp 1676037725
transform 1 0 140300 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1518
timestamp 1676037725
transform 1 0 140760 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1525
timestamp 1676037725
transform 1 0 141404 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1532
timestamp 1676037725
transform 1 0 142048 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1541
timestamp 1676037725
transform 1 0 142876 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1546
timestamp 1676037725
transform 1 0 143336 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1553
timestamp 1676037725
transform 1 0 143980 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1560
timestamp 1676037725
transform 1 0 144624 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1569
timestamp 1676037725
transform 1 0 145452 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1574
timestamp 1676037725
transform 1 0 145912 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1581
timestamp 1676037725
transform 1 0 146556 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1588
timestamp 1676037725
transform 1 0 147200 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1597
timestamp 1676037725
transform 1 0 148028 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1602
timestamp 1676037725
transform 1 0 148488 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1609
timestamp 1676037725
transform 1 0 149132 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1616
timestamp 1676037725
transform 1 0 149776 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1625
timestamp 1676037725
transform 1 0 150604 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1630
timestamp 1676037725
transform 1 0 151064 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1637
timestamp 1676037725
transform 1 0 151708 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1644
timestamp 1676037725
transform 1 0 152352 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1653
timestamp 1676037725
transform 1 0 153180 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1658
timestamp 1676037725
transform 1 0 153640 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1665
timestamp 1676037725
transform 1 0 154284 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1672
timestamp 1676037725
transform 1 0 154928 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1681
timestamp 1676037725
transform 1 0 155756 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1687
timestamp 1676037725
transform 1 0 156308 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1693
timestamp 1676037725
transform 1 0 156860 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1702
timestamp 1676037725
transform 1 0 157688 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1709
timestamp 1676037725
transform 1 0 158332 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1716
timestamp 1676037725
transform 1 0 158976 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1725
timestamp 1676037725
transform 1 0 159804 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1733
timestamp 1676037725
transform 1 0 160540 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1737
timestamp 1676037725
transform 1 0 160908 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1743
timestamp 1676037725
transform 1 0 161460 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1751
timestamp 1676037725
transform 1 0 162196 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1756
timestamp 1676037725
transform 1 0 162656 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1765
timestamp 1676037725
transform 1 0 163484 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1772
timestamp 1676037725
transform 1 0 164128 0 1 1088
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1780
timestamp 1676037725
transform 1 0 164864 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1793
timestamp 1676037725
transform 1 0 166060 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1801
timestamp 1676037725
transform 1 0 166796 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1808
timestamp 1676037725
transform 1 0 167440 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1816
timestamp 1676037725
transform 1 0 168176 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1821
timestamp 1676037725
transform 1 0 168636 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1827
timestamp 1676037725
transform 1 0 169188 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_1839
timestamp 1676037725
transform 1 0 170292 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1847
timestamp 1676037725
transform 1 0 171028 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1849
timestamp 1676037725
transform 1 0 171212 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1855
timestamp 1676037725
transform 1 0 171764 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1859
timestamp 1676037725
transform 1 0 172132 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1870
timestamp 1676037725
transform 1 0 173144 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1877
timestamp 1676037725
transform 1 0 173788 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1889
timestamp 1676037725
transform 1 0 174892 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1901
timestamp 1676037725
transform 1 0 175996 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1905
timestamp 1676037725
transform 1 0 176364 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_1917
timestamp 1676037725
transform 1 0 177468 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_1929
timestamp 1676037725
transform 1 0 178572 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1933
timestamp 1676037725
transform 1 0 178940 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1945
timestamp 1676037725
transform 1 0 180044 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1953
timestamp 1676037725
transform 1 0 180780 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1959
timestamp 1676037725
transform 1 0 181332 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1961
timestamp 1676037725
transform 1 0 181516 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_1967
timestamp 1676037725
transform 1 0 182068 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_1971
timestamp 1676037725
transform 1 0 182436 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_1982
timestamp 1676037725
transform 1 0 183448 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_1989
timestamp 1676037725
transform 1 0 184092 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_2001
timestamp 1676037725
transform 1 0 185196 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_2013
timestamp 1676037725
transform 1 0 186300 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2017
timestamp 1676037725
transform 1 0 186668 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_2029
timestamp 1676037725
transform 1 0 187772 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_2041
timestamp 1676037725
transform 1 0 188876 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2045
timestamp 1676037725
transform 1 0 189244 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2057
timestamp 1676037725
transform 1 0 190348 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2063
timestamp 1676037725
transform 1 0 190900 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_2069
timestamp 1676037725
transform 1 0 191452 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2073
timestamp 1676037725
transform 1 0 191820 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2079
timestamp 1676037725
transform 1 0 192372 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2084
timestamp 1676037725
transform 1 0 192832 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2088
timestamp 1676037725
transform 1 0 193200 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2093
timestamp 1676037725
transform 1 0 193660 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2099
timestamp 1676037725
transform 1 0 194212 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2101
timestamp 1676037725
transform 1 0 194396 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2107
timestamp 1676037725
transform 1 0 194948 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2113
timestamp 1676037725
transform 1 0 195500 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2118
timestamp 1676037725
transform 1 0 195960 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2126
timestamp 1676037725
transform 1 0 196696 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2129
timestamp 1676037725
transform 1 0 196972 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2135
timestamp 1676037725
transform 1 0 197524 0 1 1088
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_2143
timestamp 1676037725
transform 1 0 198260 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2155
timestamp 1676037725
transform 1 0 199364 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2157
timestamp 1676037725
transform 1 0 199548 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2163
timestamp 1676037725
transform 1 0 200100 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2171
timestamp 1676037725
transform 1 0 200836 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2180
timestamp 1676037725
transform 1 0 201664 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2185
timestamp 1676037725
transform 1 0 202124 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2192
timestamp 1676037725
transform 1 0 202768 0 1 1088
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_2200
timestamp 1676037725
transform 1 0 203504 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2213
timestamp 1676037725
transform 1 0 204700 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2221
timestamp 1676037725
transform 1 0 205436 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2226
timestamp 1676037725
transform 1 0 205896 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2230
timestamp 1676037725
transform 1 0 206264 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2234
timestamp 1676037725
transform 1 0 206632 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2241
timestamp 1676037725
transform 1 0 207276 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2246
timestamp 1676037725
transform 1 0 207736 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2253
timestamp 1676037725
transform 1 0 208380 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2260
timestamp 1676037725
transform 1 0 209024 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2269
timestamp 1676037725
transform 1 0 209852 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2274
timestamp 1676037725
transform 1 0 210312 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2281
timestamp 1676037725
transform 1 0 210956 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2288
timestamp 1676037725
transform 1 0 211600 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2297
timestamp 1676037725
transform 1 0 212428 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2302
timestamp 1676037725
transform 1 0 212888 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2309
timestamp 1676037725
transform 1 0 213532 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2316
timestamp 1676037725
transform 1 0 214176 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2325
timestamp 1676037725
transform 1 0 215004 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2330
timestamp 1676037725
transform 1 0 215464 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2337
timestamp 1676037725
transform 1 0 216108 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2344
timestamp 1676037725
transform 1 0 216752 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2353
timestamp 1676037725
transform 1 0 217580 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2361
timestamp 1676037725
transform 1 0 218316 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2371
timestamp 1676037725
transform 1 0 219236 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2378
timestamp 1676037725
transform 1 0 219880 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2381
timestamp 1676037725
transform 1 0 220156 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2386
timestamp 1676037725
transform 1 0 220616 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2393
timestamp 1676037725
transform 1 0 221260 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2400
timestamp 1676037725
transform 1 0 221904 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2409
timestamp 1676037725
transform 1 0 222732 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2414
timestamp 1676037725
transform 1 0 223192 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2426
timestamp 1676037725
transform 1 0 224296 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_2433
timestamp 1676037725
transform 1 0 224940 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2437
timestamp 1676037725
transform 1 0 225308 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2444
timestamp 1676037725
transform 1 0 225952 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2455
timestamp 1676037725
transform 1 0 226964 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2463
timestamp 1676037725
transform 1 0 227700 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2465
timestamp 1676037725
transform 1 0 227884 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2472
timestamp 1676037725
transform 1 0 228528 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2480
timestamp 1676037725
transform 1 0 229264 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2488
timestamp 1676037725
transform 1 0 230000 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2493
timestamp 1676037725
transform 1 0 230460 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_2499
timestamp 1676037725
transform 1 0 231012 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2516
timestamp 1676037725
transform 1 0 232576 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2521
timestamp 1676037725
transform 1 0 233036 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2527
timestamp 1676037725
transform 1 0 233588 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2535
timestamp 1676037725
transform 1 0 234324 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2543
timestamp 1676037725
transform 1 0 235060 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2547
timestamp 1676037725
transform 1 0 235428 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2549
timestamp 1676037725
transform 1 0 235612 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_2556
timestamp 1676037725
transform 1 0 236256 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2568
timestamp 1676037725
transform 1 0 237360 0 1 1088
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_2577
timestamp 1676037725
transform 1 0 238188 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2589
timestamp 1676037725
transform 1 0 239292 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2593
timestamp 1676037725
transform 1 0 239660 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2597
timestamp 1676037725
transform 1 0 240028 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2603
timestamp 1676037725
transform 1 0 240580 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2605
timestamp 1676037725
transform 1 0 240764 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_2617
timestamp 1676037725
transform 1 0 241868 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_2629
timestamp 1676037725
transform 1 0 242972 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2633
timestamp 1676037725
transform 1 0 243340 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_2645
timestamp 1676037725
transform 1 0 244444 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_2657
timestamp 1676037725
transform 1 0 245548 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2661
timestamp 1676037725
transform 1 0 245916 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2673
timestamp 1676037725
transform 1 0 247020 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2681
timestamp 1676037725
transform 1 0 247756 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2686
timestamp 1676037725
transform 1 0 248216 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2689
timestamp 1676037725
transform 1 0 248492 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2701
timestamp 1676037725
transform 1 0 249596 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2705
timestamp 1676037725
transform 1 0 249964 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2710
timestamp 1676037725
transform 1 0 250424 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2717
timestamp 1676037725
transform 1 0 251068 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2721
timestamp 1676037725
transform 1 0 251436 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_2732
timestamp 1676037725
transform 1 0 252448 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2745
timestamp 1676037725
transform 1 0 253644 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_2757
timestamp 1676037725
transform 1 0 254748 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_2769
timestamp 1676037725
transform 1 0 255852 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2773
timestamp 1676037725
transform 1 0 256220 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2785
timestamp 1676037725
transform 1 0 257324 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2794
timestamp 1676037725
transform 1 0 258152 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2801
timestamp 1676037725
transform 1 0 258796 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2813
timestamp 1676037725
transform 1 0 259900 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2821
timestamp 1676037725
transform 1 0 260636 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2827
timestamp 1676037725
transform 1 0 261188 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2829
timestamp 1676037725
transform 1 0 261372 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2835
timestamp 1676037725
transform 1 0 261924 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2843
timestamp 1676037725
transform 1 0 262660 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2851
timestamp 1676037725
transform 1 0 263396 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2855
timestamp 1676037725
transform 1 0 263764 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2857
timestamp 1676037725
transform 1 0 263948 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_2863
timestamp 1676037725
transform 1 0 264500 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2869
timestamp 1676037725
transform 1 0 265052 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2874
timestamp 1676037725
transform 1 0 265512 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2882
timestamp 1676037725
transform 1 0 266248 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2885
timestamp 1676037725
transform 1 0 266524 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2891
timestamp 1676037725
transform 1 0 267076 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2899
timestamp 1676037725
transform 1 0 267812 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2907
timestamp 1676037725
transform 1 0 268548 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_2911
timestamp 1676037725
transform 1 0 268916 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_2913
timestamp 1676037725
transform 1 0 269100 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_2920
timestamp 1676037725
transform 1 0 269744 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_2928
timestamp 1676037725
transform 1 0 270480 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_11
timestamp 1676037725
transform 1 0 2116 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_23
timestamp 1676037725
transform 1 0 3220 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_35
timestamp 1676037725
transform 1 0 4324 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_47
timestamp 1676037725
transform 1 0 5428 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_65
timestamp 1676037725
transform 1 0 7084 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_73
timestamp 1676037725
transform 1 0 7820 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_89
timestamp 1676037725
transform 1 0 9292 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_101
timestamp 1676037725
transform 1 0 10396 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_109
timestamp 1676037725
transform 1 0 11132 0 -1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_151
timestamp 1676037725
transform 1 0 14996 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_175
timestamp 1676037725
transform 1 0 17204 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_187
timestamp 1676037725
transform 1 0 18308 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_199
timestamp 1676037725
transform 1 0 19412 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_211
timestamp 1676037725
transform 1 0 20516 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_248
timestamp 1676037725
transform 1 0 23920 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_257
timestamp 1676037725
transform 1 0 24748 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_267
timestamp 1676037725
transform 1 0 25668 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_271
timestamp 1676037725
transform 1 0 26036 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_278
timestamp 1676037725
transform 1 0 26680 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_289
timestamp 1676037725
transform 1 0 27692 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_297
timestamp 1676037725
transform 1 0 28428 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_304
timestamp 1676037725
transform 1 0 29072 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_313
timestamp 1676037725
transform 1 0 29900 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_317
timestamp 1676037725
transform 1 0 30268 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_323
timestamp 1676037725
transform 1 0 30820 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_334
timestamp 1676037725
transform 1 0 31832 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_344
timestamp 1676037725
transform 1 0 32752 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_352
timestamp 1676037725
transform 1 0 33488 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_364
timestamp 1676037725
transform 1 0 34592 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_390
timestamp 1676037725
transform 1 0 36984 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_399
timestamp 1676037725
transform 1 0 37812 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_403
timestamp 1676037725
transform 1 0 38180 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_409
timestamp 1676037725
transform 1 0 38732 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_428
timestamp 1676037725
transform 1 0 40480 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_440
timestamp 1676037725
transform 1 0 41584 0 -1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_461
timestamp 1676037725
transform 1 0 43516 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_473
timestamp 1676037725
transform 1 0 44620 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_479
timestamp 1676037725
transform 1 0 45172 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_483
timestamp 1676037725
transform 1 0 45540 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_495
timestamp 1676037725
transform 1 0 46644 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_503
timestamp 1676037725
transform 1 0 47380 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_517
timestamp 1676037725
transform 1 0 48668 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_529
timestamp 1676037725
transform 1 0 49772 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_535
timestamp 1676037725
transform 1 0 50324 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_539
timestamp 1676037725
transform 1 0 50692 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_551
timestamp 1676037725
transform 1 0 51796 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_559
timestamp 1676037725
transform 1 0 52532 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_561
timestamp 1676037725
transform 1 0 52716 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_567
timestamp 1676037725
transform 1 0 53268 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_571
timestamp 1676037725
transform 1 0 53636 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_578
timestamp 1676037725
transform 1 0 54280 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_587
timestamp 1676037725
transform 1 0 55108 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_596
timestamp 1676037725
transform 1 0 55936 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_605
timestamp 1676037725
transform 1 0 56764 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_614
timestamp 1676037725
transform 1 0 57592 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_622
timestamp 1676037725
transform 1 0 58328 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_626
timestamp 1676037725
transform 1 0 58696 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_633
timestamp 1676037725
transform 1 0 59340 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_637
timestamp 1676037725
transform 1 0 59708 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_643
timestamp 1676037725
transform 1 0 60260 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_652
timestamp 1676037725
transform 1 0 61088 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_661
timestamp 1676037725
transform 1 0 61916 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_670
timestamp 1676037725
transform 1 0 62744 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_673
timestamp 1676037725
transform 1 0 63020 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_680
timestamp 1676037725
transform 1 0 63664 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_689
timestamp 1676037725
transform 1 0 64492 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_698
timestamp 1676037725
transform 1 0 65320 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_707
timestamp 1676037725
transform 1 0 66148 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_716
timestamp 1676037725
transform 1 0 66976 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_724
timestamp 1676037725
transform 1 0 67712 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_729
timestamp 1676037725
transform 1 0 68172 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_741
timestamp 1676037725
transform 1 0 69276 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_753
timestamp 1676037725
transform 1 0 70380 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_765
timestamp 1676037725
transform 1 0 71484 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_781
timestamp 1676037725
transform 1 0 72956 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_785
timestamp 1676037725
transform 1 0 73324 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_793
timestamp 1676037725
transform 1 0 74060 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_805
timestamp 1676037725
transform 1 0 75164 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_821
timestamp 1676037725
transform 1 0 76636 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_837
timestamp 1676037725
transform 1 0 78108 0 -1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_841
timestamp 1676037725
transform 1 0 78476 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_853
timestamp 1676037725
transform 1 0 79580 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_866
timestamp 1676037725
transform 1 0 80776 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_880
timestamp 1676037725
transform 1 0 82064 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_894
timestamp 1676037725
transform 1 0 83352 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_897
timestamp 1676037725
transform 1 0 83628 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_920
timestamp 1676037725
transform 1 0 85744 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_934
timestamp 1676037725
transform 1 0 87032 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_940
timestamp 1676037725
transform 1 0 87584 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_943
timestamp 1676037725
transform 1 0 87860 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_950
timestamp 1676037725
transform 1 0 88504 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_953
timestamp 1676037725
transform 1 0 88780 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_961
timestamp 1676037725
transform 1 0 89516 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_970
timestamp 1676037725
transform 1 0 90344 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_979
timestamp 1676037725
transform 1 0 91172 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_988
timestamp 1676037725
transform 1 0 92000 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_997
timestamp 1676037725
transform 1 0 92828 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1006
timestamp 1676037725
transform 1 0 93656 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1009
timestamp 1676037725
transform 1 0 93932 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1016
timestamp 1676037725
transform 1 0 94576 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1020
timestamp 1676037725
transform 1 0 94944 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1026
timestamp 1676037725
transform 1 0 95496 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1035
timestamp 1676037725
transform 1 0 96324 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1044
timestamp 1676037725
transform 1 0 97152 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1053
timestamp 1676037725
transform 1 0 97980 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1062
timestamp 1676037725
transform 1 0 98808 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_1065
timestamp 1676037725
transform 1 0 99084 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1074
timestamp 1676037725
transform 1 0 99912 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1083
timestamp 1676037725
transform 1 0 100740 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1091
timestamp 1676037725
transform 1 0 101476 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1099
timestamp 1676037725
transform 1 0 102212 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_1111
timestamp 1676037725
transform 1 0 103316 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1119
timestamp 1676037725
transform 1 0 104052 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1121
timestamp 1676037725
transform 1 0 104236 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1133
timestamp 1676037725
transform 1 0 105340 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1145
timestamp 1676037725
transform 1 0 106444 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1149
timestamp 1676037725
transform 1 0 106812 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1153
timestamp 1676037725
transform 1 0 107180 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_1165
timestamp 1676037725
transform 1 0 108284 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_1173
timestamp 1676037725
transform 1 0 109020 0 -1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1177
timestamp 1676037725
transform 1 0 109388 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1189
timestamp 1676037725
transform 1 0 110492 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1201
timestamp 1676037725
transform 1 0 111596 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1205
timestamp 1676037725
transform 1 0 111964 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1209
timestamp 1676037725
transform 1 0 112332 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_1221
timestamp 1676037725
transform 1 0 113436 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_1229
timestamp 1676037725
transform 1 0 114172 0 -1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1233
timestamp 1676037725
transform 1 0 114540 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1245
timestamp 1676037725
transform 1 0 115644 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1257
timestamp 1676037725
transform 1 0 116748 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1261
timestamp 1676037725
transform 1 0 117116 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1265
timestamp 1676037725
transform 1 0 117484 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_1277
timestamp 1676037725
transform 1 0 118588 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_1285
timestamp 1676037725
transform 1 0 119324 0 -1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1289
timestamp 1676037725
transform 1 0 119692 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1306
timestamp 1676037725
transform 1 0 121256 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1315
timestamp 1676037725
transform 1 0 122084 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1324
timestamp 1676037725
transform 1 0 122912 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1333
timestamp 1676037725
transform 1 0 123740 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1342
timestamp 1676037725
transform 1 0 124568 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1345
timestamp 1676037725
transform 1 0 124844 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1352
timestamp 1676037725
transform 1 0 125488 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1361
timestamp 1676037725
transform 1 0 126316 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1370
timestamp 1676037725
transform 1 0 127144 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1379
timestamp 1676037725
transform 1 0 127972 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1383
timestamp 1676037725
transform 1 0 128340 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1389
timestamp 1676037725
transform 1 0 128892 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1398
timestamp 1676037725
transform 1 0 129720 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1401
timestamp 1676037725
transform 1 0 129996 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1405
timestamp 1676037725
transform 1 0 130364 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1411
timestamp 1676037725
transform 1 0 130916 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1420
timestamp 1676037725
transform 1 0 131744 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1424
timestamp 1676037725
transform 1 0 132112 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_1430
timestamp 1676037725
transform 1 0 132664 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1441
timestamp 1676037725
transform 1 0 133676 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_1450
timestamp 1676037725
transform 1 0 134504 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1457
timestamp 1676037725
transform 1 0 135148 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1463
timestamp 1676037725
transform 1 0 135700 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1475
timestamp 1676037725
transform 1 0 136804 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1487
timestamp 1676037725
transform 1 0 137908 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1510
timestamp 1676037725
transform 1 0 140024 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1513
timestamp 1676037725
transform 1 0 140300 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1536
timestamp 1676037725
transform 1 0 142416 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1543
timestamp 1676037725
transform 1 0 143060 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_1555
timestamp 1676037725
transform 1 0 144164 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1564
timestamp 1676037725
transform 1 0 144992 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1569
timestamp 1676037725
transform 1 0 145452 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1581
timestamp 1676037725
transform 1 0 146556 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1593
timestamp 1676037725
transform 1 0 147660 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1605
timestamp 1676037725
transform 1 0 148764 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1620
timestamp 1676037725
transform 1 0 150144 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1625
timestamp 1676037725
transform 1 0 150604 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1637
timestamp 1676037725
transform 1 0 151708 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1649
timestamp 1676037725
transform 1 0 152812 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1661
timestamp 1676037725
transform 1 0 153916 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1673
timestamp 1676037725
transform 1 0 155020 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1678
timestamp 1676037725
transform 1 0 155480 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1681
timestamp 1676037725
transform 1 0 155756 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1687
timestamp 1676037725
transform 1 0 156308 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1700
timestamp 1676037725
transform 1 0 157504 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1713
timestamp 1676037725
transform 1 0 158700 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1722
timestamp 1676037725
transform 1 0 159528 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1731
timestamp 1676037725
transform 1 0 160356 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1735
timestamp 1676037725
transform 1 0 160724 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1737
timestamp 1676037725
transform 1 0 160908 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1744
timestamp 1676037725
transform 1 0 161552 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1753
timestamp 1676037725
transform 1 0 162380 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1762
timestamp 1676037725
transform 1 0 163208 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1771
timestamp 1676037725
transform 1 0 164036 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1780
timestamp 1676037725
transform 1 0 164864 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_1789
timestamp 1676037725
transform 1 0 165692 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1793
timestamp 1676037725
transform 1 0 166060 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1800
timestamp 1676037725
transform 1 0 166704 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1809
timestamp 1676037725
transform 1 0 167532 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1818
timestamp 1676037725
transform 1 0 168360 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1826
timestamp 1676037725
transform 1 0 169096 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_1838
timestamp 1676037725
transform 1 0 170200 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1846
timestamp 1676037725
transform 1 0 170936 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1849
timestamp 1676037725
transform 1 0 171212 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_1861
timestamp 1676037725
transform 1 0 172316 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_1867
timestamp 1676037725
transform 1 0 172868 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_1878
timestamp 1676037725
transform 1 0 173880 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_1894
timestamp 1676037725
transform 1 0 175352 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1902
timestamp 1676037725
transform 1 0 176088 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_1905
timestamp 1676037725
transform 1 0 176364 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1917
timestamp 1676037725
transform 1 0 177468 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_1931
timestamp 1676037725
transform 1 0 178756 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1945
timestamp 1676037725
transform 1 0 180044 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_1957
timestamp 1676037725
transform 1 0 181148 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_1961
timestamp 1676037725
transform 1 0 181516 0 -1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_1968
timestamp 1676037725
transform 1 0 182160 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_1990
timestamp 1676037725
transform 1 0 184184 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_2006
timestamp 1676037725
transform 1 0 185656 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2014
timestamp 1676037725
transform 1 0 186392 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2017
timestamp 1676037725
transform 1 0 186668 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2029
timestamp 1676037725
transform 1 0 187772 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2043
timestamp 1676037725
transform 1 0 189060 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2057
timestamp 1676037725
transform 1 0 190348 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_2066
timestamp 1676037725
transform 1 0 191176 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2073
timestamp 1676037725
transform 1 0 191820 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2080
timestamp 1676037725
transform 1 0 192464 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2089
timestamp 1676037725
transform 1 0 193292 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2098
timestamp 1676037725
transform 1 0 194120 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2107
timestamp 1676037725
transform 1 0 194948 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2116
timestamp 1676037725
transform 1 0 195776 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_2125
timestamp 1676037725
transform 1 0 196604 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2129
timestamp 1676037725
transform 1 0 196972 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2136
timestamp 1676037725
transform 1 0 197616 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2145
timestamp 1676037725
transform 1 0 198444 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2154
timestamp 1676037725
transform 1 0 199272 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2163
timestamp 1676037725
transform 1 0 200100 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2172
timestamp 1676037725
transform 1 0 200928 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_2181
timestamp 1676037725
transform 1 0 201756 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2185
timestamp 1676037725
transform 1 0 202124 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2192
timestamp 1676037725
transform 1 0 202768 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_2200
timestamp 1676037725
transform 1 0 203504 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_2212
timestamp 1676037725
transform 1 0 204608 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_2224
timestamp 1676037725
transform 1 0 205712 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2236
timestamp 1676037725
transform 1 0 206816 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_2241
timestamp 1676037725
transform 1 0 207276 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_2253
timestamp 1676037725
transform 1 0 208380 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_2265
timestamp 1676037725
transform 1 0 209484 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_2277
timestamp 1676037725
transform 1 0 210588 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2285
timestamp 1676037725
transform 1 0 211324 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_2290
timestamp 1676037725
transform 1 0 211784 0 -1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_2297
timestamp 1676037725
transform 1 0 212428 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_2309
timestamp 1676037725
transform 1 0 213532 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_2321
timestamp 1676037725
transform 1 0 214636 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2333
timestamp 1676037725
transform 1 0 215740 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2346
timestamp 1676037725
transform 1 0 216936 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2350
timestamp 1676037725
transform 1 0 217304 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2353
timestamp 1676037725
transform 1 0 217580 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2363
timestamp 1676037725
transform 1 0 218500 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2373
timestamp 1676037725
transform 1 0 219420 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2383
timestamp 1676037725
transform 1 0 220340 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2393
timestamp 1676037725
transform 1 0 221260 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_2400
timestamp 1676037725
transform 1 0 221904 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2409
timestamp 1676037725
transform 1 0 222732 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2417
timestamp 1676037725
transform 1 0 223468 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_2427
timestamp 1676037725
transform 1 0 224388 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2438
timestamp 1676037725
transform 1 0 225400 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2447
timestamp 1676037725
transform 1 0 226228 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_2456
timestamp 1676037725
transform 1 0 227056 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2465
timestamp 1676037725
transform 1 0 227884 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2472
timestamp 1676037725
transform 1 0 228528 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2481
timestamp 1676037725
transform 1 0 229356 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2490
timestamp 1676037725
transform 1 0 230184 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2499
timestamp 1676037725
transform 1 0 231012 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2508
timestamp 1676037725
transform 1 0 231840 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_2517
timestamp 1676037725
transform 1 0 232668 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2521
timestamp 1676037725
transform 1 0 233036 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2528
timestamp 1676037725
transform 1 0 233680 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2537
timestamp 1676037725
transform 1 0 234508 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2546
timestamp 1676037725
transform 1 0 235336 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2555
timestamp 1676037725
transform 1 0 236164 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2564
timestamp 1676037725
transform 1 0 236992 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2572
timestamp 1676037725
transform 1 0 237728 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_2577
timestamp 1676037725
transform 1 0 238188 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_2589
timestamp 1676037725
transform 1 0 239292 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_2601
timestamp 1676037725
transform 1 0 240396 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_2609
timestamp 1676037725
transform 1 0 241132 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_2620
timestamp 1676037725
transform 1 0 242144 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2633
timestamp 1676037725
transform 1 0 243340 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2645
timestamp 1676037725
transform 1 0 244444 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2659
timestamp 1676037725
transform 1 0 245732 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_2673
timestamp 1676037725
transform 1 0 247020 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_2685
timestamp 1676037725
transform 1 0 248124 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2689
timestamp 1676037725
transform 1 0 248492 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2701
timestamp 1676037725
transform 1 0 249596 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2715
timestamp 1676037725
transform 1 0 250884 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_2723
timestamp 1676037725
transform 1 0 251620 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_2729
timestamp 1676037725
transform 1 0 252172 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2740
timestamp 1676037725
transform 1 0 253184 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2745
timestamp 1676037725
transform 1 0 253644 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2757
timestamp 1676037725
transform 1 0 254748 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2771
timestamp 1676037725
transform 1 0 256036 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2785
timestamp 1676037725
transform 1 0 257324 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_2789
timestamp 1676037725
transform 1 0 257692 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2796
timestamp 1676037725
transform 1 0 258336 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2801
timestamp 1676037725
transform 1 0 258796 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2808
timestamp 1676037725
transform 1 0 259440 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2817
timestamp 1676037725
transform 1 0 260268 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2826
timestamp 1676037725
transform 1 0 261096 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2835
timestamp 1676037725
transform 1 0 261924 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2844
timestamp 1676037725
transform 1 0 262752 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_2853
timestamp 1676037725
transform 1 0 263580 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2857
timestamp 1676037725
transform 1 0 263948 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2864
timestamp 1676037725
transform 1 0 264592 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2873
timestamp 1676037725
transform 1 0 265420 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2882
timestamp 1676037725
transform 1 0 266248 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2891
timestamp 1676037725
transform 1 0 267076 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2900
timestamp 1676037725
transform 1 0 267904 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_2909
timestamp 1676037725
transform 1 0 268732 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_2913
timestamp 1676037725
transform 1 0 269100 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_2920
timestamp 1676037725
transform 1 0 269744 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_2929
timestamp 1676037725
transform 1 0 270572 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_2935
timestamp 1676037725
transform 1 0 271124 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_3
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1676037725
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1676037725
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1676037725
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1676037725
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1676037725
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1676037725
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1676037725
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1676037725
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1676037725
transform 1 0 17388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1676037725
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1676037725
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1676037725
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1676037725
transform 1 0 21436 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1676037725
transform 1 0 22540 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_245
timestamp 1676037725
transform 1 0 23644 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_263
timestamp 1676037725
transform 1 0 25300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_267
timestamp 1676037725
transform 1 0 25668 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_274
timestamp 1676037725
transform 1 0 26312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_283
timestamp 1676037725
transform 1 0 27140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_287
timestamp 1676037725
transform 1 0 27508 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_294
timestamp 1676037725
transform 1 0 28152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_302
timestamp 1676037725
transform 1 0 28888 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_333
timestamp 1676037725
transform 1 0 31740 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_343
timestamp 1676037725
transform 1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_350
timestamp 1676037725
transform 1 0 33304 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_362
timestamp 1676037725
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_377
timestamp 1676037725
transform 1 0 35788 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_385
timestamp 1676037725
transform 1 0 36524 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_405
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_417
timestamp 1676037725
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1676037725
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_445
timestamp 1676037725
transform 1 0 42044 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_457
timestamp 1676037725
transform 1 0 43148 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_469
timestamp 1676037725
transform 1 0 44252 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_475
timestamp 1676037725
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_489
timestamp 1676037725
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_501
timestamp 1676037725
transform 1 0 47196 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_513
timestamp 1676037725
transform 1 0 48300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_525
timestamp 1676037725
transform 1 0 49404 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_531
timestamp 1676037725
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_533
timestamp 1676037725
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_545
timestamp 1676037725
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_557
timestamp 1676037725
transform 1 0 52348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_569
timestamp 1676037725
transform 1 0 53452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_577
timestamp 1676037725
transform 1 0 54188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_581
timestamp 1676037725
transform 1 0 54556 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_586
timestamp 1676037725
transform 1 0 55016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_589
timestamp 1676037725
transform 1 0 55292 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_595
timestamp 1676037725
transform 1 0 55844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_607
timestamp 1676037725
transform 1 0 56948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_613
timestamp 1676037725
transform 1 0 57500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_618
timestamp 1676037725
transform 1 0 57960 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_626
timestamp 1676037725
transform 1 0 58696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_630
timestamp 1676037725
transform 1 0 59064 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_635
timestamp 1676037725
transform 1 0 59524 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_643
timestamp 1676037725
transform 1 0 60260 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_645
timestamp 1676037725
transform 1 0 60444 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_651
timestamp 1676037725
transform 1 0 60996 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_663
timestamp 1676037725
transform 1 0 62100 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_669
timestamp 1676037725
transform 1 0 62652 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_674
timestamp 1676037725
transform 1 0 63112 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_686
timestamp 1676037725
transform 1 0 64216 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_698
timestamp 1676037725
transform 1 0 65320 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_701
timestamp 1676037725
transform 1 0 65596 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_707
timestamp 1676037725
transform 1 0 66148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_711
timestamp 1676037725
transform 1 0 66516 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_715
timestamp 1676037725
transform 1 0 66884 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_727
timestamp 1676037725
transform 1 0 67988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_739
timestamp 1676037725
transform 1 0 69092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_751
timestamp 1676037725
transform 1 0 70196 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_755
timestamp 1676037725
transform 1 0 70564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_757
timestamp 1676037725
transform 1 0 70748 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_773
timestamp 1676037725
transform 1 0 72220 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_785
timestamp 1676037725
transform 1 0 73324 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_797
timestamp 1676037725
transform 1 0 74428 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_809
timestamp 1676037725
transform 1 0 75532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_813
timestamp 1676037725
transform 1 0 75900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_829
timestamp 1676037725
transform 1 0 77372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_845
timestamp 1676037725
transform 1 0 78844 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_861
timestamp 1676037725
transform 1 0 80316 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_867
timestamp 1676037725
transform 1 0 80868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_869
timestamp 1676037725
transform 1 0 81052 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_877
timestamp 1676037725
transform 1 0 81788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_890
timestamp 1676037725
transform 1 0 82984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_894
timestamp 1676037725
transform 1 0 83352 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_917
timestamp 1676037725
transform 1 0 85468 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_921
timestamp 1676037725
transform 1 0 85836 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_925
timestamp 1676037725
transform 1 0 86204 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_937
timestamp 1676037725
transform 1 0 87308 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_942
timestamp 1676037725
transform 1 0 87768 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_946
timestamp 1676037725
transform 1 0 88136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_969
timestamp 1676037725
transform 1 0 90252 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_977
timestamp 1676037725
transform 1 0 90988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_981
timestamp 1676037725
transform 1 0 91356 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_987
timestamp 1676037725
transform 1 0 91908 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_995
timestamp 1676037725
transform 1 0 92644 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1001
timestamp 1676037725
transform 1 0 93196 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1005
timestamp 1676037725
transform 1 0 93564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1010
timestamp 1676037725
transform 1 0 94024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1018
timestamp 1676037725
transform 1 0 94760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1026
timestamp 1676037725
transform 1 0 95496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1034
timestamp 1676037725
transform 1 0 96232 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1037
timestamp 1676037725
transform 1 0 96508 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1060
timestamp 1676037725
transform 1 0 98624 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1066
timestamp 1676037725
transform 1 0 99176 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_1089
timestamp 1676037725
transform 1 0 101292 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1093
timestamp 1676037725
transform 1 0 101660 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1105
timestamp 1676037725
transform 1 0 102764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1111
timestamp 1676037725
transform 1 0 103316 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1133
timestamp 1676037725
transform 1 0 105340 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_1145
timestamp 1676037725
transform 1 0 106444 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1149
timestamp 1676037725
transform 1 0 106812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1161
timestamp 1676037725
transform 1 0 107916 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1188
timestamp 1676037725
transform 1 0 110400 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1200
timestamp 1676037725
transform 1 0 111504 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1205
timestamp 1676037725
transform 1 0 111964 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1217
timestamp 1676037725
transform 1 0 113068 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1229
timestamp 1676037725
transform 1 0 114172 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1241
timestamp 1676037725
transform 1 0 115276 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1253
timestamp 1676037725
transform 1 0 116380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1259
timestamp 1676037725
transform 1 0 116932 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1261
timestamp 1676037725
transform 1 0 117116 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1273
timestamp 1676037725
transform 1 0 118220 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1285
timestamp 1676037725
transform 1 0 119324 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1297
timestamp 1676037725
transform 1 0 120428 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1309
timestamp 1676037725
transform 1 0 121532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1315
timestamp 1676037725
transform 1 0 122084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1317
timestamp 1676037725
transform 1 0 122268 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1323
timestamp 1676037725
transform 1 0 122820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1335
timestamp 1676037725
transform 1 0 123924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1341
timestamp 1676037725
transform 1 0 124476 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1346
timestamp 1676037725
transform 1 0 124936 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1358
timestamp 1676037725
transform 1 0 126040 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_1363
timestamp 1676037725
transform 1 0 126500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1371
timestamp 1676037725
transform 1 0 127236 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1373
timestamp 1676037725
transform 1 0 127420 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1379
timestamp 1676037725
transform 1 0 127972 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1387
timestamp 1676037725
transform 1 0 128708 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1403
timestamp 1676037725
transform 1 0 130180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1415
timestamp 1676037725
transform 1 0 131284 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_1420
timestamp 1676037725
transform 1 0 131744 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1429
timestamp 1676037725
transform 1 0 132572 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1435
timestamp 1676037725
transform 1 0 133124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1443
timestamp 1676037725
transform 1 0 133860 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1451
timestamp 1676037725
transform 1 0 134596 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1458
timestamp 1676037725
transform 1 0 135240 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1470
timestamp 1676037725
transform 1 0 136344 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1482
timestamp 1676037725
transform 1 0 137448 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_1485
timestamp 1676037725
transform 1 0 137724 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1493
timestamp 1676037725
transform 1 0 138460 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1496
timestamp 1676037725
transform 1 0 138736 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1519
timestamp 1676037725
transform 1 0 140852 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1523
timestamp 1676037725
transform 1 0 141220 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1535
timestamp 1676037725
transform 1 0 142324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1539
timestamp 1676037725
transform 1 0 142692 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1541
timestamp 1676037725
transform 1 0 142876 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1564
timestamp 1676037725
transform 1 0 144992 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1576
timestamp 1676037725
transform 1 0 146096 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_1588
timestamp 1676037725
transform 1 0 147200 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1597
timestamp 1676037725
transform 1 0 148028 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1620
timestamp 1676037725
transform 1 0 150144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1645
timestamp 1676037725
transform 1 0 152444 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1651
timestamp 1676037725
transform 1 0 152996 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1653
timestamp 1676037725
transform 1 0 153180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_1665
timestamp 1676037725
transform 1 0 154284 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1676
timestamp 1676037725
transform 1 0 155296 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1688
timestamp 1676037725
transform 1 0 156400 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1706
timestamp 1676037725
transform 1 0 158056 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1709
timestamp 1676037725
transform 1 0 158332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1720
timestamp 1676037725
transform 1 0 159344 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1739
timestamp 1676037725
transform 1 0 161092 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1743
timestamp 1676037725
transform 1 0 161460 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1748
timestamp 1676037725
transform 1 0 161920 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1760
timestamp 1676037725
transform 1 0 163024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1765
timestamp 1676037725
transform 1 0 163484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1771
timestamp 1676037725
transform 1 0 164036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1779
timestamp 1676037725
transform 1 0 164772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1787
timestamp 1676037725
transform 1 0 165508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1795
timestamp 1676037725
transform 1 0 166244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1803
timestamp 1676037725
transform 1 0 166980 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1809
timestamp 1676037725
transform 1 0 167532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_1815
timestamp 1676037725
transform 1 0 168084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1819
timestamp 1676037725
transform 1 0 168452 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1821
timestamp 1676037725
transform 1 0 168636 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1833
timestamp 1676037725
transform 1 0 169740 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1845
timestamp 1676037725
transform 1 0 170844 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1857
timestamp 1676037725
transform 1 0 171948 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1869
timestamp 1676037725
transform 1 0 173052 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1875
timestamp 1676037725
transform 1 0 173604 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1877
timestamp 1676037725
transform 1 0 173788 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1889
timestamp 1676037725
transform 1 0 174892 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1901
timestamp 1676037725
transform 1 0 175996 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1907
timestamp 1676037725
transform 1 0 176548 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1918
timestamp 1676037725
transform 1 0 177560 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1930
timestamp 1676037725
transform 1 0 178664 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_1933
timestamp 1676037725
transform 1 0 178940 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_1939
timestamp 1676037725
transform 1 0 179492 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1950
timestamp 1676037725
transform 1 0 180504 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1962
timestamp 1676037725
transform 1 0 181608 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1974
timestamp 1676037725
transform 1 0 182712 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_1986
timestamp 1676037725
transform 1 0 183816 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_1989
timestamp 1676037725
transform 1 0 184092 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2001
timestamp 1676037725
transform 1 0 185196 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_2013
timestamp 1676037725
transform 1 0 186300 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2019
timestamp 1676037725
transform 1 0 186852 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2030
timestamp 1676037725
transform 1 0 187864 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2042
timestamp 1676037725
transform 1 0 188968 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2045
timestamp 1676037725
transform 1 0 189244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2061
timestamp 1676037725
transform 1 0 190716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2069
timestamp 1676037725
transform 1 0 191452 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2077
timestamp 1676037725
transform 1 0 192188 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_2089
timestamp 1676037725
transform 1 0 193292 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_2097
timestamp 1676037725
transform 1 0 194028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2101
timestamp 1676037725
transform 1 0 194396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2105
timestamp 1676037725
transform 1 0 194764 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_2110
timestamp 1676037725
transform 1 0 195224 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_2118
timestamp 1676037725
transform 1 0 195960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2125
timestamp 1676037725
transform 1 0 196604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2129
timestamp 1676037725
transform 1 0 196972 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_2135
timestamp 1676037725
transform 1 0 197524 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2143
timestamp 1676037725
transform 1 0 198260 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_2148
timestamp 1676037725
transform 1 0 198720 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2157
timestamp 1676037725
transform 1 0 199548 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2163
timestamp 1676037725
transform 1 0 200100 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2179
timestamp 1676037725
transform 1 0 201572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2188
timestamp 1676037725
transform 1 0 202400 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2196
timestamp 1676037725
transform 1 0 203136 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2210
timestamp 1676037725
transform 1 0 204424 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2213
timestamp 1676037725
transform 1 0 204700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2236
timestamp 1676037725
transform 1 0 206816 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2240
timestamp 1676037725
transform 1 0 207184 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2252
timestamp 1676037725
transform 1 0 208288 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2264
timestamp 1676037725
transform 1 0 209392 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2269
timestamp 1676037725
transform 1 0 209852 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2292
timestamp 1676037725
transform 1 0 211968 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2304
timestamp 1676037725
transform 1 0 213072 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_2316
timestamp 1676037725
transform 1 0 214176 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_2325
timestamp 1676037725
transform 1 0 215004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_2333
timestamp 1676037725
transform 1 0 215740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2344
timestamp 1676037725
transform 1 0 216752 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2348
timestamp 1676037725
transform 1 0 217120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2358
timestamp 1676037725
transform 1 0 218040 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2362
timestamp 1676037725
transform 1 0 218408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2372
timestamp 1676037725
transform 1 0 219328 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2376
timestamp 1676037725
transform 1 0 219696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_2381
timestamp 1676037725
transform 1 0 220156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2386
timestamp 1676037725
transform 1 0 220616 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2396
timestamp 1676037725
transform 1 0 221536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2408
timestamp 1676037725
transform 1 0 222640 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2420
timestamp 1676037725
transform 1 0 223744 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2426
timestamp 1676037725
transform 1 0 224296 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2430
timestamp 1676037725
transform 1 0 224664 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2434
timestamp 1676037725
transform 1 0 225032 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2445
timestamp 1676037725
transform 1 0 226044 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2451
timestamp 1676037725
transform 1 0 226596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_2459
timestamp 1676037725
transform 1 0 227332 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2471
timestamp 1676037725
transform 1 0 228436 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2479
timestamp 1676037725
transform 1 0 229172 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2491
timestamp 1676037725
transform 1 0 230276 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_2493
timestamp 1676037725
transform 1 0 230460 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2499
timestamp 1676037725
transform 1 0 231012 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2504
timestamp 1676037725
transform 1 0 231472 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2512
timestamp 1676037725
transform 1 0 232208 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2520
timestamp 1676037725
transform 1 0 232944 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2532
timestamp 1676037725
transform 1 0 234048 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2544
timestamp 1676037725
transform 1 0 235152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2549
timestamp 1676037725
transform 1 0 235612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2555
timestamp 1676037725
transform 1 0 236164 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2563
timestamp 1676037725
transform 1 0 236900 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2575
timestamp 1676037725
transform 1 0 238004 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2587
timestamp 1676037725
transform 1 0 239108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2599
timestamp 1676037725
transform 1 0 240212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2603
timestamp 1676037725
transform 1 0 240580 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2605
timestamp 1676037725
transform 1 0 240764 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2617
timestamp 1676037725
transform 1 0 241868 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2629
timestamp 1676037725
transform 1 0 242972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2633
timestamp 1676037725
transform 1 0 243340 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2644
timestamp 1676037725
transform 1 0 244352 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2656
timestamp 1676037725
transform 1 0 245456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2661
timestamp 1676037725
transform 1 0 245916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2665
timestamp 1676037725
transform 1 0 246284 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2676
timestamp 1676037725
transform 1 0 247296 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2688
timestamp 1676037725
transform 1 0 248400 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2700
timestamp 1676037725
transform 1 0 249504 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2712
timestamp 1676037725
transform 1 0 250608 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2717
timestamp 1676037725
transform 1 0 251068 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2729
timestamp 1676037725
transform 1 0 252172 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2741
timestamp 1676037725
transform 1 0 253276 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2753
timestamp 1676037725
transform 1 0 254380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_2765
timestamp 1676037725
transform 1 0 255484 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2771
timestamp 1676037725
transform 1 0 256036 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2773
timestamp 1676037725
transform 1 0 256220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2777
timestamp 1676037725
transform 1 0 256588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2788
timestamp 1676037725
transform 1 0 257600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2798
timestamp 1676037725
transform 1 0 258520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2807
timestamp 1676037725
transform 1 0 259348 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2815
timestamp 1676037725
transform 1 0 260084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2827
timestamp 1676037725
transform 1 0 261188 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2829
timestamp 1676037725
transform 1 0 261372 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_2835
timestamp 1676037725
transform 1 0 261924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_2847
timestamp 1676037725
transform 1 0 263028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2855
timestamp 1676037725
transform 1 0 263764 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2862
timestamp 1676037725
transform 1 0 264408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_2870
timestamp 1676037725
transform 1 0 265144 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_2878
timestamp 1676037725
transform 1 0 265880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_2882
timestamp 1676037725
transform 1 0 266248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_2885
timestamp 1676037725
transform 1 0 266524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2894
timestamp 1676037725
transform 1 0 267352 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2901
timestamp 1676037725
transform 1 0 267996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2908
timestamp 1676037725
transform 1 0 268640 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2917
timestamp 1676037725
transform 1 0 269468 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_2925
timestamp 1676037725
transform 1 0 270204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_2933
timestamp 1676037725
transform 1 0 270940 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_256
timestamp 1676037725
transform 1 0 24656 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_260
timestamp 1676037725
transform 1 0 25024 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_267
timestamp 1676037725
transform 1 0 25668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_276
timestamp 1676037725
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_290
timestamp 1676037725
transform 1 0 27784 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_296
timestamp 1676037725
transform 1 0 28336 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_308
timestamp 1676037725
transform 1 0 29440 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_320
timestamp 1676037725
transform 1 0 30544 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_332
timestamp 1676037725
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_415
timestamp 1676037725
transform 1 0 39284 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_437
timestamp 1676037725
transform 1 0 41308 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_445
timestamp 1676037725
transform 1 0 42044 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_461
timestamp 1676037725
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_473
timestamp 1676037725
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_485
timestamp 1676037725
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_497
timestamp 1676037725
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_503
timestamp 1676037725
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_517
timestamp 1676037725
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_529
timestamp 1676037725
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_541
timestamp 1676037725
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_553
timestamp 1676037725
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_559
timestamp 1676037725
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_561
timestamp 1676037725
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_573
timestamp 1676037725
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_585
timestamp 1676037725
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_597
timestamp 1676037725
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_609
timestamp 1676037725
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_615
timestamp 1676037725
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_617
timestamp 1676037725
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_629
timestamp 1676037725
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_641
timestamp 1676037725
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_653
timestamp 1676037725
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_665
timestamp 1676037725
transform 1 0 62284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_671
timestamp 1676037725
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_673
timestamp 1676037725
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_685
timestamp 1676037725
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_697
timestamp 1676037725
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_709
timestamp 1676037725
transform 1 0 66332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_721
timestamp 1676037725
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_727
timestamp 1676037725
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_729
timestamp 1676037725
transform 1 0 68172 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_741
timestamp 1676037725
transform 1 0 69276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_753
timestamp 1676037725
transform 1 0 70380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_765
timestamp 1676037725
transform 1 0 71484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_777
timestamp 1676037725
transform 1 0 72588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_783
timestamp 1676037725
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_785
timestamp 1676037725
transform 1 0 73324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_797
timestamp 1676037725
transform 1 0 74428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_809
timestamp 1676037725
transform 1 0 75532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_821
timestamp 1676037725
transform 1 0 76636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_833
timestamp 1676037725
transform 1 0 77740 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_839
timestamp 1676037725
transform 1 0 78292 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_841
timestamp 1676037725
transform 1 0 78476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_853
timestamp 1676037725
transform 1 0 79580 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_865
timestamp 1676037725
transform 1 0 80684 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_877
timestamp 1676037725
transform 1 0 81788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_890
timestamp 1676037725
transform 1 0 82984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_894
timestamp 1676037725
transform 1 0 83352 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_897
timestamp 1676037725
transform 1 0 83628 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_902
timestamp 1676037725
transform 1 0 84088 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_925
timestamp 1676037725
transform 1 0 86204 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_950
timestamp 1676037725
transform 1 0 88504 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_953
timestamp 1676037725
transform 1 0 88780 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_961
timestamp 1676037725
transform 1 0 89516 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_965
timestamp 1676037725
transform 1 0 89884 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_988
timestamp 1676037725
transform 1 0 92000 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_992
timestamp 1676037725
transform 1 0 92368 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1004
timestamp 1676037725
transform 1 0 93472 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_1009
timestamp 1676037725
transform 1 0 93932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1033
timestamp 1676037725
transform 1 0 96140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1039
timestamp 1676037725
transform 1 0 96692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1062
timestamp 1676037725
transform 1 0 98808 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_1065
timestamp 1676037725
transform 1 0 99084 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1092
timestamp 1676037725
transform 1 0 101568 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1114
timestamp 1676037725
transform 1 0 103592 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1118
timestamp 1676037725
transform 1 0 103960 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1121
timestamp 1676037725
transform 1 0 104236 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1144
timestamp 1676037725
transform 1 0 106352 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1148
timestamp 1676037725
transform 1 0 106720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_1173
timestamp 1676037725
transform 1 0 109020 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_1177
timestamp 1676037725
transform 1 0 109388 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1185
timestamp 1676037725
transform 1 0 110124 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1207
timestamp 1676037725
transform 1 0 112148 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1219
timestamp 1676037725
transform 1 0 113252 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1231
timestamp 1676037725
transform 1 0 114356 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1233
timestamp 1676037725
transform 1 0 114540 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1245
timestamp 1676037725
transform 1 0 115644 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1248
timestamp 1676037725
transform 1 0 115920 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1252
timestamp 1676037725
transform 1 0 116288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1275
timestamp 1676037725
transform 1 0 118404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_1279
timestamp 1676037725
transform 1 0 118772 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1287
timestamp 1676037725
transform 1 0 119508 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_1289
timestamp 1676037725
transform 1 0 119692 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1297
timestamp 1676037725
transform 1 0 120428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1301
timestamp 1676037725
transform 1 0 120796 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1305
timestamp 1676037725
transform 1 0 121164 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1328
timestamp 1676037725
transform 1 0 123280 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1332
timestamp 1676037725
transform 1 0 123648 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1345
timestamp 1676037725
transform 1 0 124844 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1357
timestamp 1676037725
transform 1 0 125948 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1369
timestamp 1676037725
transform 1 0 127052 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1381
timestamp 1676037725
transform 1 0 128156 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_1393
timestamp 1676037725
transform 1 0 129260 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1399
timestamp 1676037725
transform 1 0 129812 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1401
timestamp 1676037725
transform 1 0 129996 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1413
timestamp 1676037725
transform 1 0 131100 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1425
timestamp 1676037725
transform 1 0 132204 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1437
timestamp 1676037725
transform 1 0 133308 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_1449
timestamp 1676037725
transform 1 0 134412 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1455
timestamp 1676037725
transform 1 0 134964 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1457
timestamp 1676037725
transform 1 0 135148 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1469
timestamp 1676037725
transform 1 0 136252 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1481
timestamp 1676037725
transform 1 0 137356 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1506
timestamp 1676037725
transform 1 0 139656 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1510
timestamp 1676037725
transform 1 0 140024 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1513
timestamp 1676037725
transform 1 0 140300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1536
timestamp 1676037725
transform 1 0 142416 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_1561
timestamp 1676037725
transform 1 0 144716 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1567
timestamp 1676037725
transform 1 0 145268 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1569
timestamp 1676037725
transform 1 0 145452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1592
timestamp 1676037725
transform 1 0 147568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_1617
timestamp 1676037725
transform 1 0 149868 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1623
timestamp 1676037725
transform 1 0 150420 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1625
timestamp 1676037725
transform 1 0 150604 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1648
timestamp 1676037725
transform 1 0 152720 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1660
timestamp 1676037725
transform 1 0 153824 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_1672
timestamp 1676037725
transform 1 0 154928 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1681
timestamp 1676037725
transform 1 0 155756 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_1725
timestamp 1676037725
transform 1 0 159804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1730
timestamp 1676037725
transform 1 0 160264 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1734
timestamp 1676037725
transform 1 0 160632 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1737
timestamp 1676037725
transform 1 0 160908 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1755
timestamp 1676037725
transform 1 0 162564 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1763
timestamp 1676037725
transform 1 0 163300 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1775
timestamp 1676037725
transform 1 0 164404 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_1787
timestamp 1676037725
transform 1 0 165508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1791
timestamp 1676037725
transform 1 0 165876 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1793
timestamp 1676037725
transform 1 0 166060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_1805
timestamp 1676037725
transform 1 0 167164 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1814
timestamp 1676037725
transform 1 0 167992 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1826
timestamp 1676037725
transform 1 0 169096 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_1838
timestamp 1676037725
transform 1 0 170200 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_1846
timestamp 1676037725
transform 1 0 170936 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1849
timestamp 1676037725
transform 1 0 171212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1861
timestamp 1676037725
transform 1 0 172316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1873
timestamp 1676037725
transform 1 0 173420 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1885
timestamp 1676037725
transform 1 0 174524 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_1897
timestamp 1676037725
transform 1 0 175628 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1903
timestamp 1676037725
transform 1 0 176180 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1905
timestamp 1676037725
transform 1 0 176364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1917
timestamp 1676037725
transform 1 0 177468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1929
timestamp 1676037725
transform 1 0 178572 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1941
timestamp 1676037725
transform 1 0 179676 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_1953
timestamp 1676037725
transform 1 0 180780 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_1959
timestamp 1676037725
transform 1 0 181332 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1961
timestamp 1676037725
transform 1 0 181516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1973
timestamp 1676037725
transform 1 0 182620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1985
timestamp 1676037725
transform 1 0 183724 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_1997
timestamp 1676037725
transform 1 0 184828 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2009
timestamp 1676037725
transform 1 0 185932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2015
timestamp 1676037725
transform 1 0 186484 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2017
timestamp 1676037725
transform 1 0 186668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2029
timestamp 1676037725
transform 1 0 187772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2041
timestamp 1676037725
transform 1 0 188876 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2053
timestamp 1676037725
transform 1 0 189980 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2065
timestamp 1676037725
transform 1 0 191084 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2071
timestamp 1676037725
transform 1 0 191636 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2073
timestamp 1676037725
transform 1 0 191820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2085
timestamp 1676037725
transform 1 0 192924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2097
timestamp 1676037725
transform 1 0 194028 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2109
timestamp 1676037725
transform 1 0 195132 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2121
timestamp 1676037725
transform 1 0 196236 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2127
timestamp 1676037725
transform 1 0 196788 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2129
timestamp 1676037725
transform 1 0 196972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2141
timestamp 1676037725
transform 1 0 198076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2153
timestamp 1676037725
transform 1 0 199180 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2165
timestamp 1676037725
transform 1 0 200284 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2177
timestamp 1676037725
transform 1 0 201388 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2183
timestamp 1676037725
transform 1 0 201940 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2185
timestamp 1676037725
transform 1 0 202124 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2190
timestamp 1676037725
transform 1 0 202584 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2202
timestamp 1676037725
transform 1 0 203688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2205
timestamp 1676037725
transform 1 0 203964 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2228
timestamp 1676037725
transform 1 0 206080 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2241
timestamp 1676037725
transform 1 0 207276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2245
timestamp 1676037725
transform 1 0 207644 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2267
timestamp 1676037725
transform 1 0 209668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2292
timestamp 1676037725
transform 1 0 211968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2297
timestamp 1676037725
transform 1 0 212428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2320
timestamp 1676037725
transform 1 0 214544 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2324
timestamp 1676037725
transform 1 0 214912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2328
timestamp 1676037725
transform 1 0 215280 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2350
timestamp 1676037725
transform 1 0 217304 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2353
timestamp 1676037725
transform 1 0 217580 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2363
timestamp 1676037725
transform 1 0 218500 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2375
timestamp 1676037725
transform 1 0 219604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_2387
timestamp 1676037725
transform 1 0 220708 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2395
timestamp 1676037725
transform 1 0 221444 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2404
timestamp 1676037725
transform 1 0 222272 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2409
timestamp 1676037725
transform 1 0 222732 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2417
timestamp 1676037725
transform 1 0 223468 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2424
timestamp 1676037725
transform 1 0 224112 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2436
timestamp 1676037725
transform 1 0 225216 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2442
timestamp 1676037725
transform 1 0 225768 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2452
timestamp 1676037725
transform 1 0 226688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2460
timestamp 1676037725
transform 1 0 227424 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2465
timestamp 1676037725
transform 1 0 227884 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2471
timestamp 1676037725
transform 1 0 228436 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2483
timestamp 1676037725
transform 1 0 229540 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2495
timestamp 1676037725
transform 1 0 230644 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2507
timestamp 1676037725
transform 1 0 231748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2519
timestamp 1676037725
transform 1 0 232852 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2521
timestamp 1676037725
transform 1 0 233036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2533
timestamp 1676037725
transform 1 0 234140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2545
timestamp 1676037725
transform 1 0 235244 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2554
timestamp 1676037725
transform 1 0 236072 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_2566
timestamp 1676037725
transform 1 0 237176 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2574
timestamp 1676037725
transform 1 0 237912 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2577
timestamp 1676037725
transform 1 0 238188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2589
timestamp 1676037725
transform 1 0 239292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2601
timestamp 1676037725
transform 1 0 240396 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2613
timestamp 1676037725
transform 1 0 241500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2625
timestamp 1676037725
transform 1 0 242604 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2631
timestamp 1676037725
transform 1 0 243156 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2633
timestamp 1676037725
transform 1 0 243340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2645
timestamp 1676037725
transform 1 0 244444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2657
timestamp 1676037725
transform 1 0 245548 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2669
timestamp 1676037725
transform 1 0 246652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2681
timestamp 1676037725
transform 1 0 247756 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2687
timestamp 1676037725
transform 1 0 248308 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2689
timestamp 1676037725
transform 1 0 248492 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2701
timestamp 1676037725
transform 1 0 249596 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2713
timestamp 1676037725
transform 1 0 250700 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2725
timestamp 1676037725
transform 1 0 251804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2737
timestamp 1676037725
transform 1 0 252908 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2743
timestamp 1676037725
transform 1 0 253460 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2745
timestamp 1676037725
transform 1 0 253644 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2757
timestamp 1676037725
transform 1 0 254748 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2769
timestamp 1676037725
transform 1 0 255852 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2781
timestamp 1676037725
transform 1 0 256956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_2787
timestamp 1676037725
transform 1 0 257508 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_2792
timestamp 1676037725
transform 1 0 257968 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2801
timestamp 1676037725
transform 1 0 258796 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2807
timestamp 1676037725
transform 1 0 259348 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2817
timestamp 1676037725
transform 1 0 260268 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2829
timestamp 1676037725
transform 1 0 261372 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2841
timestamp 1676037725
transform 1 0 262476 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_2853
timestamp 1676037725
transform 1 0 263580 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_2857
timestamp 1676037725
transform 1 0 263948 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_2869
timestamp 1676037725
transform 1 0 265052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2875
timestamp 1676037725
transform 1 0 265604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2882
timestamp 1676037725
transform 1 0 266248 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2889
timestamp 1676037725
transform 1 0 266892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2896
timestamp 1676037725
transform 1 0 267536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_2903
timestamp 1676037725
transform 1 0 268180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2910
timestamp 1676037725
transform 1 0 268824 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_2913
timestamp 1676037725
transform 1 0 269100 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_2925
timestamp 1676037725
transform 1 0 270204 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_2934
timestamp 1676037725
transform 1 0 271032 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_264
timestamp 1676037725
transform 1 0 25392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_272
timestamp 1676037725
transform 1 0 26128 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_280
timestamp 1676037725
transform 1 0 26864 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_288
timestamp 1676037725
transform 1 0 27600 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_300
timestamp 1676037725
transform 1 0 28704 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_380
timestamp 1676037725
transform 1 0 36064 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_400
timestamp 1676037725
transform 1 0 37904 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_412
timestamp 1676037725
transform 1 0 39008 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_430
timestamp 1676037725
transform 1 0 40664 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_452
timestamp 1676037725
transform 1 0 42688 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_464
timestamp 1676037725
transform 1 0 43792 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_491
timestamp 1676037725
transform 1 0 46276 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_511
timestamp 1676037725
transform 1 0 48116 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_523
timestamp 1676037725
transform 1 0 49220 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_531
timestamp 1676037725
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_533
timestamp 1676037725
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_545
timestamp 1676037725
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_557
timestamp 1676037725
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_569
timestamp 1676037725
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_581
timestamp 1676037725
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_587
timestamp 1676037725
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_589
timestamp 1676037725
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_601
timestamp 1676037725
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_613
timestamp 1676037725
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_625
timestamp 1676037725
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_637
timestamp 1676037725
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_643
timestamp 1676037725
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_645
timestamp 1676037725
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_657
timestamp 1676037725
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_669
timestamp 1676037725
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_681
timestamp 1676037725
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_693
timestamp 1676037725
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_699
timestamp 1676037725
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_701
timestamp 1676037725
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_713
timestamp 1676037725
transform 1 0 66700 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_722
timestamp 1676037725
transform 1 0 67528 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_734
timestamp 1676037725
transform 1 0 68632 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_746
timestamp 1676037725
transform 1 0 69736 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_754
timestamp 1676037725
transform 1 0 70472 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_757
timestamp 1676037725
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_769
timestamp 1676037725
transform 1 0 71852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_781
timestamp 1676037725
transform 1 0 72956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_793
timestamp 1676037725
transform 1 0 74060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_805
timestamp 1676037725
transform 1 0 75164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_811
timestamp 1676037725
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_813
timestamp 1676037725
transform 1 0 75900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_825
timestamp 1676037725
transform 1 0 77004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_837
timestamp 1676037725
transform 1 0 78108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_849
timestamp 1676037725
transform 1 0 79212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_861
timestamp 1676037725
transform 1 0 80316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_867
timestamp 1676037725
transform 1 0 80868 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_869
timestamp 1676037725
transform 1 0 81052 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_881
timestamp 1676037725
transform 1 0 82156 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_889
timestamp 1676037725
transform 1 0 82892 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_893
timestamp 1676037725
transform 1 0 83260 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_916
timestamp 1676037725
transform 1 0 85376 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_920
timestamp 1676037725
transform 1 0 85744 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_925
timestamp 1676037725
transform 1 0 86204 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_937
timestamp 1676037725
transform 1 0 87308 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_943
timestamp 1676037725
transform 1 0 87860 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_948
timestamp 1676037725
transform 1 0 88320 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_954
timestamp 1676037725
transform 1 0 88872 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_957
timestamp 1676037725
transform 1 0 89148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_969
timestamp 1676037725
transform 1 0 90252 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_977
timestamp 1676037725
transform 1 0 90988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_981
timestamp 1676037725
transform 1 0 91356 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_1006
timestamp 1676037725
transform 1 0 93656 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_1031
timestamp 1676037725
transform 1 0 95956 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1035
timestamp 1676037725
transform 1 0 96324 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1037
timestamp 1676037725
transform 1 0 96508 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1059
timestamp 1676037725
transform 1 0 98532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1063
timestamp 1676037725
transform 1 0 98900 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1067
timestamp 1676037725
transform 1 0 99268 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1090
timestamp 1676037725
transform 1 0 101384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_1093
timestamp 1676037725
transform 1 0 101660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_1117
timestamp 1676037725
transform 1 0 103868 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1123
timestamp 1676037725
transform 1 0 104420 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1146
timestamp 1676037725
transform 1 0 106536 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1149
timestamp 1676037725
transform 1 0 106812 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1153
timestamp 1676037725
transform 1 0 107180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_1165
timestamp 1676037725
transform 1 0 108284 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1173
timestamp 1676037725
transform 1 0 109020 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_1195
timestamp 1676037725
transform 1 0 111044 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1203
timestamp 1676037725
transform 1 0 111780 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1205
timestamp 1676037725
transform 1 0 111964 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1217
timestamp 1676037725
transform 1 0 113068 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_1229
timestamp 1676037725
transform 1 0 114172 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1258
timestamp 1676037725
transform 1 0 116840 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1261
timestamp 1676037725
transform 1 0 117116 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_1273
timestamp 1676037725
transform 1 0 118220 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1281
timestamp 1676037725
transform 1 0 118956 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1304
timestamp 1676037725
transform 1 0 121072 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1317
timestamp 1676037725
transform 1 0 122268 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1325
timestamp 1676037725
transform 1 0 123004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1337
timestamp 1676037725
transform 1 0 124108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1349
timestamp 1676037725
transform 1 0 125212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_1361
timestamp 1676037725
transform 1 0 126316 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_1369
timestamp 1676037725
transform 1 0 127052 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1373
timestamp 1676037725
transform 1 0 127420 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1385
timestamp 1676037725
transform 1 0 128524 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1397
timestamp 1676037725
transform 1 0 129628 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1409
timestamp 1676037725
transform 1 0 130732 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1421
timestamp 1676037725
transform 1 0 131836 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1427
timestamp 1676037725
transform 1 0 132388 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1429
timestamp 1676037725
transform 1 0 132572 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1441
timestamp 1676037725
transform 1 0 133676 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1453
timestamp 1676037725
transform 1 0 134780 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1465
timestamp 1676037725
transform 1 0 135884 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1477
timestamp 1676037725
transform 1 0 136988 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1483
timestamp 1676037725
transform 1 0 137540 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_1485
timestamp 1676037725
transform 1 0 137724 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1493
timestamp 1676037725
transform 1 0 138460 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1496
timestamp 1676037725
transform 1 0 138736 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1519
timestamp 1676037725
transform 1 0 140852 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_1531
timestamp 1676037725
transform 1 0 141956 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1539
timestamp 1676037725
transform 1 0 142692 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1541
timestamp 1676037725
transform 1 0 142876 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_1564
timestamp 1676037725
transform 1 0 144992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1589
timestamp 1676037725
transform 1 0 147292 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1595
timestamp 1676037725
transform 1 0 147844 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1597
timestamp 1676037725
transform 1 0 148028 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1620
timestamp 1676037725
transform 1 0 150144 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1632
timestamp 1676037725
transform 1 0 151248 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_1644
timestamp 1676037725
transform 1 0 152352 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1653
timestamp 1676037725
transform 1 0 153180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_1665
timestamp 1676037725
transform 1 0 154284 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1673
timestamp 1676037725
transform 1 0 155020 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1679
timestamp 1676037725
transform 1 0 155572 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1701
timestamp 1676037725
transform 1 0 157596 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1707
timestamp 1676037725
transform 1 0 158148 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1730
timestamp 1676037725
transform 1 0 160264 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_1734
timestamp 1676037725
transform 1 0 160632 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1757
timestamp 1676037725
transform 1 0 162748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1763
timestamp 1676037725
transform 1 0 163300 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1765
timestamp 1676037725
transform 1 0 163484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1777
timestamp 1676037725
transform 1 0 164588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1789
timestamp 1676037725
transform 1 0 165692 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1801
timestamp 1676037725
transform 1 0 166796 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1813
timestamp 1676037725
transform 1 0 167900 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1819
timestamp 1676037725
transform 1 0 168452 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1821
timestamp 1676037725
transform 1 0 168636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1833
timestamp 1676037725
transform 1 0 169740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1845
timestamp 1676037725
transform 1 0 170844 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1857
timestamp 1676037725
transform 1 0 171948 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1869
timestamp 1676037725
transform 1 0 173052 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1875
timestamp 1676037725
transform 1 0 173604 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1877
timestamp 1676037725
transform 1 0 173788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1889
timestamp 1676037725
transform 1 0 174892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1901
timestamp 1676037725
transform 1 0 175996 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1913
timestamp 1676037725
transform 1 0 177100 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1925
timestamp 1676037725
transform 1 0 178204 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1931
timestamp 1676037725
transform 1 0 178756 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1933
timestamp 1676037725
transform 1 0 178940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1945
timestamp 1676037725
transform 1 0 180044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1957
timestamp 1676037725
transform 1 0 181148 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1969
timestamp 1676037725
transform 1 0 182252 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_1981
timestamp 1676037725
transform 1 0 183356 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_1987
timestamp 1676037725
transform 1 0 183908 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_1989
timestamp 1676037725
transform 1 0 184092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2001
timestamp 1676037725
transform 1 0 185196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2013
timestamp 1676037725
transform 1 0 186300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2025
timestamp 1676037725
transform 1 0 187404 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_2037
timestamp 1676037725
transform 1 0 188508 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2043
timestamp 1676037725
transform 1 0 189060 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2045
timestamp 1676037725
transform 1 0 189244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2057
timestamp 1676037725
transform 1 0 190348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2069
timestamp 1676037725
transform 1 0 191452 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2081
timestamp 1676037725
transform 1 0 192556 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_2093
timestamp 1676037725
transform 1 0 193660 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2099
timestamp 1676037725
transform 1 0 194212 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2101
timestamp 1676037725
transform 1 0 194396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2113
timestamp 1676037725
transform 1 0 195500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2125
timestamp 1676037725
transform 1 0 196604 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2137
timestamp 1676037725
transform 1 0 197708 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_2149
timestamp 1676037725
transform 1 0 198812 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2155
timestamp 1676037725
transform 1 0 199364 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2157
timestamp 1676037725
transform 1 0 199548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2169
timestamp 1676037725
transform 1 0 200652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2181
timestamp 1676037725
transform 1 0 201756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_2193
timestamp 1676037725
transform 1 0 202860 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_2201
timestamp 1676037725
transform 1 0 203596 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2206
timestamp 1676037725
transform 1 0 204056 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2210
timestamp 1676037725
transform 1 0 204424 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2213
timestamp 1676037725
transform 1 0 204700 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2236
timestamp 1676037725
transform 1 0 206816 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2261
timestamp 1676037725
transform 1 0 209116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_2265
timestamp 1676037725
transform 1 0 209484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2269
timestamp 1676037725
transform 1 0 209852 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_2273
timestamp 1676037725
transform 1 0 210220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2318
timestamp 1676037725
transform 1 0 214360 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2322
timestamp 1676037725
transform 1 0 214728 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2325
timestamp 1676037725
transform 1 0 215004 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2348
timestamp 1676037725
transform 1 0 217120 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_2373
timestamp 1676037725
transform 1 0 219420 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2379
timestamp 1676037725
transform 1 0 219972 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2381
timestamp 1676037725
transform 1 0 220156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2393
timestamp 1676037725
transform 1 0 221260 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2405
timestamp 1676037725
transform 1 0 222364 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2410
timestamp 1676037725
transform 1 0 222824 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2422
timestamp 1676037725
transform 1 0 223928 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2434
timestamp 1676037725
transform 1 0 225032 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2437
timestamp 1676037725
transform 1 0 225308 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2460
timestamp 1676037725
transform 1 0 227424 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2464
timestamp 1676037725
transform 1 0 227792 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2476
timestamp 1676037725
transform 1 0 228896 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2488
timestamp 1676037725
transform 1 0 230000 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2493
timestamp 1676037725
transform 1 0 230460 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2499
timestamp 1676037725
transform 1 0 231012 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2511
timestamp 1676037725
transform 1 0 232116 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2523
timestamp 1676037725
transform 1 0 233220 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2535
timestamp 1676037725
transform 1 0 234324 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2547
timestamp 1676037725
transform 1 0 235428 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2549
timestamp 1676037725
transform 1 0 235612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2561
timestamp 1676037725
transform 1 0 236716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2573
timestamp 1676037725
transform 1 0 237820 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2585
timestamp 1676037725
transform 1 0 238924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_2597
timestamp 1676037725
transform 1 0 240028 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2603
timestamp 1676037725
transform 1 0 240580 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2605
timestamp 1676037725
transform 1 0 240764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2617
timestamp 1676037725
transform 1 0 241868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2629
timestamp 1676037725
transform 1 0 242972 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2641
timestamp 1676037725
transform 1 0 244076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_2653
timestamp 1676037725
transform 1 0 245180 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2659
timestamp 1676037725
transform 1 0 245732 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2661
timestamp 1676037725
transform 1 0 245916 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2673
timestamp 1676037725
transform 1 0 247020 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2685
timestamp 1676037725
transform 1 0 248124 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2697
timestamp 1676037725
transform 1 0 249228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_2709
timestamp 1676037725
transform 1 0 250332 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2715
timestamp 1676037725
transform 1 0 250884 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_2717
timestamp 1676037725
transform 1 0 251068 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2725
timestamp 1676037725
transform 1 0 251804 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2733
timestamp 1676037725
transform 1 0 252540 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2745
timestamp 1676037725
transform 1 0 253644 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2757
timestamp 1676037725
transform 1 0 254748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_2769
timestamp 1676037725
transform 1 0 255852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2773
timestamp 1676037725
transform 1 0 256220 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2777
timestamp 1676037725
transform 1 0 256588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_2789
timestamp 1676037725
transform 1 0 257692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2798
timestamp 1676037725
transform 1 0 258520 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2808
timestamp 1676037725
transform 1 0 259440 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2818
timestamp 1676037725
transform 1 0 260360 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_2822
timestamp 1676037725
transform 1 0 260728 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2829
timestamp 1676037725
transform 1 0 261372 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2841
timestamp 1676037725
transform 1 0 262476 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_2853
timestamp 1676037725
transform 1 0 263580 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_2865
timestamp 1676037725
transform 1 0 264684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2871
timestamp 1676037725
transform 1 0 265236 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2875
timestamp 1676037725
transform 1 0 265604 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_2882
timestamp 1676037725
transform 1 0 266248 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_2885
timestamp 1676037725
transform 1 0 266524 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_2891
timestamp 1676037725
transform 1 0 267076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2895
timestamp 1676037725
transform 1 0 267444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2902
timestamp 1676037725
transform 1 0 268088 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2909
timestamp 1676037725
transform 1 0 268732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2917
timestamp 1676037725
transform 1 0 269468 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2925
timestamp 1676037725
transform 1 0 270204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_2932
timestamp 1676037725
transform 1 0 270848 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_267
timestamp 1676037725
transform 1 0 25668 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_272
timestamp 1676037725
transform 1 0 26128 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_417
timestamp 1676037725
transform 1 0 39468 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_425
timestamp 1676037725
transform 1 0 40204 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_445
timestamp 1676037725
transform 1 0 42044 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_473
timestamp 1676037725
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_485
timestamp 1676037725
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_497
timestamp 1676037725
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_503
timestamp 1676037725
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_514
timestamp 1676037725
transform 1 0 48392 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_536
timestamp 1676037725
transform 1 0 50416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_558
timestamp 1676037725
transform 1 0 52440 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_561
timestamp 1676037725
transform 1 0 52716 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_567
timestamp 1676037725
transform 1 0 53268 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_579
timestamp 1676037725
transform 1 0 54372 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_591
timestamp 1676037725
transform 1 0 55476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_603
timestamp 1676037725
transform 1 0 56580 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_615
timestamp 1676037725
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_617
timestamp 1676037725
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_629
timestamp 1676037725
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_641
timestamp 1676037725
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_653
timestamp 1676037725
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_665
timestamp 1676037725
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_671
timestamp 1676037725
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_673
timestamp 1676037725
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_685
timestamp 1676037725
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_697
timestamp 1676037725
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_709
timestamp 1676037725
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_721
timestamp 1676037725
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_727
timestamp 1676037725
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_729
timestamp 1676037725
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_741
timestamp 1676037725
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_753
timestamp 1676037725
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_765
timestamp 1676037725
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_777
timestamp 1676037725
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_783
timestamp 1676037725
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_785
timestamp 1676037725
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_797
timestamp 1676037725
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_809
timestamp 1676037725
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_821
timestamp 1676037725
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_833
timestamp 1676037725
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_839
timestamp 1676037725
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_841
timestamp 1676037725
transform 1 0 78476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_853
timestamp 1676037725
transform 1 0 79580 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_867
timestamp 1676037725
transform 1 0 80868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_871
timestamp 1676037725
transform 1 0 81236 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_894
timestamp 1676037725
transform 1 0 83352 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_897
timestamp 1676037725
transform 1 0 83628 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_901
timestamp 1676037725
transform 1 0 83996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_907
timestamp 1676037725
transform 1 0 84548 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_930
timestamp 1676037725
transform 1 0 86664 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_934
timestamp 1676037725
transform 1 0 87032 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_946
timestamp 1676037725
transform 1 0 88136 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_953
timestamp 1676037725
transform 1 0 88780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_965
timestamp 1676037725
transform 1 0 89884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_977
timestamp 1676037725
transform 1 0 90988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_989
timestamp 1676037725
transform 1 0 92092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_1001
timestamp 1676037725
transform 1 0 93196 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1007
timestamp 1676037725
transform 1 0 93748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_1009
timestamp 1676037725
transform 1 0 93932 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1034
timestamp 1676037725
transform 1 0 96232 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1046
timestamp 1676037725
transform 1 0 97336 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1058
timestamp 1676037725
transform 1 0 98440 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1062
timestamp 1676037725
transform 1 0 98808 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_1065
timestamp 1676037725
transform 1 0 99084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1089
timestamp 1676037725
transform 1 0 101292 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1093
timestamp 1676037725
transform 1 0 101660 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1105
timestamp 1676037725
transform 1 0 102764 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1117
timestamp 1676037725
transform 1 0 103868 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1121
timestamp 1676037725
transform 1 0 104236 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_1125
timestamp 1676037725
transform 1 0 104604 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_1149
timestamp 1676037725
transform 1 0 106812 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1174
timestamp 1676037725
transform 1 0 109112 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1177
timestamp 1676037725
transform 1 0 109388 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1189
timestamp 1676037725
transform 1 0 110492 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_1201
timestamp 1676037725
transform 1 0 111596 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1230
timestamp 1676037725
transform 1 0 114264 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1233
timestamp 1676037725
transform 1 0 114540 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1255
timestamp 1676037725
transform 1 0 116564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1259
timestamp 1676037725
transform 1 0 116932 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1263
timestamp 1676037725
transform 1 0 117300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1286
timestamp 1676037725
transform 1 0 119416 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1289
timestamp 1676037725
transform 1 0 119692 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_1293
timestamp 1676037725
transform 1 0 120060 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1301
timestamp 1676037725
transform 1 0 120796 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1305
timestamp 1676037725
transform 1 0 121164 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1309
timestamp 1676037725
transform 1 0 121532 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1332
timestamp 1676037725
transform 1 0 123648 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_1336
timestamp 1676037725
transform 1 0 124016 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1345
timestamp 1676037725
transform 1 0 124844 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1357
timestamp 1676037725
transform 1 0 125948 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1369
timestamp 1676037725
transform 1 0 127052 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1381
timestamp 1676037725
transform 1 0 128156 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_1393
timestamp 1676037725
transform 1 0 129260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1399
timestamp 1676037725
transform 1 0 129812 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1401
timestamp 1676037725
transform 1 0 129996 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1413
timestamp 1676037725
transform 1 0 131100 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1425
timestamp 1676037725
transform 1 0 132204 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1437
timestamp 1676037725
transform 1 0 133308 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_1449
timestamp 1676037725
transform 1 0 134412 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1455
timestamp 1676037725
transform 1 0 134964 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1457
timestamp 1676037725
transform 1 0 135148 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1469
timestamp 1676037725
transform 1 0 136252 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1481
timestamp 1676037725
transform 1 0 137356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1493
timestamp 1676037725
transform 1 0 138460 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_1505
timestamp 1676037725
transform 1 0 139564 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1511
timestamp 1676037725
transform 1 0 140116 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1513
timestamp 1676037725
transform 1 0 140300 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1527
timestamp 1676037725
transform 1 0 141588 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1550
timestamp 1676037725
transform 1 0 143704 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_1554
timestamp 1676037725
transform 1 0 144072 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1562
timestamp 1676037725
transform 1 0 144808 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1566
timestamp 1676037725
transform 1 0 145176 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1569
timestamp 1676037725
transform 1 0 145452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1592
timestamp 1676037725
transform 1 0 147568 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_1617
timestamp 1676037725
transform 1 0 149868 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1623
timestamp 1676037725
transform 1 0 150420 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1625
timestamp 1676037725
transform 1 0 150604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_1658
timestamp 1676037725
transform 1 0 153640 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1666
timestamp 1676037725
transform 1 0 154376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1674
timestamp 1676037725
transform 1 0 155112 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1678
timestamp 1676037725
transform 1 0 155480 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1681
timestamp 1676037725
transform 1 0 155756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_1693
timestamp 1676037725
transform 1 0 156860 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1701
timestamp 1676037725
transform 1 0 157596 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1704
timestamp 1676037725
transform 1 0 157872 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_1729
timestamp 1676037725
transform 1 0 160172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1734
timestamp 1676037725
transform 1 0 160632 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1737
timestamp 1676037725
transform 1 0 160908 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1760
timestamp 1676037725
transform 1 0 163024 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_1764
timestamp 1676037725
transform 1 0 163392 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1768
timestamp 1676037725
transform 1 0 163760 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1780
timestamp 1676037725
transform 1 0 164864 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1793
timestamp 1676037725
transform 1 0 166060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1805
timestamp 1676037725
transform 1 0 167164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1817
timestamp 1676037725
transform 1 0 168268 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1829
timestamp 1676037725
transform 1 0 169372 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_1841
timestamp 1676037725
transform 1 0 170476 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1847
timestamp 1676037725
transform 1 0 171028 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1849
timestamp 1676037725
transform 1 0 171212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1861
timestamp 1676037725
transform 1 0 172316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1873
timestamp 1676037725
transform 1 0 173420 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1885
timestamp 1676037725
transform 1 0 174524 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_1897
timestamp 1676037725
transform 1 0 175628 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1903
timestamp 1676037725
transform 1 0 176180 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1905
timestamp 1676037725
transform 1 0 176364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1917
timestamp 1676037725
transform 1 0 177468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1929
timestamp 1676037725
transform 1 0 178572 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1941
timestamp 1676037725
transform 1 0 179676 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_1953
timestamp 1676037725
transform 1 0 180780 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_1959
timestamp 1676037725
transform 1 0 181332 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1961
timestamp 1676037725
transform 1 0 181516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1973
timestamp 1676037725
transform 1 0 182620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1985
timestamp 1676037725
transform 1 0 183724 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_1997
timestamp 1676037725
transform 1 0 184828 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_2009
timestamp 1676037725
transform 1 0 185932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2015
timestamp 1676037725
transform 1 0 186484 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2017
timestamp 1676037725
transform 1 0 186668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2029
timestamp 1676037725
transform 1 0 187772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_2041
timestamp 1676037725
transform 1 0 188876 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_2049
timestamp 1676037725
transform 1 0 189612 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2058
timestamp 1676037725
transform 1 0 190440 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2070
timestamp 1676037725
transform 1 0 191544 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2073
timestamp 1676037725
transform 1 0 191820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2085
timestamp 1676037725
transform 1 0 192924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2097
timestamp 1676037725
transform 1 0 194028 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2109
timestamp 1676037725
transform 1 0 195132 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_2121
timestamp 1676037725
transform 1 0 196236 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2127
timestamp 1676037725
transform 1 0 196788 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2129
timestamp 1676037725
transform 1 0 196972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2141
timestamp 1676037725
transform 1 0 198076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2153
timestamp 1676037725
transform 1 0 199180 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2165
timestamp 1676037725
transform 1 0 200284 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_2177
timestamp 1676037725
transform 1 0 201388 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2183
timestamp 1676037725
transform 1 0 201940 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2185
timestamp 1676037725
transform 1 0 202124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2197
timestamp 1676037725
transform 1 0 203228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2209
timestamp 1676037725
transform 1 0 204332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_2221
timestamp 1676037725
transform 1 0 205436 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_2229
timestamp 1676037725
transform 1 0 206172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2234
timestamp 1676037725
transform 1 0 206632 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2238
timestamp 1676037725
transform 1 0 207000 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2241
timestamp 1676037725
transform 1 0 207276 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2264
timestamp 1676037725
transform 1 0 209392 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2289
timestamp 1676037725
transform 1 0 211692 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_2293
timestamp 1676037725
transform 1 0 212060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2297
timestamp 1676037725
transform 1 0 212428 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2322
timestamp 1676037725
transform 1 0 214728 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_2345
timestamp 1676037725
transform 1 0 216844 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2351
timestamp 1676037725
transform 1 0 217396 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2353
timestamp 1676037725
transform 1 0 217580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2365
timestamp 1676037725
transform 1 0 218684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2377
timestamp 1676037725
transform 1 0 219788 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2389
timestamp 1676037725
transform 1 0 220892 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_2401
timestamp 1676037725
transform 1 0 221996 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2407
timestamp 1676037725
transform 1 0 222548 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2409
timestamp 1676037725
transform 1 0 222732 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2421
timestamp 1676037725
transform 1 0 223836 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2424
timestamp 1676037725
transform 1 0 224112 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2447
timestamp 1676037725
transform 1 0 226228 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_2457
timestamp 1676037725
transform 1 0 227148 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2462
timestamp 1676037725
transform 1 0 227608 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2465
timestamp 1676037725
transform 1 0 227884 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2488
timestamp 1676037725
transform 1 0 230000 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2496
timestamp 1676037725
transform 1 0 230736 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2508
timestamp 1676037725
transform 1 0 231840 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2521
timestamp 1676037725
transform 1 0 233036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2533
timestamp 1676037725
transform 1 0 234140 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_2545
timestamp 1676037725
transform 1 0 235244 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2554
timestamp 1676037725
transform 1 0 236072 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_2566
timestamp 1676037725
transform 1 0 237176 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2574
timestamp 1676037725
transform 1 0 237912 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2577
timestamp 1676037725
transform 1 0 238188 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_2589
timestamp 1676037725
transform 1 0 239292 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_2597
timestamp 1676037725
transform 1 0 240028 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2606
timestamp 1676037725
transform 1 0 240856 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2618
timestamp 1676037725
transform 1 0 241960 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_2626
timestamp 1676037725
transform 1 0 242696 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2633
timestamp 1676037725
transform 1 0 243340 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2637
timestamp 1676037725
transform 1 0 243708 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2644
timestamp 1676037725
transform 1 0 244352 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2656
timestamp 1676037725
transform 1 0 245456 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2668
timestamp 1676037725
transform 1 0 246560 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_2680
timestamp 1676037725
transform 1 0 247664 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2689
timestamp 1676037725
transform 1 0 248492 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2701
timestamp 1676037725
transform 1 0 249596 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2713
timestamp 1676037725
transform 1 0 250700 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2716
timestamp 1676037725
transform 1 0 250976 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2720
timestamp 1676037725
transform 1 0 251344 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2724
timestamp 1676037725
transform 1 0 251712 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2735
timestamp 1676037725
transform 1 0 252724 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2739
timestamp 1676037725
transform 1 0 253092 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2743
timestamp 1676037725
transform 1 0 253460 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2745
timestamp 1676037725
transform 1 0 253644 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2756
timestamp 1676037725
transform 1 0 254656 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2760
timestamp 1676037725
transform 1 0 255024 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_2764
timestamp 1676037725
transform 1 0 255392 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2769
timestamp 1676037725
transform 1 0 255852 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_2773
timestamp 1676037725
transform 1 0 256220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2784
timestamp 1676037725
transform 1 0 257232 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2796
timestamp 1676037725
transform 1 0 258336 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_2801
timestamp 1676037725
transform 1 0 258796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_2806
timestamp 1676037725
transform 1 0 259256 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2821
timestamp 1676037725
transform 1 0 260636 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2829
timestamp 1676037725
transform 1 0 261372 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_2841
timestamp 1676037725
transform 1 0 262476 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_2853
timestamp 1676037725
transform 1 0 263580 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2857
timestamp 1676037725
transform 1 0 263948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_2861
timestamp 1676037725
transform 1 0 264316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2865
timestamp 1676037725
transform 1 0 264684 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2872
timestamp 1676037725
transform 1 0 265328 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2879
timestamp 1676037725
transform 1 0 265972 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2886
timestamp 1676037725
transform 1 0 266616 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2893
timestamp 1676037725
transform 1 0 267260 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2901
timestamp 1676037725
transform 1 0 267996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2910
timestamp 1676037725
transform 1 0 268824 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2913
timestamp 1676037725
transform 1 0 269100 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2919
timestamp 1676037725
transform 1 0 269652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_2927
timestamp 1676037725
transform 1 0 270388 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_2934
timestamp 1676037725
transform 1 0 271032 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1676037725
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1676037725
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1676037725
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1676037725
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1676037725
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_425
timestamp 1676037725
transform 1 0 40204 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_429
timestamp 1676037725
transform 1 0 40572 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_449
timestamp 1676037725
transform 1 0 42412 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_471
timestamp 1676037725
transform 1 0 44436 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_475
timestamp 1676037725
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_481
timestamp 1676037725
transform 1 0 45356 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_493
timestamp 1676037725
transform 1 0 46460 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_497
timestamp 1676037725
transform 1 0 46828 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_500
timestamp 1676037725
transform 1 0 47104 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_520
timestamp 1676037725
transform 1 0 48944 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_533
timestamp 1676037725
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_545
timestamp 1676037725
transform 1 0 51244 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_551
timestamp 1676037725
transform 1 0 51796 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_570
timestamp 1676037725
transform 1 0 53544 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_582
timestamp 1676037725
transform 1 0 54648 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_589
timestamp 1676037725
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_601
timestamp 1676037725
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_613
timestamp 1676037725
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_625
timestamp 1676037725
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_637
timestamp 1676037725
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_643
timestamp 1676037725
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_645
timestamp 1676037725
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_657
timestamp 1676037725
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_669
timestamp 1676037725
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_681
timestamp 1676037725
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_693
timestamp 1676037725
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_699
timestamp 1676037725
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_701
timestamp 1676037725
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_713
timestamp 1676037725
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_725
timestamp 1676037725
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_737
timestamp 1676037725
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_749
timestamp 1676037725
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_755
timestamp 1676037725
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_757
timestamp 1676037725
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_769
timestamp 1676037725
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_781
timestamp 1676037725
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_793
timestamp 1676037725
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_805
timestamp 1676037725
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_811
timestamp 1676037725
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_813
timestamp 1676037725
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_825
timestamp 1676037725
transform 1 0 77004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_837
timestamp 1676037725
transform 1 0 78108 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_849
timestamp 1676037725
transform 1 0 79212 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_857
timestamp 1676037725
transform 1 0 79948 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_862
timestamp 1676037725
transform 1 0 80408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_866
timestamp 1676037725
transform 1 0 80776 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_869
timestamp 1676037725
transform 1 0 81052 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_874
timestamp 1676037725
transform 1 0 81512 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_897
timestamp 1676037725
transform 1 0 83628 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_922
timestamp 1676037725
transform 1 0 85928 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_925
timestamp 1676037725
transform 1 0 86204 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_929
timestamp 1676037725
transform 1 0 86572 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_933
timestamp 1676037725
transform 1 0 86940 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_937
timestamp 1676037725
transform 1 0 87308 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_941
timestamp 1676037725
transform 1 0 87676 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_964
timestamp 1676037725
transform 1 0 89792 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_968
timestamp 1676037725
transform 1 0 90160 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_972
timestamp 1676037725
transform 1 0 90528 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_976
timestamp 1676037725
transform 1 0 90896 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_981
timestamp 1676037725
transform 1 0 91356 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1017
timestamp 1676037725
transform 1 0 94668 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_1027
timestamp 1676037725
transform 1 0 95588 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1035
timestamp 1676037725
transform 1 0 96324 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1037
timestamp 1676037725
transform 1 0 96508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1049
timestamp 1676037725
transform 1 0 97612 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_1061
timestamp 1676037725
transform 1 0 98716 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1067
timestamp 1676037725
transform 1 0 99268 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1078
timestamp 1676037725
transform 1 0 100280 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1090
timestamp 1676037725
transform 1 0 101384 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1093
timestamp 1676037725
transform 1 0 101660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1105
timestamp 1676037725
transform 1 0 102764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1117
timestamp 1676037725
transform 1 0 103868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1129
timestamp 1676037725
transform 1 0 104972 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_1141
timestamp 1676037725
transform 1 0 106076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1147
timestamp 1676037725
transform 1 0 106628 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1149
timestamp 1676037725
transform 1 0 106812 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1172
timestamp 1676037725
transform 1 0 108928 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1176
timestamp 1676037725
transform 1 0 109296 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1179
timestamp 1676037725
transform 1 0 109572 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1202
timestamp 1676037725
transform 1 0 111688 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1205
timestamp 1676037725
transform 1 0 111964 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_1217
timestamp 1676037725
transform 1 0 113068 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1222
timestamp 1676037725
transform 1 0 113528 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1226
timestamp 1676037725
transform 1 0 113896 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1249
timestamp 1676037725
transform 1 0 116012 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_1253
timestamp 1676037725
transform 1 0 116380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1259
timestamp 1676037725
transform 1 0 116932 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1261
timestamp 1676037725
transform 1 0 117116 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1294
timestamp 1676037725
transform 1 0 120152 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1298
timestamp 1676037725
transform 1 0 120520 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_1306
timestamp 1676037725
transform 1 0 121256 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1314
timestamp 1676037725
transform 1 0 121992 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1317
timestamp 1676037725
transform 1 0 122268 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1340
timestamp 1676037725
transform 1 0 124384 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1344
timestamp 1676037725
transform 1 0 124752 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1356
timestamp 1676037725
transform 1 0 125856 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1368
timestamp 1676037725
transform 1 0 126960 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1373
timestamp 1676037725
transform 1 0 127420 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1385
timestamp 1676037725
transform 1 0 128524 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1397
timestamp 1676037725
transform 1 0 129628 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1409
timestamp 1676037725
transform 1 0 130732 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_1421
timestamp 1676037725
transform 1 0 131836 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1427
timestamp 1676037725
transform 1 0 132388 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1429
timestamp 1676037725
transform 1 0 132572 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1441
timestamp 1676037725
transform 1 0 133676 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1453
timestamp 1676037725
transform 1 0 134780 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1465
timestamp 1676037725
transform 1 0 135884 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_1477
timestamp 1676037725
transform 1 0 136988 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1483
timestamp 1676037725
transform 1 0 137540 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1485
timestamp 1676037725
transform 1 0 137724 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1497
timestamp 1676037725
transform 1 0 138828 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1509
timestamp 1676037725
transform 1 0 139932 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1521
timestamp 1676037725
transform 1 0 141036 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_1533
timestamp 1676037725
transform 1 0 142140 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1538
timestamp 1676037725
transform 1 0 142600 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1541
timestamp 1676037725
transform 1 0 142876 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1564
timestamp 1676037725
transform 1 0 144992 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1568
timestamp 1676037725
transform 1 0 145360 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1580
timestamp 1676037725
transform 1 0 146464 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1592
timestamp 1676037725
transform 1 0 147568 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1597
timestamp 1676037725
transform 1 0 148028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1609
timestamp 1676037725
transform 1 0 149132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_1621
timestamp 1676037725
transform 1 0 150236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_1645
timestamp 1676037725
transform 1 0 152444 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1651
timestamp 1676037725
transform 1 0 152996 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1674
timestamp 1676037725
transform 1 0 155112 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_1678
timestamp 1676037725
transform 1 0 155480 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1682
timestamp 1676037725
transform 1 0 155848 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1704
timestamp 1676037725
transform 1 0 157872 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1730
timestamp 1676037725
transform 1 0 160264 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1734
timestamp 1676037725
transform 1 0 160632 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_1759
timestamp 1676037725
transform 1 0 162932 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1763
timestamp 1676037725
transform 1 0 163300 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1765
timestamp 1676037725
transform 1 0 163484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1777
timestamp 1676037725
transform 1 0 164588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1789
timestamp 1676037725
transform 1 0 165692 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1801
timestamp 1676037725
transform 1 0 166796 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_1813
timestamp 1676037725
transform 1 0 167900 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1819
timestamp 1676037725
transform 1 0 168452 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1821
timestamp 1676037725
transform 1 0 168636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1833
timestamp 1676037725
transform 1 0 169740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1845
timestamp 1676037725
transform 1 0 170844 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1857
timestamp 1676037725
transform 1 0 171948 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_1869
timestamp 1676037725
transform 1 0 173052 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1875
timestamp 1676037725
transform 1 0 173604 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1877
timestamp 1676037725
transform 1 0 173788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1889
timestamp 1676037725
transform 1 0 174892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1901
timestamp 1676037725
transform 1 0 175996 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1913
timestamp 1676037725
transform 1 0 177100 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_1925
timestamp 1676037725
transform 1 0 178204 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1931
timestamp 1676037725
transform 1 0 178756 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1933
timestamp 1676037725
transform 1 0 178940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1945
timestamp 1676037725
transform 1 0 180044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1957
timestamp 1676037725
transform 1 0 181148 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1969
timestamp 1676037725
transform 1 0 182252 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_1981
timestamp 1676037725
transform 1 0 183356 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_1987
timestamp 1676037725
transform 1 0 183908 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_1989
timestamp 1676037725
transform 1 0 184092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2001
timestamp 1676037725
transform 1 0 185196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2013
timestamp 1676037725
transform 1 0 186300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2025
timestamp 1676037725
transform 1 0 187404 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_2037
timestamp 1676037725
transform 1 0 188508 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2043
timestamp 1676037725
transform 1 0 189060 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2045
timestamp 1676037725
transform 1 0 189244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2057
timestamp 1676037725
transform 1 0 190348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2069
timestamp 1676037725
transform 1 0 191452 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2081
timestamp 1676037725
transform 1 0 192556 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_2093
timestamp 1676037725
transform 1 0 193660 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2099
timestamp 1676037725
transform 1 0 194212 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2101
timestamp 1676037725
transform 1 0 194396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2113
timestamp 1676037725
transform 1 0 195500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2125
timestamp 1676037725
transform 1 0 196604 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2137
timestamp 1676037725
transform 1 0 197708 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_2149
timestamp 1676037725
transform 1 0 198812 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2155
timestamp 1676037725
transform 1 0 199364 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2157
timestamp 1676037725
transform 1 0 199548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2169
timestamp 1676037725
transform 1 0 200652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2181
timestamp 1676037725
transform 1 0 201756 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2193
timestamp 1676037725
transform 1 0 202860 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_2205
timestamp 1676037725
transform 1 0 203964 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2211
timestamp 1676037725
transform 1 0 204516 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2213
timestamp 1676037725
transform 1 0 204700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2225
timestamp 1676037725
transform 1 0 205804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2237
timestamp 1676037725
transform 1 0 206908 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2249
timestamp 1676037725
transform 1 0 208012 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_2261
timestamp 1676037725
transform 1 0 209116 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2267
timestamp 1676037725
transform 1 0 209668 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2269
timestamp 1676037725
transform 1 0 209852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2281
timestamp 1676037725
transform 1 0 210956 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_2293
timestamp 1676037725
transform 1 0 212060 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_2317
timestamp 1676037725
transform 1 0 214268 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2323
timestamp 1676037725
transform 1 0 214820 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2325
timestamp 1676037725
transform 1 0 215004 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2348
timestamp 1676037725
transform 1 0 217120 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2352
timestamp 1676037725
transform 1 0 217488 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2364
timestamp 1676037725
transform 1 0 218592 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2378
timestamp 1676037725
transform 1 0 219880 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2381
timestamp 1676037725
transform 1 0 220156 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2385
timestamp 1676037725
transform 1 0 220524 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2407
timestamp 1676037725
transform 1 0 222548 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2411
timestamp 1676037725
transform 1 0 222916 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2415
timestamp 1676037725
transform 1 0 223284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_2427
timestamp 1676037725
transform 1 0 224388 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2432
timestamp 1676037725
transform 1 0 224848 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2437
timestamp 1676037725
transform 1 0 225308 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2441
timestamp 1676037725
transform 1 0 225676 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2444
timestamp 1676037725
transform 1 0 225952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2448
timestamp 1676037725
transform 1 0 226320 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2471
timestamp 1676037725
transform 1 0 228436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_2486
timestamp 1676037725
transform 1 0 229816 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2493
timestamp 1676037725
transform 1 0 230460 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2505
timestamp 1676037725
transform 1 0 231564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2517
timestamp 1676037725
transform 1 0 232668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2529
timestamp 1676037725
transform 1 0 233772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_2541
timestamp 1676037725
transform 1 0 234876 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2547
timestamp 1676037725
transform 1 0 235428 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2549
timestamp 1676037725
transform 1 0 235612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2561
timestamp 1676037725
transform 1 0 236716 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2573
timestamp 1676037725
transform 1 0 237820 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2577
timestamp 1676037725
transform 1 0 238188 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2580
timestamp 1676037725
transform 1 0 238464 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2584
timestamp 1676037725
transform 1 0 238832 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2594
timestamp 1676037725
transform 1 0 239752 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2598
timestamp 1676037725
transform 1 0 240120 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2602
timestamp 1676037725
transform 1 0 240488 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2605
timestamp 1676037725
transform 1 0 240764 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2615
timestamp 1676037725
transform 1 0 241684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2619
timestamp 1676037725
transform 1 0 242052 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2623
timestamp 1676037725
transform 1 0 242420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2633
timestamp 1676037725
transform 1 0 243340 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2637
timestamp 1676037725
transform 1 0 243708 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2647
timestamp 1676037725
transform 1 0 244628 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_2657
timestamp 1676037725
transform 1 0 245548 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2661
timestamp 1676037725
transform 1 0 245916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2673
timestamp 1676037725
transform 1 0 247020 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2685
timestamp 1676037725
transform 1 0 248124 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2697
timestamp 1676037725
transform 1 0 249228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_2709
timestamp 1676037725
transform 1 0 250332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2714
timestamp 1676037725
transform 1 0 250792 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2717
timestamp 1676037725
transform 1 0 251068 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2727
timestamp 1676037725
transform 1 0 251988 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2731
timestamp 1676037725
transform 1 0 252356 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2743
timestamp 1676037725
transform 1 0 253460 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2746
timestamp 1676037725
transform 1 0 253736 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2750
timestamp 1676037725
transform 1 0 254104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2761
timestamp 1676037725
transform 1 0 255116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_2765
timestamp 1676037725
transform 1 0 255484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2770
timestamp 1676037725
transform 1 0 255944 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2773
timestamp 1676037725
transform 1 0 256220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2777
timestamp 1676037725
transform 1 0 256588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2780
timestamp 1676037725
transform 1 0 256864 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2790
timestamp 1676037725
transform 1 0 257784 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2802
timestamp 1676037725
transform 1 0 258888 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2808
timestamp 1676037725
transform 1 0 259440 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2824
timestamp 1676037725
transform 1 0 260912 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_2829
timestamp 1676037725
transform 1 0 261372 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_2841
timestamp 1676037725
transform 1 0 262476 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2850
timestamp 1676037725
transform 1 0 263304 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_2863
timestamp 1676037725
transform 1 0 264500 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2869
timestamp 1676037725
transform 1 0 265052 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2873
timestamp 1676037725
transform 1 0 265420 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2882
timestamp 1676037725
transform 1 0 266248 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_2885
timestamp 1676037725
transform 1 0 266524 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2891
timestamp 1676037725
transform 1 0 267076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2898
timestamp 1676037725
transform 1 0 267720 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2911
timestamp 1676037725
transform 1 0 268916 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_2920
timestamp 1676037725
transform 1 0 269744 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_2929
timestamp 1676037725
transform 1 0 270572 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_2935
timestamp 1676037725
transform 1 0 271124 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_413
timestamp 1676037725
transform 1 0 39100 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_425
timestamp 1676037725
transform 1 0 40204 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_437
timestamp 1676037725
transform 1 0 41308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_446
timestamp 1676037725
transform 1 0 42136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_454
timestamp 1676037725
transform 1 0 42872 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_475
timestamp 1676037725
transform 1 0 44804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_483
timestamp 1676037725
transform 1 0 45540 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_502
timestamp 1676037725
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_513
timestamp 1676037725
transform 1 0 48300 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_525
timestamp 1676037725
transform 1 0 49404 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_533
timestamp 1676037725
transform 1 0 50140 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_554
timestamp 1676037725
transform 1 0 52072 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_561
timestamp 1676037725
transform 1 0 52716 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_569
timestamp 1676037725
transform 1 0 53452 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_573
timestamp 1676037725
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_585
timestamp 1676037725
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_597
timestamp 1676037725
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_609
timestamp 1676037725
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_615
timestamp 1676037725
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_617
timestamp 1676037725
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_629
timestamp 1676037725
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_641
timestamp 1676037725
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_653
timestamp 1676037725
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_665
timestamp 1676037725
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_671
timestamp 1676037725
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_673
timestamp 1676037725
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_685
timestamp 1676037725
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_697
timestamp 1676037725
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_709
timestamp 1676037725
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_721
timestamp 1676037725
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_727
timestamp 1676037725
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_729
timestamp 1676037725
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_741
timestamp 1676037725
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_753
timestamp 1676037725
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_765
timestamp 1676037725
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_777
timestamp 1676037725
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_783
timestamp 1676037725
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_785
timestamp 1676037725
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_797
timestamp 1676037725
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_809
timestamp 1676037725
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_821
timestamp 1676037725
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_833
timestamp 1676037725
transform 1 0 77740 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_839
timestamp 1676037725
transform 1 0 78292 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_841
timestamp 1676037725
transform 1 0 78476 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_853
timestamp 1676037725
transform 1 0 79580 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_857
timestamp 1676037725
transform 1 0 79948 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_869
timestamp 1676037725
transform 1 0 81052 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_894
timestamp 1676037725
transform 1 0 83352 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_897
timestamp 1676037725
transform 1 0 83628 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_901
timestamp 1676037725
transform 1 0 83996 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_905
timestamp 1676037725
transform 1 0 84364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_930
timestamp 1676037725
transform 1 0 86664 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_938
timestamp 1676037725
transform 1 0 87400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_942
timestamp 1676037725
transform 1 0 87768 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_946
timestamp 1676037725
transform 1 0 88136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_950
timestamp 1676037725
transform 1 0 88504 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_953
timestamp 1676037725
transform 1 0 88780 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_958
timestamp 1676037725
transform 1 0 89240 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_981
timestamp 1676037725
transform 1 0 91356 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1006
timestamp 1676037725
transform 1 0 93656 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1009
timestamp 1676037725
transform 1 0 93932 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1013
timestamp 1676037725
transform 1 0 94300 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1017
timestamp 1676037725
transform 1 0 94668 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1021
timestamp 1676037725
transform 1 0 95036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1033
timestamp 1676037725
transform 1 0 96140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1045
timestamp 1676037725
transform 1 0 97244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_1057
timestamp 1676037725
transform 1 0 98348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1063
timestamp 1676037725
transform 1 0 98900 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1065
timestamp 1676037725
transform 1 0 99084 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_1077
timestamp 1676037725
transform 1 0 100188 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1085
timestamp 1676037725
transform 1 0 100924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1089
timestamp 1676037725
transform 1 0 101292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1101
timestamp 1676037725
transform 1 0 102396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_1113
timestamp 1676037725
transform 1 0 103500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1119
timestamp 1676037725
transform 1 0 104052 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1121
timestamp 1676037725
transform 1 0 104236 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1133
timestamp 1676037725
transform 1 0 105340 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1139
timestamp 1676037725
transform 1 0 105892 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1162
timestamp 1676037725
transform 1 0 108008 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_1166
timestamp 1676037725
transform 1 0 108376 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1174
timestamp 1676037725
transform 1 0 109112 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1177
timestamp 1676037725
transform 1 0 109388 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_1189
timestamp 1676037725
transform 1 0 110492 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1197
timestamp 1676037725
transform 1 0 111228 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1201
timestamp 1676037725
transform 1 0 111596 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1224
timestamp 1676037725
transform 1 0 113712 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1230
timestamp 1676037725
transform 1 0 114264 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1233
timestamp 1676037725
transform 1 0 114540 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1237
timestamp 1676037725
transform 1 0 114908 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1260
timestamp 1676037725
transform 1 0 117024 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_1285
timestamp 1676037725
transform 1 0 119324 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1289
timestamp 1676037725
transform 1 0 119692 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1314
timestamp 1676037725
transform 1 0 121992 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1320
timestamp 1676037725
transform 1 0 122544 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1332
timestamp 1676037725
transform 1 0 123648 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1345
timestamp 1676037725
transform 1 0 124844 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1357
timestamp 1676037725
transform 1 0 125948 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1369
timestamp 1676037725
transform 1 0 127052 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1381
timestamp 1676037725
transform 1 0 128156 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_1393
timestamp 1676037725
transform 1 0 129260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1399
timestamp 1676037725
transform 1 0 129812 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1401
timestamp 1676037725
transform 1 0 129996 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1413
timestamp 1676037725
transform 1 0 131100 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1425
timestamp 1676037725
transform 1 0 132204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1437
timestamp 1676037725
transform 1 0 133308 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_1449
timestamp 1676037725
transform 1 0 134412 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1455
timestamp 1676037725
transform 1 0 134964 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1457
timestamp 1676037725
transform 1 0 135148 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1469
timestamp 1676037725
transform 1 0 136252 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1481
timestamp 1676037725
transform 1 0 137356 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1493
timestamp 1676037725
transform 1 0 138460 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_1505
timestamp 1676037725
transform 1 0 139564 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1511
timestamp 1676037725
transform 1 0 140116 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1513
timestamp 1676037725
transform 1 0 140300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1525
timestamp 1676037725
transform 1 0 141404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1537
timestamp 1676037725
transform 1 0 142508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1549
timestamp 1676037725
transform 1 0 143612 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_1561
timestamp 1676037725
transform 1 0 144716 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1567
timestamp 1676037725
transform 1 0 145268 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1569
timestamp 1676037725
transform 1 0 145452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1581
timestamp 1676037725
transform 1 0 146556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1593
timestamp 1676037725
transform 1 0 147660 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1605
timestamp 1676037725
transform 1 0 148764 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_1617
timestamp 1676037725
transform 1 0 149868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1622
timestamp 1676037725
transform 1 0 150328 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1646
timestamp 1676037725
transform 1 0 152536 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1650
timestamp 1676037725
transform 1 0 152904 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_1673
timestamp 1676037725
transform 1 0 155020 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1678
timestamp 1676037725
transform 1 0 155480 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1681
timestamp 1676037725
transform 1 0 155756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_1693
timestamp 1676037725
transform 1 0 156860 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1701
timestamp 1676037725
transform 1 0 157596 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1704
timestamp 1676037725
transform 1 0 157872 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1729
timestamp 1676037725
transform 1 0 160172 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_1733
timestamp 1676037725
transform 1 0 160540 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1737
timestamp 1676037725
transform 1 0 160908 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_1741
timestamp 1676037725
transform 1 0 161276 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1746
timestamp 1676037725
transform 1 0 161736 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1752
timestamp 1676037725
transform 1 0 162288 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1764
timestamp 1676037725
transform 1 0 163392 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1776
timestamp 1676037725
transform 1 0 164496 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_1788
timestamp 1676037725
transform 1 0 165600 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1793
timestamp 1676037725
transform 1 0 166060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1805
timestamp 1676037725
transform 1 0 167164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1817
timestamp 1676037725
transform 1 0 168268 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1829
timestamp 1676037725
transform 1 0 169372 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_1841
timestamp 1676037725
transform 1 0 170476 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1847
timestamp 1676037725
transform 1 0 171028 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1849
timestamp 1676037725
transform 1 0 171212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1861
timestamp 1676037725
transform 1 0 172316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1873
timestamp 1676037725
transform 1 0 173420 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1885
timestamp 1676037725
transform 1 0 174524 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_1897
timestamp 1676037725
transform 1 0 175628 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1903
timestamp 1676037725
transform 1 0 176180 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1905
timestamp 1676037725
transform 1 0 176364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1917
timestamp 1676037725
transform 1 0 177468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1929
timestamp 1676037725
transform 1 0 178572 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1941
timestamp 1676037725
transform 1 0 179676 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_1953
timestamp 1676037725
transform 1 0 180780 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_1959
timestamp 1676037725
transform 1 0 181332 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_1961
timestamp 1676037725
transform 1 0 181516 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1976
timestamp 1676037725
transform 1 0 182896 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_1988
timestamp 1676037725
transform 1 0 184000 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2000
timestamp 1676037725
transform 1 0 185104 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2012
timestamp 1676037725
transform 1 0 186208 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2017
timestamp 1676037725
transform 1 0 186668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2029
timestamp 1676037725
transform 1 0 187772 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2035
timestamp 1676037725
transform 1 0 188324 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2038
timestamp 1676037725
transform 1 0 188600 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2047
timestamp 1676037725
transform 1 0 189428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2059
timestamp 1676037725
transform 1 0 190532 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2071
timestamp 1676037725
transform 1 0 191636 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2073
timestamp 1676037725
transform 1 0 191820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2085
timestamp 1676037725
transform 1 0 192924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2097
timestamp 1676037725
transform 1 0 194028 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2109
timestamp 1676037725
transform 1 0 195132 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2121
timestamp 1676037725
transform 1 0 196236 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2127
timestamp 1676037725
transform 1 0 196788 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2129
timestamp 1676037725
transform 1 0 196972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2141
timestamp 1676037725
transform 1 0 198076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2153
timestamp 1676037725
transform 1 0 199180 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2165
timestamp 1676037725
transform 1 0 200284 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2177
timestamp 1676037725
transform 1 0 201388 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2183
timestamp 1676037725
transform 1 0 201940 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2185
timestamp 1676037725
transform 1 0 202124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2197
timestamp 1676037725
transform 1 0 203228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2209
timestamp 1676037725
transform 1 0 204332 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2221
timestamp 1676037725
transform 1 0 205436 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2233
timestamp 1676037725
transform 1 0 206540 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2239
timestamp 1676037725
transform 1 0 207092 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2241
timestamp 1676037725
transform 1 0 207276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2253
timestamp 1676037725
transform 1 0 208380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2265
timestamp 1676037725
transform 1 0 209484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2277
timestamp 1676037725
transform 1 0 210588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2289
timestamp 1676037725
transform 1 0 211692 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2295
timestamp 1676037725
transform 1 0 212244 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2297
timestamp 1676037725
transform 1 0 212428 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2309
timestamp 1676037725
transform 1 0 213532 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2313
timestamp 1676037725
transform 1 0 213900 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2335
timestamp 1676037725
transform 1 0 215924 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2347
timestamp 1676037725
transform 1 0 217028 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2351
timestamp 1676037725
transform 1 0 217396 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2353
timestamp 1676037725
transform 1 0 217580 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2361
timestamp 1676037725
transform 1 0 218316 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2365
timestamp 1676037725
transform 1 0 218684 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2369
timestamp 1676037725
transform 1 0 219052 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2392
timestamp 1676037725
transform 1 0 221168 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2396
timestamp 1676037725
transform 1 0 221536 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2400
timestamp 1676037725
transform 1 0 221904 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2406
timestamp 1676037725
transform 1 0 222456 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2409
timestamp 1676037725
transform 1 0 222732 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2431
timestamp 1676037725
transform 1 0 224756 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2435
timestamp 1676037725
transform 1 0 225124 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2439
timestamp 1676037725
transform 1 0 225492 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2462
timestamp 1676037725
transform 1 0 227608 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2465
timestamp 1676037725
transform 1 0 227884 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2485
timestamp 1676037725
transform 1 0 229724 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2494
timestamp 1676037725
transform 1 0 230552 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2505
timestamp 1676037725
transform 1 0 231564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_2517
timestamp 1676037725
transform 1 0 232668 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2521
timestamp 1676037725
transform 1 0 233036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2533
timestamp 1676037725
transform 1 0 234140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2545
timestamp 1676037725
transform 1 0 235244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2557
timestamp 1676037725
transform 1 0 236348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2569
timestamp 1676037725
transform 1 0 237452 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2575
timestamp 1676037725
transform 1 0 238004 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2577
timestamp 1676037725
transform 1 0 238188 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2585
timestamp 1676037725
transform 1 0 238924 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2595
timestamp 1676037725
transform 1 0 239844 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2603
timestamp 1676037725
transform 1 0 240580 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2615
timestamp 1676037725
transform 1 0 241684 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2619
timestamp 1676037725
transform 1 0 242052 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2623
timestamp 1676037725
transform 1 0 242420 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2627
timestamp 1676037725
transform 1 0 242788 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2631
timestamp 1676037725
transform 1 0 243156 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2633
timestamp 1676037725
transform 1 0 243340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2645
timestamp 1676037725
transform 1 0 244444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2657
timestamp 1676037725
transform 1 0 245548 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2669
timestamp 1676037725
transform 1 0 246652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2681
timestamp 1676037725
transform 1 0 247756 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2687
timestamp 1676037725
transform 1 0 248308 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2689
timestamp 1676037725
transform 1 0 248492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2701
timestamp 1676037725
transform 1 0 249596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2713
timestamp 1676037725
transform 1 0 250700 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2725
timestamp 1676037725
transform 1 0 251804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2737
timestamp 1676037725
transform 1 0 252908 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2743
timestamp 1676037725
transform 1 0 253460 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2745
timestamp 1676037725
transform 1 0 253644 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2757
timestamp 1676037725
transform 1 0 254748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2769
timestamp 1676037725
transform 1 0 255852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_2781
timestamp 1676037725
transform 1 0 256956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2793
timestamp 1676037725
transform 1 0 258060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2799
timestamp 1676037725
transform 1 0 258612 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_2801
timestamp 1676037725
transform 1 0 258796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2806
timestamp 1676037725
transform 1 0 259256 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2810
timestamp 1676037725
transform 1 0 259624 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_2814
timestamp 1676037725
transform 1 0 259992 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2826
timestamp 1676037725
transform 1 0 261096 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_2835
timestamp 1676037725
transform 1 0 261924 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2843
timestamp 1676037725
transform 1 0 262660 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2854
timestamp 1676037725
transform 1 0 263672 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2857
timestamp 1676037725
transform 1 0 263948 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_2868
timestamp 1676037725
transform 1 0 264960 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2876
timestamp 1676037725
transform 1 0 265696 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2883
timestamp 1676037725
transform 1 0 266340 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2892
timestamp 1676037725
transform 1 0 267168 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2900
timestamp 1676037725
transform 1 0 267904 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_2909
timestamp 1676037725
transform 1 0 268732 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_2913
timestamp 1676037725
transform 1 0 269100 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_2920
timestamp 1676037725
transform 1 0 269744 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_2929
timestamp 1676037725
transform 1 0 270572 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_2935
timestamp 1676037725
transform 1 0 271124 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1676037725
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 1676037725
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_441
timestamp 1676037725
transform 1 0 41676 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_450
timestamp 1676037725
transform 1 0 42504 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_454
timestamp 1676037725
transform 1 0 42872 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_474
timestamp 1676037725
transform 1 0 44712 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_489
timestamp 1676037725
transform 1 0 46092 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_510
timestamp 1676037725
transform 1 0 48024 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_522
timestamp 1676037725
transform 1 0 49128 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_530
timestamp 1676037725
transform 1 0 49864 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_533
timestamp 1676037725
transform 1 0 50140 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_553
timestamp 1676037725
transform 1 0 51980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_565
timestamp 1676037725
transform 1 0 53084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_577
timestamp 1676037725
transform 1 0 54188 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_585
timestamp 1676037725
transform 1 0 54924 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_589
timestamp 1676037725
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_601
timestamp 1676037725
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_613
timestamp 1676037725
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_625
timestamp 1676037725
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_637
timestamp 1676037725
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_643
timestamp 1676037725
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_645
timestamp 1676037725
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_657
timestamp 1676037725
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_669
timestamp 1676037725
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_681
timestamp 1676037725
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_693
timestamp 1676037725
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_699
timestamp 1676037725
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_701
timestamp 1676037725
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_713
timestamp 1676037725
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_725
timestamp 1676037725
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_737
timestamp 1676037725
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_749
timestamp 1676037725
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_755
timestamp 1676037725
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_757
timestamp 1676037725
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_769
timestamp 1676037725
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_781
timestamp 1676037725
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_793
timestamp 1676037725
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_805
timestamp 1676037725
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_811
timestamp 1676037725
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_813
timestamp 1676037725
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_825
timestamp 1676037725
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_837
timestamp 1676037725
transform 1 0 78108 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_845
timestamp 1676037725
transform 1 0 78844 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_853
timestamp 1676037725
transform 1 0 79580 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_865
timestamp 1676037725
transform 1 0 80684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_869
timestamp 1676037725
transform 1 0 81052 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_876
timestamp 1676037725
transform 1 0 81696 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_880
timestamp 1676037725
transform 1 0 82064 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_888
timestamp 1676037725
transform 1 0 82800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_892
timestamp 1676037725
transform 1 0 83168 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_915
timestamp 1676037725
transform 1 0 85284 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_919
timestamp 1676037725
transform 1 0 85652 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_923
timestamp 1676037725
transform 1 0 86020 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_925
timestamp 1676037725
transform 1 0 86204 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_929
timestamp 1676037725
transform 1 0 86572 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_946
timestamp 1676037725
transform 1 0 88136 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_958
timestamp 1676037725
transform 1 0 89240 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_970
timestamp 1676037725
transform 1 0 90344 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_978
timestamp 1676037725
transform 1 0 91080 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_981
timestamp 1676037725
transform 1 0 91356 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_993
timestamp 1676037725
transform 1 0 92460 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1016
timestamp 1676037725
transform 1 0 94576 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_1028
timestamp 1676037725
transform 1 0 95680 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1037
timestamp 1676037725
transform 1 0 96508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1049
timestamp 1676037725
transform 1 0 97612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1061
timestamp 1676037725
transform 1 0 98716 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1073
timestamp 1676037725
transform 1 0 99820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1077
timestamp 1676037725
transform 1 0 100188 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1080
timestamp 1676037725
transform 1 0 100464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1087
timestamp 1676037725
transform 1 0 101108 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1091
timestamp 1676037725
transform 1 0 101476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_1093
timestamp 1676037725
transform 1 0 101660 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1112
timestamp 1676037725
transform 1 0 103408 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1124
timestamp 1676037725
transform 1 0 104512 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1136
timestamp 1676037725
transform 1 0 105616 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1149
timestamp 1676037725
transform 1 0 106812 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1161
timestamp 1676037725
transform 1 0 107916 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1167
timestamp 1676037725
transform 1 0 108468 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1171
timestamp 1676037725
transform 1 0 108836 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1194
timestamp 1676037725
transform 1 0 110952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1198
timestamp 1676037725
transform 1 0 111320 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1202
timestamp 1676037725
transform 1 0 111688 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1205
timestamp 1676037725
transform 1 0 111964 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1209
timestamp 1676037725
transform 1 0 112332 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1212
timestamp 1676037725
transform 1 0 112608 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1216
timestamp 1676037725
transform 1 0 112976 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1239
timestamp 1676037725
transform 1 0 115092 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1243
timestamp 1676037725
transform 1 0 115460 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1247
timestamp 1676037725
transform 1 0 115828 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1259
timestamp 1676037725
transform 1 0 116932 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1261
timestamp 1676037725
transform 1 0 117116 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_1273
timestamp 1676037725
transform 1 0 118220 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1283
timestamp 1676037725
transform 1 0 119140 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1287
timestamp 1676037725
transform 1 0 119508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1291
timestamp 1676037725
transform 1 0 119876 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1314
timestamp 1676037725
transform 1 0 121992 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1317
timestamp 1676037725
transform 1 0 122268 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1321
timestamp 1676037725
transform 1 0 122636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1333
timestamp 1676037725
transform 1 0 123740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1345
timestamp 1676037725
transform 1 0 124844 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1352
timestamp 1676037725
transform 1 0 125488 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_1364
timestamp 1676037725
transform 1 0 126592 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1373
timestamp 1676037725
transform 1 0 127420 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1385
timestamp 1676037725
transform 1 0 128524 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1397
timestamp 1676037725
transform 1 0 129628 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1408
timestamp 1676037725
transform 1 0 130640 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_1420
timestamp 1676037725
transform 1 0 131744 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1429
timestamp 1676037725
transform 1 0 132572 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1441
timestamp 1676037725
transform 1 0 133676 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1453
timestamp 1676037725
transform 1 0 134780 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1465
timestamp 1676037725
transform 1 0 135884 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_1477
timestamp 1676037725
transform 1 0 136988 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1483
timestamp 1676037725
transform 1 0 137540 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1485
timestamp 1676037725
transform 1 0 137724 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1497
timestamp 1676037725
transform 1 0 138828 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1509
timestamp 1676037725
transform 1 0 139932 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1521
timestamp 1676037725
transform 1 0 141036 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_1533
timestamp 1676037725
transform 1 0 142140 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1539
timestamp 1676037725
transform 1 0 142692 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1541
timestamp 1676037725
transform 1 0 142876 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1564
timestamp 1676037725
transform 1 0 144992 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1576
timestamp 1676037725
transform 1 0 146096 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1588
timestamp 1676037725
transform 1 0 147200 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1594
timestamp 1676037725
transform 1 0 147752 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1597
timestamp 1676037725
transform 1 0 148028 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1620
timestamp 1676037725
transform 1 0 150144 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1624
timestamp 1676037725
transform 1 0 150512 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1628
timestamp 1676037725
transform 1 0 150880 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1642
timestamp 1676037725
transform 1 0 152168 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1646
timestamp 1676037725
transform 1 0 152536 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1650
timestamp 1676037725
transform 1 0 152904 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1653
timestamp 1676037725
transform 1 0 153180 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1676
timestamp 1676037725
transform 1 0 155296 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1701
timestamp 1676037725
transform 1 0 157596 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_1705
timestamp 1676037725
transform 1 0 157964 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1709
timestamp 1676037725
transform 1 0 158332 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1713
timestamp 1676037725
transform 1 0 158700 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1717
timestamp 1676037725
transform 1 0 159068 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_1721
timestamp 1676037725
transform 1 0 159436 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1727
timestamp 1676037725
transform 1 0 159988 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1730
timestamp 1676037725
transform 1 0 160264 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1734
timestamp 1676037725
transform 1 0 160632 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1738
timestamp 1676037725
transform 1 0 161000 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_1742
timestamp 1676037725
transform 1 0 161368 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1754
timestamp 1676037725
transform 1 0 162472 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_1760
timestamp 1676037725
transform 1 0 163024 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1765
timestamp 1676037725
transform 1 0 163484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1777
timestamp 1676037725
transform 1 0 164588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1789
timestamp 1676037725
transform 1 0 165692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1801
timestamp 1676037725
transform 1 0 166796 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_1813
timestamp 1676037725
transform 1 0 167900 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1819
timestamp 1676037725
transform 1 0 168452 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1821
timestamp 1676037725
transform 1 0 168636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1833
timestamp 1676037725
transform 1 0 169740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1845
timestamp 1676037725
transform 1 0 170844 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1857
timestamp 1676037725
transform 1 0 171948 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_1869
timestamp 1676037725
transform 1 0 173052 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1875
timestamp 1676037725
transform 1 0 173604 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1877
timestamp 1676037725
transform 1 0 173788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1889
timestamp 1676037725
transform 1 0 174892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1901
timestamp 1676037725
transform 1 0 175996 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1913
timestamp 1676037725
transform 1 0 177100 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_1925
timestamp 1676037725
transform 1 0 178204 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_1931
timestamp 1676037725
transform 1 0 178756 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1933
timestamp 1676037725
transform 1 0 178940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1945
timestamp 1676037725
transform 1 0 180044 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_1949
timestamp 1676037725
transform 1 0 180412 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_1956
timestamp 1676037725
transform 1 0 181056 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_1977
timestamp 1676037725
transform 1 0 182988 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_1985
timestamp 1676037725
transform 1 0 183724 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_1989
timestamp 1676037725
transform 1 0 184092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2001
timestamp 1676037725
transform 1 0 185196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2013
timestamp 1676037725
transform 1 0 186300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2025
timestamp 1676037725
transform 1 0 187404 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2037
timestamp 1676037725
transform 1 0 188508 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2043
timestamp 1676037725
transform 1 0 189060 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2045
timestamp 1676037725
transform 1 0 189244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2057
timestamp 1676037725
transform 1 0 190348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2069
timestamp 1676037725
transform 1 0 191452 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2081
timestamp 1676037725
transform 1 0 192556 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2093
timestamp 1676037725
transform 1 0 193660 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2099
timestamp 1676037725
transform 1 0 194212 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2101
timestamp 1676037725
transform 1 0 194396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2113
timestamp 1676037725
transform 1 0 195500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2125
timestamp 1676037725
transform 1 0 196604 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2137
timestamp 1676037725
transform 1 0 197708 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2149
timestamp 1676037725
transform 1 0 198812 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2155
timestamp 1676037725
transform 1 0 199364 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2157
timestamp 1676037725
transform 1 0 199548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2169
timestamp 1676037725
transform 1 0 200652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2181
timestamp 1676037725
transform 1 0 201756 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2193
timestamp 1676037725
transform 1 0 202860 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2205
timestamp 1676037725
transform 1 0 203964 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2211
timestamp 1676037725
transform 1 0 204516 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2213
timestamp 1676037725
transform 1 0 204700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2225
timestamp 1676037725
transform 1 0 205804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2237
timestamp 1676037725
transform 1 0 206908 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2249
timestamp 1676037725
transform 1 0 208012 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2261
timestamp 1676037725
transform 1 0 209116 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2267
timestamp 1676037725
transform 1 0 209668 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2269
timestamp 1676037725
transform 1 0 209852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2281
timestamp 1676037725
transform 1 0 210956 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2295
timestamp 1676037725
transform 1 0 212244 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2299
timestamp 1676037725
transform 1 0 212612 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2322
timestamp 1676037725
transform 1 0 214728 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2325
timestamp 1676037725
transform 1 0 215004 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2350
timestamp 1676037725
transform 1 0 217304 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2362
timestamp 1676037725
transform 1 0 218408 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2374
timestamp 1676037725
transform 1 0 219512 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_2381
timestamp 1676037725
transform 1 0 220156 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2389
timestamp 1676037725
transform 1 0 220892 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2393
timestamp 1676037725
transform 1 0 221260 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2397
timestamp 1676037725
transform 1 0 221628 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2420
timestamp 1676037725
transform 1 0 223744 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2424
timestamp 1676037725
transform 1 0 224112 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2428
timestamp 1676037725
transform 1 0 224480 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2434
timestamp 1676037725
transform 1 0 225032 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2437
timestamp 1676037725
transform 1 0 225308 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2460
timestamp 1676037725
transform 1 0 227424 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_2464
timestamp 1676037725
transform 1 0 227792 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2474
timestamp 1676037725
transform 1 0 228712 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2488
timestamp 1676037725
transform 1 0 230000 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2493
timestamp 1676037725
transform 1 0 230460 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2500
timestamp 1676037725
transform 1 0 231104 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2509
timestamp 1676037725
transform 1 0 231932 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2517
timestamp 1676037725
transform 1 0 232668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2529
timestamp 1676037725
transform 1 0 233772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2541
timestamp 1676037725
transform 1 0 234876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2547
timestamp 1676037725
transform 1 0 235428 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2549
timestamp 1676037725
transform 1 0 235612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2561
timestamp 1676037725
transform 1 0 236716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2573
timestamp 1676037725
transform 1 0 237820 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2585
timestamp 1676037725
transform 1 0 238924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2597
timestamp 1676037725
transform 1 0 240028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2603
timestamp 1676037725
transform 1 0 240580 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2605
timestamp 1676037725
transform 1 0 240764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2617
timestamp 1676037725
transform 1 0 241868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2629
timestamp 1676037725
transform 1 0 242972 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2641
timestamp 1676037725
transform 1 0 244076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2653
timestamp 1676037725
transform 1 0 245180 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2659
timestamp 1676037725
transform 1 0 245732 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2661
timestamp 1676037725
transform 1 0 245916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2673
timestamp 1676037725
transform 1 0 247020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2685
timestamp 1676037725
transform 1 0 248124 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2697
timestamp 1676037725
transform 1 0 249228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2709
timestamp 1676037725
transform 1 0 250332 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2715
timestamp 1676037725
transform 1 0 250884 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2717
timestamp 1676037725
transform 1 0 251068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2729
timestamp 1676037725
transform 1 0 252172 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2741
timestamp 1676037725
transform 1 0 253276 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2753
timestamp 1676037725
transform 1 0 254380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_2765
timestamp 1676037725
transform 1 0 255484 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2771
timestamp 1676037725
transform 1 0 256036 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2773
timestamp 1676037725
transform 1 0 256220 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_2785
timestamp 1676037725
transform 1 0 257324 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2797
timestamp 1676037725
transform 1 0 258428 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2801
timestamp 1676037725
transform 1 0 258796 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2811
timestamp 1676037725
transform 1 0 259716 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2824
timestamp 1676037725
transform 1 0 260912 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2829
timestamp 1676037725
transform 1 0 261372 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2840
timestamp 1676037725
transform 1 0 262384 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2853
timestamp 1676037725
transform 1 0 263580 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2866
timestamp 1676037725
transform 1 0 264776 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2875
timestamp 1676037725
transform 1 0 265604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2882
timestamp 1676037725
transform 1 0 266248 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_2885
timestamp 1676037725
transform 1 0 266524 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_2896
timestamp 1676037725
transform 1 0 267536 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2913
timestamp 1676037725
transform 1 0 269100 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2922
timestamp 1676037725
transform 1 0 269928 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_2931
timestamp 1676037725
transform 1 0 270756 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_2935
timestamp 1676037725
transform 1 0 271124 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1676037725
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 1676037725
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_429
timestamp 1676037725
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_441
timestamp 1676037725
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_469
timestamp 1676037725
transform 1 0 44252 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_473
timestamp 1676037725
transform 1 0 44620 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_493
timestamp 1676037725
transform 1 0 46460 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_497
timestamp 1676037725
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_503
timestamp 1676037725
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_517
timestamp 1676037725
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_529
timestamp 1676037725
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_541
timestamp 1676037725
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_553
timestamp 1676037725
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_559
timestamp 1676037725
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_561
timestamp 1676037725
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_573
timestamp 1676037725
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_585
timestamp 1676037725
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_597
timestamp 1676037725
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_609
timestamp 1676037725
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_615
timestamp 1676037725
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_617
timestamp 1676037725
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_629
timestamp 1676037725
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_641
timestamp 1676037725
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_653
timestamp 1676037725
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_665
timestamp 1676037725
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_671
timestamp 1676037725
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_673
timestamp 1676037725
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_685
timestamp 1676037725
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_697
timestamp 1676037725
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_709
timestamp 1676037725
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_721
timestamp 1676037725
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_727
timestamp 1676037725
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_729
timestamp 1676037725
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_741
timestamp 1676037725
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_753
timestamp 1676037725
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_765
timestamp 1676037725
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_777
timestamp 1676037725
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_783
timestamp 1676037725
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_785
timestamp 1676037725
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_797
timestamp 1676037725
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_809
timestamp 1676037725
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_821
timestamp 1676037725
transform 1 0 76636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_833
timestamp 1676037725
transform 1 0 77740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_839
timestamp 1676037725
transform 1 0 78292 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_841
timestamp 1676037725
transform 1 0 78476 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_854
timestamp 1676037725
transform 1 0 79672 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_866
timestamp 1676037725
transform 1 0 80776 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_878
timestamp 1676037725
transform 1 0 81880 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_890
timestamp 1676037725
transform 1 0 82984 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_897
timestamp 1676037725
transform 1 0 83628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_909
timestamp 1676037725
transform 1 0 84732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_921
timestamp 1676037725
transform 1 0 85836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_933
timestamp 1676037725
transform 1 0 86940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_945
timestamp 1676037725
transform 1 0 88044 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_951
timestamp 1676037725
transform 1 0 88596 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_953
timestamp 1676037725
transform 1 0 88780 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_965
timestamp 1676037725
transform 1 0 89884 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_973
timestamp 1676037725
transform 1 0 90620 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_977
timestamp 1676037725
transform 1 0 90988 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_981
timestamp 1676037725
transform 1 0 91356 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1004
timestamp 1676037725
transform 1 0 93472 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1009
timestamp 1676037725
transform 1 0 93932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1021
timestamp 1676037725
transform 1 0 95036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1033
timestamp 1676037725
transform 1 0 96140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1045
timestamp 1676037725
transform 1 0 97244 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_1057
timestamp 1676037725
transform 1 0 98348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1063
timestamp 1676037725
transform 1 0 98900 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_1065
timestamp 1676037725
transform 1 0 99084 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1071
timestamp 1676037725
transform 1 0 99636 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1079
timestamp 1676037725
transform 1 0 100372 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_1091
timestamp 1676037725
transform 1 0 101476 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1115
timestamp 1676037725
transform 1 0 103684 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1119
timestamp 1676037725
transform 1 0 104052 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1121
timestamp 1676037725
transform 1 0 104236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1133
timestamp 1676037725
transform 1 0 105340 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1145
timestamp 1676037725
transform 1 0 106444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1149
timestamp 1676037725
transform 1 0 106812 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1171
timestamp 1676037725
transform 1 0 108836 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1175
timestamp 1676037725
transform 1 0 109204 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1177
timestamp 1676037725
transform 1 0 109388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1189
timestamp 1676037725
transform 1 0 110492 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1214
timestamp 1676037725
transform 1 0 112792 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_1226
timestamp 1676037725
transform 1 0 113896 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1233
timestamp 1676037725
transform 1 0 114540 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1245
timestamp 1676037725
transform 1 0 115644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1257
timestamp 1676037725
transform 1 0 116748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1269
timestamp 1676037725
transform 1 0 117852 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_1281
timestamp 1676037725
transform 1 0 118956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_1286
timestamp 1676037725
transform 1 0 119416 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_1289
timestamp 1676037725
transform 1 0 119692 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1296
timestamp 1676037725
transform 1 0 120336 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1307
timestamp 1676037725
transform 1 0 121348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1319
timestamp 1676037725
transform 1 0 122452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1331
timestamp 1676037725
transform 1 0 123556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1343
timestamp 1676037725
transform 1 0 124660 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_1345
timestamp 1676037725
transform 1 0 124844 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1356
timestamp 1676037725
transform 1 0 125856 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1368
timestamp 1676037725
transform 1 0 126960 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1380
timestamp 1676037725
transform 1 0 128064 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_1392
timestamp 1676037725
transform 1 0 129168 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_1401
timestamp 1676037725
transform 1 0 129996 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1409
timestamp 1676037725
transform 1 0 130732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1421
timestamp 1676037725
transform 1 0 131836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1433
timestamp 1676037725
transform 1 0 132940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_1445
timestamp 1676037725
transform 1 0 134044 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_1453
timestamp 1676037725
transform 1 0 134780 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1457
timestamp 1676037725
transform 1 0 135148 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1469
timestamp 1676037725
transform 1 0 136252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1481
timestamp 1676037725
transform 1 0 137356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1493
timestamp 1676037725
transform 1 0 138460 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_1505
timestamp 1676037725
transform 1 0 139564 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1511
timestamp 1676037725
transform 1 0 140116 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1513
timestamp 1676037725
transform 1 0 140300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1525
timestamp 1676037725
transform 1 0 141404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1537
timestamp 1676037725
transform 1 0 142508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1549
timestamp 1676037725
transform 1 0 143612 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_1561
timestamp 1676037725
transform 1 0 144716 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1567
timestamp 1676037725
transform 1 0 145268 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_1569
timestamp 1676037725
transform 1 0 145452 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_1577
timestamp 1676037725
transform 1 0 146188 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1601
timestamp 1676037725
transform 1 0 148396 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_1621
timestamp 1676037725
transform 1 0 150236 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_1625
timestamp 1676037725
transform 1 0 150604 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1648
timestamp 1676037725
transform 1 0 152720 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1660
timestamp 1676037725
transform 1 0 153824 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_1672
timestamp 1676037725
transform 1 0 154928 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_1681
timestamp 1676037725
transform 1 0 155756 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_1689
timestamp 1676037725
transform 1 0 156492 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1699
timestamp 1676037725
transform 1 0 157412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1711
timestamp 1676037725
transform 1 0 158516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1723
timestamp 1676037725
transform 1 0 159620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1735
timestamp 1676037725
transform 1 0 160724 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_1737
timestamp 1676037725
transform 1 0 160908 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1745
timestamp 1676037725
transform 1 0 161644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1757
timestamp 1676037725
transform 1 0 162748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1769
timestamp 1676037725
transform 1 0 163852 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_1781
timestamp 1676037725
transform 1 0 164956 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_1789
timestamp 1676037725
transform 1 0 165692 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1793
timestamp 1676037725
transform 1 0 166060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1805
timestamp 1676037725
transform 1 0 167164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1817
timestamp 1676037725
transform 1 0 168268 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1829
timestamp 1676037725
transform 1 0 169372 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_1841
timestamp 1676037725
transform 1 0 170476 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1847
timestamp 1676037725
transform 1 0 171028 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1849
timestamp 1676037725
transform 1 0 171212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1861
timestamp 1676037725
transform 1 0 172316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1873
timestamp 1676037725
transform 1 0 173420 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1885
timestamp 1676037725
transform 1 0 174524 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_1897
timestamp 1676037725
transform 1 0 175628 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1903
timestamp 1676037725
transform 1 0 176180 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1905
timestamp 1676037725
transform 1 0 176364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1917
timestamp 1676037725
transform 1 0 177468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1929
timestamp 1676037725
transform 1 0 178572 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1941
timestamp 1676037725
transform 1 0 179676 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_1953
timestamp 1676037725
transform 1 0 180780 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_1959
timestamp 1676037725
transform 1 0 181332 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_1961
timestamp 1676037725
transform 1 0 181516 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1973
timestamp 1676037725
transform 1 0 182620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1985
timestamp 1676037725
transform 1 0 183724 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_1997
timestamp 1676037725
transform 1 0 184828 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2009
timestamp 1676037725
transform 1 0 185932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2015
timestamp 1676037725
transform 1 0 186484 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2017
timestamp 1676037725
transform 1 0 186668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2029
timestamp 1676037725
transform 1 0 187772 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2041
timestamp 1676037725
transform 1 0 188876 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2047
timestamp 1676037725
transform 1 0 189428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2059
timestamp 1676037725
transform 1 0 190532 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2071
timestamp 1676037725
transform 1 0 191636 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2073
timestamp 1676037725
transform 1 0 191820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2085
timestamp 1676037725
transform 1 0 192924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2097
timestamp 1676037725
transform 1 0 194028 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2109
timestamp 1676037725
transform 1 0 195132 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2121
timestamp 1676037725
transform 1 0 196236 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2127
timestamp 1676037725
transform 1 0 196788 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2129
timestamp 1676037725
transform 1 0 196972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2141
timestamp 1676037725
transform 1 0 198076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2153
timestamp 1676037725
transform 1 0 199180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2165
timestamp 1676037725
transform 1 0 200284 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2177
timestamp 1676037725
transform 1 0 201388 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2183
timestamp 1676037725
transform 1 0 201940 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2185
timestamp 1676037725
transform 1 0 202124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2197
timestamp 1676037725
transform 1 0 203228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2209
timestamp 1676037725
transform 1 0 204332 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2221
timestamp 1676037725
transform 1 0 205436 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2233
timestamp 1676037725
transform 1 0 206540 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2239
timestamp 1676037725
transform 1 0 207092 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_2241
timestamp 1676037725
transform 1 0 207276 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2265
timestamp 1676037725
transform 1 0 209484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2277
timestamp 1676037725
transform 1 0 210588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2289
timestamp 1676037725
transform 1 0 211692 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2295
timestamp 1676037725
transform 1 0 212244 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2297
timestamp 1676037725
transform 1 0 212428 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2309
timestamp 1676037725
transform 1 0 213532 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2315
timestamp 1676037725
transform 1 0 214084 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2337
timestamp 1676037725
transform 1 0 216108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_2349
timestamp 1676037725
transform 1 0 217212 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2353
timestamp 1676037725
transform 1 0 217580 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2376
timestamp 1676037725
transform 1 0 219696 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2380
timestamp 1676037725
transform 1 0 220064 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2403
timestamp 1676037725
transform 1 0 222180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2407
timestamp 1676037725
transform 1 0 222548 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2409
timestamp 1676037725
transform 1 0 222732 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2413
timestamp 1676037725
transform 1 0 223100 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2417
timestamp 1676037725
transform 1 0 223468 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2440
timestamp 1676037725
transform 1 0 225584 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2444
timestamp 1676037725
transform 1 0 225952 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_2456
timestamp 1676037725
transform 1 0 227056 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2465
timestamp 1676037725
transform 1 0 227884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2477
timestamp 1676037725
transform 1 0 228988 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2495
timestamp 1676037725
transform 1 0 230644 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_2510
timestamp 1676037725
transform 1 0 232024 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2518
timestamp 1676037725
transform 1 0 232760 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2521
timestamp 1676037725
transform 1 0 233036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2533
timestamp 1676037725
transform 1 0 234140 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_2545
timestamp 1676037725
transform 1 0 235244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2553
timestamp 1676037725
transform 1 0 235980 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2563
timestamp 1676037725
transform 1 0 236900 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2575
timestamp 1676037725
transform 1 0 238004 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2577
timestamp 1676037725
transform 1 0 238188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2589
timestamp 1676037725
transform 1 0 239292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2601
timestamp 1676037725
transform 1 0 240396 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2613
timestamp 1676037725
transform 1 0 241500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2625
timestamp 1676037725
transform 1 0 242604 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2631
timestamp 1676037725
transform 1 0 243156 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2633
timestamp 1676037725
transform 1 0 243340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2645
timestamp 1676037725
transform 1 0 244444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2657
timestamp 1676037725
transform 1 0 245548 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2669
timestamp 1676037725
transform 1 0 246652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2681
timestamp 1676037725
transform 1 0 247756 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2687
timestamp 1676037725
transform 1 0 248308 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2689
timestamp 1676037725
transform 1 0 248492 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2701
timestamp 1676037725
transform 1 0 249596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2713
timestamp 1676037725
transform 1 0 250700 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2725
timestamp 1676037725
transform 1 0 251804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2737
timestamp 1676037725
transform 1 0 252908 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2743
timestamp 1676037725
transform 1 0 253460 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2745
timestamp 1676037725
transform 1 0 253644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2757
timestamp 1676037725
transform 1 0 254748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2769
timestamp 1676037725
transform 1 0 255852 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2781
timestamp 1676037725
transform 1 0 256956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2793
timestamp 1676037725
transform 1 0 258060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2799
timestamp 1676037725
transform 1 0 258612 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2801
timestamp 1676037725
transform 1 0 258796 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_2813
timestamp 1676037725
transform 1 0 259900 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2825
timestamp 1676037725
transform 1 0 261004 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2835
timestamp 1676037725
transform 1 0 261924 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_2844
timestamp 1676037725
transform 1 0 262752 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2850
timestamp 1676037725
transform 1 0 263304 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2854
timestamp 1676037725
transform 1 0 263672 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2857
timestamp 1676037725
transform 1 0 263948 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2868
timestamp 1676037725
transform 1 0 264960 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2881
timestamp 1676037725
transform 1 0 266156 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2894
timestamp 1676037725
transform 1 0 267352 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2907
timestamp 1676037725
transform 1 0 268548 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_2911
timestamp 1676037725
transform 1 0 268916 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_2913
timestamp 1676037725
transform 1 0 269100 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_2924
timestamp 1676037725
transform 1 0 270112 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_2933
timestamp 1676037725
transform 1 0 270940 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1676037725
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1676037725
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1676037725
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_270
timestamp 1676037725
transform 1 0 25944 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_280
timestamp 1676037725
transform 1 0 26864 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_292
timestamp 1676037725
transform 1 0 27968 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_304
timestamp 1676037725
transform 1 0 29072 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1676037725
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_401
timestamp 1676037725
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_413
timestamp 1676037725
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_469
timestamp 1676037725
transform 1 0 44252 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_473
timestamp 1676037725
transform 1 0 44620 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_489
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_501
timestamp 1676037725
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_513
timestamp 1676037725
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_531
timestamp 1676037725
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_533
timestamp 1676037725
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_545
timestamp 1676037725
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_557
timestamp 1676037725
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_569
timestamp 1676037725
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_581
timestamp 1676037725
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_587
timestamp 1676037725
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_589
timestamp 1676037725
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_601
timestamp 1676037725
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_613
timestamp 1676037725
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_625
timestamp 1676037725
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_637
timestamp 1676037725
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_643
timestamp 1676037725
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_645
timestamp 1676037725
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_657
timestamp 1676037725
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_669
timestamp 1676037725
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_681
timestamp 1676037725
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_693
timestamp 1676037725
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_699
timestamp 1676037725
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_701
timestamp 1676037725
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_713
timestamp 1676037725
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_725
timestamp 1676037725
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_737
timestamp 1676037725
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_749
timestamp 1676037725
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_755
timestamp 1676037725
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_757
timestamp 1676037725
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_769
timestamp 1676037725
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_781
timestamp 1676037725
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_793
timestamp 1676037725
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_805
timestamp 1676037725
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_811
timestamp 1676037725
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_813
timestamp 1676037725
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_825
timestamp 1676037725
transform 1 0 77004 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_837
timestamp 1676037725
transform 1 0 78108 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_845
timestamp 1676037725
transform 1 0 78844 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_852
timestamp 1676037725
transform 1 0 79488 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_864
timestamp 1676037725
transform 1 0 80592 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_869
timestamp 1676037725
transform 1 0 81052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_881
timestamp 1676037725
transform 1 0 82156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_893
timestamp 1676037725
transform 1 0 83260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_905
timestamp 1676037725
transform 1 0 84364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_917
timestamp 1676037725
transform 1 0 85468 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_923
timestamp 1676037725
transform 1 0 86020 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_925
timestamp 1676037725
transform 1 0 86204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_937
timestamp 1676037725
transform 1 0 87308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_949
timestamp 1676037725
transform 1 0 88412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_961
timestamp 1676037725
transform 1 0 89516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_973
timestamp 1676037725
transform 1 0 90620 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_979
timestamp 1676037725
transform 1 0 91172 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_981
timestamp 1676037725
transform 1 0 91356 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_993
timestamp 1676037725
transform 1 0 92460 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1012
timestamp 1676037725
transform 1 0 94208 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1024
timestamp 1676037725
transform 1 0 95312 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1037
timestamp 1676037725
transform 1 0 96508 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_1049
timestamp 1676037725
transform 1 0 97612 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_1057
timestamp 1676037725
transform 1 0 98348 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1062
timestamp 1676037725
transform 1 0 98808 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1066
timestamp 1676037725
transform 1 0 99176 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_1089
timestamp 1676037725
transform 1 0 101292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1093
timestamp 1676037725
transform 1 0 101660 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1097
timestamp 1676037725
transform 1 0 102028 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1107
timestamp 1676037725
transform 1 0 102948 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1119
timestamp 1676037725
transform 1 0 104052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1131
timestamp 1676037725
transform 1 0 105156 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1143
timestamp 1676037725
transform 1 0 106260 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1147
timestamp 1676037725
transform 1 0 106628 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_1149
timestamp 1676037725
transform 1 0 106812 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1157
timestamp 1676037725
transform 1 0 107548 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1161
timestamp 1676037725
transform 1 0 107916 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1184
timestamp 1676037725
transform 1 0 110032 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1188
timestamp 1676037725
transform 1 0 110400 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1200
timestamp 1676037725
transform 1 0 111504 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1205
timestamp 1676037725
transform 1 0 111964 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1209
timestamp 1676037725
transform 1 0 112332 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1231
timestamp 1676037725
transform 1 0 114356 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1235
timestamp 1676037725
transform 1 0 114724 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1239
timestamp 1676037725
transform 1 0 115092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_1251
timestamp 1676037725
transform 1 0 116196 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1259
timestamp 1676037725
transform 1 0 116932 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1261
timestamp 1676037725
transform 1 0 117116 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1273
timestamp 1676037725
transform 1 0 118220 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1285
timestamp 1676037725
transform 1 0 119324 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1297
timestamp 1676037725
transform 1 0 120428 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1309
timestamp 1676037725
transform 1 0 121532 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1315
timestamp 1676037725
transform 1 0 122084 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1317
timestamp 1676037725
transform 1 0 122268 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1329
timestamp 1676037725
transform 1 0 123372 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1341
timestamp 1676037725
transform 1 0 124476 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1353
timestamp 1676037725
transform 1 0 125580 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1365
timestamp 1676037725
transform 1 0 126684 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1371
timestamp 1676037725
transform 1 0 127236 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1373
timestamp 1676037725
transform 1 0 127420 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1385
timestamp 1676037725
transform 1 0 128524 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1397
timestamp 1676037725
transform 1 0 129628 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1409
timestamp 1676037725
transform 1 0 130732 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1421
timestamp 1676037725
transform 1 0 131836 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1427
timestamp 1676037725
transform 1 0 132388 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1429
timestamp 1676037725
transform 1 0 132572 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1441
timestamp 1676037725
transform 1 0 133676 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1453
timestamp 1676037725
transform 1 0 134780 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1465
timestamp 1676037725
transform 1 0 135884 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1477
timestamp 1676037725
transform 1 0 136988 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1483
timestamp 1676037725
transform 1 0 137540 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1485
timestamp 1676037725
transform 1 0 137724 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1497
timestamp 1676037725
transform 1 0 138828 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1509
timestamp 1676037725
transform 1 0 139932 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1515
timestamp 1676037725
transform 1 0 140484 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1538
timestamp 1676037725
transform 1 0 142600 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1541
timestamp 1676037725
transform 1 0 142876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1553
timestamp 1676037725
transform 1 0 143980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_1565
timestamp 1676037725
transform 1 0 145084 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1594
timestamp 1676037725
transform 1 0 147752 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_1597
timestamp 1676037725
transform 1 0 148028 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1620
timestamp 1676037725
transform 1 0 150144 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1645
timestamp 1676037725
transform 1 0 152444 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1651
timestamp 1676037725
transform 1 0 152996 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1653
timestamp 1676037725
transform 1 0 153180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1665
timestamp 1676037725
transform 1 0 154284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1677
timestamp 1676037725
transform 1 0 155388 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1689
timestamp 1676037725
transform 1 0 156492 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1701
timestamp 1676037725
transform 1 0 157596 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1707
timestamp 1676037725
transform 1 0 158148 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1709
timestamp 1676037725
transform 1 0 158332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1721
timestamp 1676037725
transform 1 0 159436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1733
timestamp 1676037725
transform 1 0 160540 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1745
timestamp 1676037725
transform 1 0 161644 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1757
timestamp 1676037725
transform 1 0 162748 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1763
timestamp 1676037725
transform 1 0 163300 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1765
timestamp 1676037725
transform 1 0 163484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1777
timestamp 1676037725
transform 1 0 164588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1789
timestamp 1676037725
transform 1 0 165692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1801
timestamp 1676037725
transform 1 0 166796 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1813
timestamp 1676037725
transform 1 0 167900 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1819
timestamp 1676037725
transform 1 0 168452 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1821
timestamp 1676037725
transform 1 0 168636 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_1834
timestamp 1676037725
transform 1 0 169832 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1844
timestamp 1676037725
transform 1 0 170752 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1856
timestamp 1676037725
transform 1 0 171856 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_1868
timestamp 1676037725
transform 1 0 172960 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1877
timestamp 1676037725
transform 1 0 173788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1889
timestamp 1676037725
transform 1 0 174892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1901
timestamp 1676037725
transform 1 0 175996 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1913
timestamp 1676037725
transform 1 0 177100 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1925
timestamp 1676037725
transform 1 0 178204 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1931
timestamp 1676037725
transform 1 0 178756 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1933
timestamp 1676037725
transform 1 0 178940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1945
timestamp 1676037725
transform 1 0 180044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1957
timestamp 1676037725
transform 1 0 181148 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1969
timestamp 1676037725
transform 1 0 182252 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_1981
timestamp 1676037725
transform 1 0 183356 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_1987
timestamp 1676037725
transform 1 0 183908 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_1989
timestamp 1676037725
transform 1 0 184092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2001
timestamp 1676037725
transform 1 0 185196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2013
timestamp 1676037725
transform 1 0 186300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2025
timestamp 1676037725
transform 1 0 187404 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2037
timestamp 1676037725
transform 1 0 188508 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2043
timestamp 1676037725
transform 1 0 189060 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_2045
timestamp 1676037725
transform 1 0 189244 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2056
timestamp 1676037725
transform 1 0 190256 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2068
timestamp 1676037725
transform 1 0 191360 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2080
timestamp 1676037725
transform 1 0 192464 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_2092
timestamp 1676037725
transform 1 0 193568 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2101
timestamp 1676037725
transform 1 0 194396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2113
timestamp 1676037725
transform 1 0 195500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2125
timestamp 1676037725
transform 1 0 196604 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2137
timestamp 1676037725
transform 1 0 197708 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2149
timestamp 1676037725
transform 1 0 198812 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2155
timestamp 1676037725
transform 1 0 199364 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2157
timestamp 1676037725
transform 1 0 199548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2169
timestamp 1676037725
transform 1 0 200652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2181
timestamp 1676037725
transform 1 0 201756 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2193
timestamp 1676037725
transform 1 0 202860 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2205
timestamp 1676037725
transform 1 0 203964 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2211
timestamp 1676037725
transform 1 0 204516 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2213
timestamp 1676037725
transform 1 0 204700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2225
timestamp 1676037725
transform 1 0 205804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2237
timestamp 1676037725
transform 1 0 206908 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2249
timestamp 1676037725
transform 1 0 208012 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2261
timestamp 1676037725
transform 1 0 209116 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2267
timestamp 1676037725
transform 1 0 209668 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2269
timestamp 1676037725
transform 1 0 209852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2294
timestamp 1676037725
transform 1 0 212152 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2319
timestamp 1676037725
transform 1 0 214452 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2323
timestamp 1676037725
transform 1 0 214820 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_2325
timestamp 1676037725
transform 1 0 215004 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2330
timestamp 1676037725
transform 1 0 215464 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2353
timestamp 1676037725
transform 1 0 217580 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2378
timestamp 1676037725
transform 1 0 219880 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2402
timestamp 1676037725
transform 1 0 222088 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2406
timestamp 1676037725
transform 1 0 222456 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_2429
timestamp 1676037725
transform 1 0 224572 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2434
timestamp 1676037725
transform 1 0 225032 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2437
timestamp 1676037725
transform 1 0 225308 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2460
timestamp 1676037725
transform 1 0 227424 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2464
timestamp 1676037725
transform 1 0 227792 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2468
timestamp 1676037725
transform 1 0 228160 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_2480
timestamp 1676037725
transform 1 0 229264 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2490
timestamp 1676037725
transform 1 0 230184 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2493
timestamp 1676037725
transform 1 0 230460 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2497
timestamp 1676037725
transform 1 0 230828 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2510
timestamp 1676037725
transform 1 0 232024 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2522
timestamp 1676037725
transform 1 0 233128 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2534
timestamp 1676037725
transform 1 0 234232 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2546
timestamp 1676037725
transform 1 0 235336 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2558
timestamp 1676037725
transform 1 0 236440 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2562
timestamp 1676037725
transform 1 0 236808 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2569
timestamp 1676037725
transform 1 0 237452 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2581
timestamp 1676037725
transform 1 0 238556 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_2593
timestamp 1676037725
transform 1 0 239660 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_2601
timestamp 1676037725
transform 1 0 240396 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2605
timestamp 1676037725
transform 1 0 240764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2617
timestamp 1676037725
transform 1 0 241868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2629
timestamp 1676037725
transform 1 0 242972 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2641
timestamp 1676037725
transform 1 0 244076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2653
timestamp 1676037725
transform 1 0 245180 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2659
timestamp 1676037725
transform 1 0 245732 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2661
timestamp 1676037725
transform 1 0 245916 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2673
timestamp 1676037725
transform 1 0 247020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2685
timestamp 1676037725
transform 1 0 248124 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2697
timestamp 1676037725
transform 1 0 249228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2709
timestamp 1676037725
transform 1 0 250332 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2715
timestamp 1676037725
transform 1 0 250884 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2717
timestamp 1676037725
transform 1 0 251068 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2729
timestamp 1676037725
transform 1 0 252172 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2741
timestamp 1676037725
transform 1 0 253276 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2753
timestamp 1676037725
transform 1 0 254380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2765
timestamp 1676037725
transform 1 0 255484 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2771
timestamp 1676037725
transform 1 0 256036 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2773
timestamp 1676037725
transform 1 0 256220 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2785
timestamp 1676037725
transform 1 0 257324 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_2797
timestamp 1676037725
transform 1 0 258428 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2809
timestamp 1676037725
transform 1 0 259532 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2815
timestamp 1676037725
transform 1 0 260084 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2819
timestamp 1676037725
transform 1 0 260452 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_2826
timestamp 1676037725
transform 1 0 261096 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2829
timestamp 1676037725
transform 1 0 261372 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2835
timestamp 1676037725
transform 1 0 261924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2839
timestamp 1676037725
transform 1 0 262292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2846
timestamp 1676037725
transform 1 0 262936 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2854
timestamp 1676037725
transform 1 0 263672 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2862
timestamp 1676037725
transform 1 0 264408 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2870
timestamp 1676037725
transform 1 0 265144 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2878
timestamp 1676037725
transform 1 0 265880 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_2885
timestamp 1676037725
transform 1 0 266524 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_2891
timestamp 1676037725
transform 1 0 267076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2897
timestamp 1676037725
transform 1 0 267628 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2910
timestamp 1676037725
transform 1 0 268824 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_2924
timestamp 1676037725
transform 1 0 270112 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_2933
timestamp 1676037725
transform 1 0 270940 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_253
timestamp 1676037725
transform 1 0 24380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_258
timestamp 1676037725
transform 1 0 24840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_267
timestamp 1676037725
transform 1 0 25668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_276
timestamp 1676037725
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_289
timestamp 1676037725
transform 1 0 27692 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_294
timestamp 1676037725
transform 1 0 28152 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_306
timestamp 1676037725
transform 1 0 29256 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_318
timestamp 1676037725
transform 1 0 30360 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_330
timestamp 1676037725
transform 1 0 31464 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1676037725
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1676037725
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1676037725
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1676037725
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1676037725
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1676037725
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 1676037725
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_429
timestamp 1676037725
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 1676037725
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1676037725
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_454
timestamp 1676037725
transform 1 0 42872 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_458
timestamp 1676037725
transform 1 0 43240 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_470
timestamp 1676037725
transform 1 0 44344 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_482
timestamp 1676037725
transform 1 0 45448 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_494
timestamp 1676037725
transform 1 0 46552 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_502
timestamp 1676037725
transform 1 0 47288 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_517
timestamp 1676037725
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_529
timestamp 1676037725
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_541
timestamp 1676037725
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_553
timestamp 1676037725
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_559
timestamp 1676037725
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_561
timestamp 1676037725
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_573
timestamp 1676037725
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_585
timestamp 1676037725
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_597
timestamp 1676037725
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_609
timestamp 1676037725
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_615
timestamp 1676037725
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_617
timestamp 1676037725
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_629
timestamp 1676037725
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_641
timestamp 1676037725
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_653
timestamp 1676037725
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_665
timestamp 1676037725
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_671
timestamp 1676037725
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_673
timestamp 1676037725
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_685
timestamp 1676037725
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_697
timestamp 1676037725
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_709
timestamp 1676037725
transform 1 0 66332 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_717
timestamp 1676037725
transform 1 0 67068 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_723
timestamp 1676037725
transform 1 0 67620 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_727
timestamp 1676037725
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_729
timestamp 1676037725
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_741
timestamp 1676037725
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_753
timestamp 1676037725
transform 1 0 70380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_765
timestamp 1676037725
transform 1 0 71484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_777
timestamp 1676037725
transform 1 0 72588 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_783
timestamp 1676037725
transform 1 0 73140 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_785
timestamp 1676037725
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_797
timestamp 1676037725
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_809
timestamp 1676037725
transform 1 0 75532 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_821
timestamp 1676037725
transform 1 0 76636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_833
timestamp 1676037725
transform 1 0 77740 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_839
timestamp 1676037725
transform 1 0 78292 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_841
timestamp 1676037725
transform 1 0 78476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_853
timestamp 1676037725
transform 1 0 79580 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_865
timestamp 1676037725
transform 1 0 80684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_877
timestamp 1676037725
transform 1 0 81788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_889
timestamp 1676037725
transform 1 0 82892 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_895
timestamp 1676037725
transform 1 0 83444 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_897
timestamp 1676037725
transform 1 0 83628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_909
timestamp 1676037725
transform 1 0 84732 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_921
timestamp 1676037725
transform 1 0 85836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_933
timestamp 1676037725
transform 1 0 86940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_945
timestamp 1676037725
transform 1 0 88044 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_951
timestamp 1676037725
transform 1 0 88596 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_953
timestamp 1676037725
transform 1 0 88780 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_965
timestamp 1676037725
transform 1 0 89884 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_977
timestamp 1676037725
transform 1 0 90988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_989
timestamp 1676037725
transform 1 0 92092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1001
timestamp 1676037725
transform 1 0 93196 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1007
timestamp 1676037725
transform 1 0 93748 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1009
timestamp 1676037725
transform 1 0 93932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1021
timestamp 1676037725
transform 1 0 95036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1033
timestamp 1676037725
transform 1 0 96140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1045
timestamp 1676037725
transform 1 0 97244 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1057
timestamp 1676037725
transform 1 0 98348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1063
timestamp 1676037725
transform 1 0 98900 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_1065
timestamp 1676037725
transform 1 0 99084 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1073
timestamp 1676037725
transform 1 0 99820 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1078
timestamp 1676037725
transform 1 0 100280 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1090
timestamp 1676037725
transform 1 0 101384 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1102
timestamp 1676037725
transform 1 0 102488 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1114
timestamp 1676037725
transform 1 0 103592 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1121
timestamp 1676037725
transform 1 0 104236 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_1133
timestamp 1676037725
transform 1 0 105340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1143
timestamp 1676037725
transform 1 0 106260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1170
timestamp 1676037725
transform 1 0 108744 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1174
timestamp 1676037725
transform 1 0 109112 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1177
timestamp 1676037725
transform 1 0 109388 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1200
timestamp 1676037725
transform 1 0 111504 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1220
timestamp 1676037725
transform 1 0 113344 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1233
timestamp 1676037725
transform 1 0 114540 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1245
timestamp 1676037725
transform 1 0 115644 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1257
timestamp 1676037725
transform 1 0 116748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1269
timestamp 1676037725
transform 1 0 117852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1281
timestamp 1676037725
transform 1 0 118956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1287
timestamp 1676037725
transform 1 0 119508 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1289
timestamp 1676037725
transform 1 0 119692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_1301
timestamp 1676037725
transform 1 0 120796 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1308
timestamp 1676037725
transform 1 0 121440 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1320
timestamp 1676037725
transform 1 0 122544 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1332
timestamp 1676037725
transform 1 0 123648 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1345
timestamp 1676037725
transform 1 0 124844 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1357
timestamp 1676037725
transform 1 0 125948 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1369
timestamp 1676037725
transform 1 0 127052 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1381
timestamp 1676037725
transform 1 0 128156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1393
timestamp 1676037725
transform 1 0 129260 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1399
timestamp 1676037725
transform 1 0 129812 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1401
timestamp 1676037725
transform 1 0 129996 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1413
timestamp 1676037725
transform 1 0 131100 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1425
timestamp 1676037725
transform 1 0 132204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1437
timestamp 1676037725
transform 1 0 133308 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1449
timestamp 1676037725
transform 1 0 134412 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1455
timestamp 1676037725
transform 1 0 134964 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1457
timestamp 1676037725
transform 1 0 135148 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1469
timestamp 1676037725
transform 1 0 136252 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1481
timestamp 1676037725
transform 1 0 137356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1493
timestamp 1676037725
transform 1 0 138460 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1505
timestamp 1676037725
transform 1 0 139564 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1511
timestamp 1676037725
transform 1 0 140116 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1513
timestamp 1676037725
transform 1 0 140300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1525
timestamp 1676037725
transform 1 0 141404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1537
timestamp 1676037725
transform 1 0 142508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1549
timestamp 1676037725
transform 1 0 143612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1561
timestamp 1676037725
transform 1 0 144716 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1567
timestamp 1676037725
transform 1 0 145268 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1569
timestamp 1676037725
transform 1 0 145452 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1592
timestamp 1676037725
transform 1 0 147568 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1596
timestamp 1676037725
transform 1 0 147936 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1608
timestamp 1676037725
transform 1 0 149040 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_1620
timestamp 1676037725
transform 1 0 150144 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1625
timestamp 1676037725
transform 1 0 150604 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1629
timestamp 1676037725
transform 1 0 150972 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1652
timestamp 1676037725
transform 1 0 153088 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1656
timestamp 1676037725
transform 1 0 153456 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1668
timestamp 1676037725
transform 1 0 154560 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1681
timestamp 1676037725
transform 1 0 155756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1693
timestamp 1676037725
transform 1 0 156860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1705
timestamp 1676037725
transform 1 0 157964 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1717
timestamp 1676037725
transform 1 0 159068 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1729
timestamp 1676037725
transform 1 0 160172 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1735
timestamp 1676037725
transform 1 0 160724 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1737
timestamp 1676037725
transform 1 0 160908 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_1743
timestamp 1676037725
transform 1 0 161460 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_1751
timestamp 1676037725
transform 1 0 162196 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_1757
timestamp 1676037725
transform 1 0 162748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_1765
timestamp 1676037725
transform 1 0 163484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_1773
timestamp 1676037725
transform 1 0 164220 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_1781
timestamp 1676037725
transform 1 0 164956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_1789
timestamp 1676037725
transform 1 0 165692 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1793
timestamp 1676037725
transform 1 0 166060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1805
timestamp 1676037725
transform 1 0 167164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_1817
timestamp 1676037725
transform 1 0 168268 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1825
timestamp 1676037725
transform 1 0 169004 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1829
timestamp 1676037725
transform 1 0 169372 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1841
timestamp 1676037725
transform 1 0 170476 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1847
timestamp 1676037725
transform 1 0 171028 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1849
timestamp 1676037725
transform 1 0 171212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1861
timestamp 1676037725
transform 1 0 172316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1873
timestamp 1676037725
transform 1 0 173420 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1885
timestamp 1676037725
transform 1 0 174524 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1897
timestamp 1676037725
transform 1 0 175628 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1903
timestamp 1676037725
transform 1 0 176180 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1905
timestamp 1676037725
transform 1 0 176364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1917
timestamp 1676037725
transform 1 0 177468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1929
timestamp 1676037725
transform 1 0 178572 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1941
timestamp 1676037725
transform 1 0 179676 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_1953
timestamp 1676037725
transform 1 0 180780 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_1959
timestamp 1676037725
transform 1 0 181332 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1961
timestamp 1676037725
transform 1 0 181516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1973
timestamp 1676037725
transform 1 0 182620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1985
timestamp 1676037725
transform 1 0 183724 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_1997
timestamp 1676037725
transform 1 0 184828 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2009
timestamp 1676037725
transform 1 0 185932 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2015
timestamp 1676037725
transform 1 0 186484 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2017
timestamp 1676037725
transform 1 0 186668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2029
timestamp 1676037725
transform 1 0 187772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2041
timestamp 1676037725
transform 1 0 188876 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2053
timestamp 1676037725
transform 1 0 189980 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2065
timestamp 1676037725
transform 1 0 191084 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2071
timestamp 1676037725
transform 1 0 191636 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2073
timestamp 1676037725
transform 1 0 191820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2085
timestamp 1676037725
transform 1 0 192924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2097
timestamp 1676037725
transform 1 0 194028 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2109
timestamp 1676037725
transform 1 0 195132 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2121
timestamp 1676037725
transform 1 0 196236 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2127
timestamp 1676037725
transform 1 0 196788 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2129
timestamp 1676037725
transform 1 0 196972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2141
timestamp 1676037725
transform 1 0 198076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2153
timestamp 1676037725
transform 1 0 199180 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2165
timestamp 1676037725
transform 1 0 200284 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2177
timestamp 1676037725
transform 1 0 201388 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2183
timestamp 1676037725
transform 1 0 201940 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2185
timestamp 1676037725
transform 1 0 202124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2197
timestamp 1676037725
transform 1 0 203228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2209
timestamp 1676037725
transform 1 0 204332 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2221
timestamp 1676037725
transform 1 0 205436 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2233
timestamp 1676037725
transform 1 0 206540 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2239
timestamp 1676037725
transform 1 0 207092 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2241
timestamp 1676037725
transform 1 0 207276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2253
timestamp 1676037725
transform 1 0 208380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2265
timestamp 1676037725
transform 1 0 209484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2277
timestamp 1676037725
transform 1 0 210588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2289
timestamp 1676037725
transform 1 0 211692 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2295
timestamp 1676037725
transform 1 0 212244 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2297
timestamp 1676037725
transform 1 0 212428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2309
timestamp 1676037725
transform 1 0 213532 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2317
timestamp 1676037725
transform 1 0 214268 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2346
timestamp 1676037725
transform 1 0 216936 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2350
timestamp 1676037725
transform 1 0 217304 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2353
timestamp 1676037725
transform 1 0 217580 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2376
timestamp 1676037725
transform 1 0 219696 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2380
timestamp 1676037725
transform 1 0 220064 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2384
timestamp 1676037725
transform 1 0 220432 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2406
timestamp 1676037725
transform 1 0 222456 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2409
timestamp 1676037725
transform 1 0 222732 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2432
timestamp 1676037725
transform 1 0 224848 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2436
timestamp 1676037725
transform 1 0 225216 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2448
timestamp 1676037725
transform 1 0 226320 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2460
timestamp 1676037725
transform 1 0 227424 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2465
timestamp 1676037725
transform 1 0 227884 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2477
timestamp 1676037725
transform 1 0 228988 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2486
timestamp 1676037725
transform 1 0 229816 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2496
timestamp 1676037725
transform 1 0 230736 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2509
timestamp 1676037725
transform 1 0 231932 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_2517
timestamp 1676037725
transform 1 0 232668 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2521
timestamp 1676037725
transform 1 0 233036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2533
timestamp 1676037725
transform 1 0 234140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2550
timestamp 1676037725
transform 1 0 235704 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2563
timestamp 1676037725
transform 1 0 236900 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2572
timestamp 1676037725
transform 1 0 237728 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2577
timestamp 1676037725
transform 1 0 238188 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2584
timestamp 1676037725
transform 1 0 238832 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2588
timestamp 1676037725
transform 1 0 239200 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2600
timestamp 1676037725
transform 1 0 240304 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2612
timestamp 1676037725
transform 1 0 241408 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_2624
timestamp 1676037725
transform 1 0 242512 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2633
timestamp 1676037725
transform 1 0 243340 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2645
timestamp 1676037725
transform 1 0 244444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2657
timestamp 1676037725
transform 1 0 245548 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2669
timestamp 1676037725
transform 1 0 246652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2681
timestamp 1676037725
transform 1 0 247756 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2687
timestamp 1676037725
transform 1 0 248308 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2689
timestamp 1676037725
transform 1 0 248492 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2701
timestamp 1676037725
transform 1 0 249596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2713
timestamp 1676037725
transform 1 0 250700 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2725
timestamp 1676037725
transform 1 0 251804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2737
timestamp 1676037725
transform 1 0 252908 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2743
timestamp 1676037725
transform 1 0 253460 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2745
timestamp 1676037725
transform 1 0 253644 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2757
timestamp 1676037725
transform 1 0 254748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2769
timestamp 1676037725
transform 1 0 255852 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_2781
timestamp 1676037725
transform 1 0 256956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2793
timestamp 1676037725
transform 1 0 258060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2799
timestamp 1676037725
transform 1 0 258612 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_2801
timestamp 1676037725
transform 1 0 258796 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2809
timestamp 1676037725
transform 1 0 259532 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2813
timestamp 1676037725
transform 1 0 259900 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2820
timestamp 1676037725
transform 1 0 260544 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2827
timestamp 1676037725
transform 1 0 261188 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2835
timestamp 1676037725
transform 1 0 261924 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2843
timestamp 1676037725
transform 1 0 262660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2851
timestamp 1676037725
transform 1 0 263396 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2855
timestamp 1676037725
transform 1 0 263764 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2857
timestamp 1676037725
transform 1 0 263948 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2863
timestamp 1676037725
transform 1 0 264500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2870
timestamp 1676037725
transform 1 0 265144 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2879
timestamp 1676037725
transform 1 0 265972 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2888
timestamp 1676037725
transform 1 0 266800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_2897
timestamp 1676037725
transform 1 0 267628 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_2903
timestamp 1676037725
transform 1 0 268180 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2910
timestamp 1676037725
transform 1 0 268824 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2913
timestamp 1676037725
transform 1 0 269100 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_2920
timestamp 1676037725
transform 1 0 269744 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_2934
timestamp 1676037725
transform 1 0 271032 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1676037725
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1676037725
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_257
timestamp 1676037725
transform 1 0 24748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_263
timestamp 1676037725
transform 1 0 25300 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_267
timestamp 1676037725
transform 1 0 25668 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_271
timestamp 1676037725
transform 1 0 26036 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_274
timestamp 1676037725
transform 1 0 26312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_281
timestamp 1676037725
transform 1 0 26956 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_290
timestamp 1676037725
transform 1 0 27784 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_298
timestamp 1676037725
transform 1 0 28520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_306
timestamp 1676037725
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1676037725
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1676037725
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1676037725
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1676037725
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1676037725
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 1676037725
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_401
timestamp 1676037725
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_413
timestamp 1676037725
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 1676037725
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_445
timestamp 1676037725
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_457
timestamp 1676037725
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_469
timestamp 1676037725
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_475
timestamp 1676037725
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_489
timestamp 1676037725
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_501
timestamp 1676037725
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_513
timestamp 1676037725
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_525
timestamp 1676037725
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_531
timestamp 1676037725
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_533
timestamp 1676037725
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_545
timestamp 1676037725
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_557
timestamp 1676037725
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_569
timestamp 1676037725
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_581
timestamp 1676037725
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_587
timestamp 1676037725
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_589
timestamp 1676037725
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_601
timestamp 1676037725
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_613
timestamp 1676037725
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_625
timestamp 1676037725
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_637
timestamp 1676037725
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_643
timestamp 1676037725
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_645
timestamp 1676037725
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_657
timestamp 1676037725
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_669
timestamp 1676037725
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_681
timestamp 1676037725
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_693
timestamp 1676037725
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_699
timestamp 1676037725
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_701
timestamp 1676037725
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_713
timestamp 1676037725
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_725
timestamp 1676037725
transform 1 0 67804 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_737
timestamp 1676037725
transform 1 0 68908 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_749
timestamp 1676037725
transform 1 0 70012 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_755
timestamp 1676037725
transform 1 0 70564 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_757
timestamp 1676037725
transform 1 0 70748 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_769
timestamp 1676037725
transform 1 0 71852 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_781
timestamp 1676037725
transform 1 0 72956 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_793
timestamp 1676037725
transform 1 0 74060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_805
timestamp 1676037725
transform 1 0 75164 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_811
timestamp 1676037725
transform 1 0 75716 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_813
timestamp 1676037725
transform 1 0 75900 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_825
timestamp 1676037725
transform 1 0 77004 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_837
timestamp 1676037725
transform 1 0 78108 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_849
timestamp 1676037725
transform 1 0 79212 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_861
timestamp 1676037725
transform 1 0 80316 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_867
timestamp 1676037725
transform 1 0 80868 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_869
timestamp 1676037725
transform 1 0 81052 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_881
timestamp 1676037725
transform 1 0 82156 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_893
timestamp 1676037725
transform 1 0 83260 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_905
timestamp 1676037725
transform 1 0 84364 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_917
timestamp 1676037725
transform 1 0 85468 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_923
timestamp 1676037725
transform 1 0 86020 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_925
timestamp 1676037725
transform 1 0 86204 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_937
timestamp 1676037725
transform 1 0 87308 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_949
timestamp 1676037725
transform 1 0 88412 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_965
timestamp 1676037725
transform 1 0 89884 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_977
timestamp 1676037725
transform 1 0 90988 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_981
timestamp 1676037725
transform 1 0 91356 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_993
timestamp 1676037725
transform 1 0 92460 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_999
timestamp 1676037725
transform 1 0 93012 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1004
timestamp 1676037725
transform 1 0 93472 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1016
timestamp 1676037725
transform 1 0 94576 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_1028
timestamp 1676037725
transform 1 0 95680 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1037
timestamp 1676037725
transform 1 0 96508 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1049
timestamp 1676037725
transform 1 0 97612 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1061
timestamp 1676037725
transform 1 0 98716 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1067
timestamp 1676037725
transform 1 0 99268 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_1072
timestamp 1676037725
transform 1 0 99728 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1079
timestamp 1676037725
transform 1 0 100372 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1091
timestamp 1676037725
transform 1 0 101476 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1093
timestamp 1676037725
transform 1 0 101660 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_1105
timestamp 1676037725
transform 1 0 102764 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_1113
timestamp 1676037725
transform 1 0 103500 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_1118
timestamp 1676037725
transform 1 0 103960 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_1122
timestamp 1676037725
transform 1 0 104328 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_1145
timestamp 1676037725
transform 1 0 106444 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_1149
timestamp 1676037725
transform 1 0 106812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1157
timestamp 1676037725
transform 1 0 107548 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_1162
timestamp 1676037725
transform 1 0 108008 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1170
timestamp 1676037725
transform 1 0 108744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_1177
timestamp 1676037725
transform 1 0 109388 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1185
timestamp 1676037725
transform 1 0 110124 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1197
timestamp 1676037725
transform 1 0 111228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1203
timestamp 1676037725
transform 1 0 111780 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1205
timestamp 1676037725
transform 1 0 111964 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1217
timestamp 1676037725
transform 1 0 113068 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1229
timestamp 1676037725
transform 1 0 114172 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1241
timestamp 1676037725
transform 1 0 115276 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1253
timestamp 1676037725
transform 1 0 116380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1259
timestamp 1676037725
transform 1 0 116932 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1261
timestamp 1676037725
transform 1 0 117116 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1273
timestamp 1676037725
transform 1 0 118220 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1285
timestamp 1676037725
transform 1 0 119324 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1297
timestamp 1676037725
transform 1 0 120428 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1309
timestamp 1676037725
transform 1 0 121532 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1315
timestamp 1676037725
transform 1 0 122084 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1317
timestamp 1676037725
transform 1 0 122268 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1329
timestamp 1676037725
transform 1 0 123372 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1341
timestamp 1676037725
transform 1 0 124476 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1353
timestamp 1676037725
transform 1 0 125580 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1365
timestamp 1676037725
transform 1 0 126684 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1371
timestamp 1676037725
transform 1 0 127236 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1373
timestamp 1676037725
transform 1 0 127420 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1385
timestamp 1676037725
transform 1 0 128524 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1397
timestamp 1676037725
transform 1 0 129628 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1409
timestamp 1676037725
transform 1 0 130732 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1421
timestamp 1676037725
transform 1 0 131836 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1427
timestamp 1676037725
transform 1 0 132388 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_1429
timestamp 1676037725
transform 1 0 132572 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1436
timestamp 1676037725
transform 1 0 133216 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1448
timestamp 1676037725
transform 1 0 134320 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1460
timestamp 1676037725
transform 1 0 135424 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1472
timestamp 1676037725
transform 1 0 136528 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1485
timestamp 1676037725
transform 1 0 137724 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1497
timestamp 1676037725
transform 1 0 138828 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1509
timestamp 1676037725
transform 1 0 139932 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1521
timestamp 1676037725
transform 1 0 141036 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1533
timestamp 1676037725
transform 1 0 142140 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1539
timestamp 1676037725
transform 1 0 142692 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1541
timestamp 1676037725
transform 1 0 142876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1553
timestamp 1676037725
transform 1 0 143980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1565
timestamp 1676037725
transform 1 0 145084 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1577
timestamp 1676037725
transform 1 0 146188 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1589
timestamp 1676037725
transform 1 0 147292 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1595
timestamp 1676037725
transform 1 0 147844 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1597
timestamp 1676037725
transform 1 0 148028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1609
timestamp 1676037725
transform 1 0 149132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1621
timestamp 1676037725
transform 1 0 150236 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1633
timestamp 1676037725
transform 1 0 151340 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1645
timestamp 1676037725
transform 1 0 152444 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1651
timestamp 1676037725
transform 1 0 152996 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1653
timestamp 1676037725
transform 1 0 153180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1665
timestamp 1676037725
transform 1 0 154284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1677
timestamp 1676037725
transform 1 0 155388 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1689
timestamp 1676037725
transform 1 0 156492 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1701
timestamp 1676037725
transform 1 0 157596 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1707
timestamp 1676037725
transform 1 0 158148 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1709
timestamp 1676037725
transform 1 0 158332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1721
timestamp 1676037725
transform 1 0 159436 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1727
timestamp 1676037725
transform 1 0 159988 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_1732
timestamp 1676037725
transform 1 0 160448 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_1740
timestamp 1676037725
transform 1 0 161184 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_1747
timestamp 1676037725
transform 1 0 161828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_1755
timestamp 1676037725
transform 1 0 162564 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1763
timestamp 1676037725
transform 1 0 163300 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_1765
timestamp 1676037725
transform 1 0 163484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_1772
timestamp 1676037725
transform 1 0 164128 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_1781
timestamp 1676037725
transform 1 0 164956 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_1790
timestamp 1676037725
transform 1 0 165784 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_1798
timestamp 1676037725
transform 1 0 166520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_1806
timestamp 1676037725
transform 1 0 167256 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1814
timestamp 1676037725
transform 1 0 167992 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_1821
timestamp 1676037725
transform 1 0 168636 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_1827
timestamp 1676037725
transform 1 0 169188 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1834
timestamp 1676037725
transform 1 0 169832 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1846
timestamp 1676037725
transform 1 0 170936 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1858
timestamp 1676037725
transform 1 0 172040 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1870
timestamp 1676037725
transform 1 0 173144 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1877
timestamp 1676037725
transform 1 0 173788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1889
timestamp 1676037725
transform 1 0 174892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1901
timestamp 1676037725
transform 1 0 175996 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1913
timestamp 1676037725
transform 1 0 177100 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1925
timestamp 1676037725
transform 1 0 178204 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1931
timestamp 1676037725
transform 1 0 178756 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1933
timestamp 1676037725
transform 1 0 178940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1945
timestamp 1676037725
transform 1 0 180044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1957
timestamp 1676037725
transform 1 0 181148 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1969
timestamp 1676037725
transform 1 0 182252 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_1981
timestamp 1676037725
transform 1 0 183356 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_1987
timestamp 1676037725
transform 1 0 183908 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_1989
timestamp 1676037725
transform 1 0 184092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2001
timestamp 1676037725
transform 1 0 185196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2013
timestamp 1676037725
transform 1 0 186300 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2025
timestamp 1676037725
transform 1 0 187404 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2037
timestamp 1676037725
transform 1 0 188508 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2043
timestamp 1676037725
transform 1 0 189060 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2045
timestamp 1676037725
transform 1 0 189244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2057
timestamp 1676037725
transform 1 0 190348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2069
timestamp 1676037725
transform 1 0 191452 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2081
timestamp 1676037725
transform 1 0 192556 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2093
timestamp 1676037725
transform 1 0 193660 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2099
timestamp 1676037725
transform 1 0 194212 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2101
timestamp 1676037725
transform 1 0 194396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2113
timestamp 1676037725
transform 1 0 195500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2125
timestamp 1676037725
transform 1 0 196604 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2137
timestamp 1676037725
transform 1 0 197708 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2149
timestamp 1676037725
transform 1 0 198812 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2155
timestamp 1676037725
transform 1 0 199364 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2157
timestamp 1676037725
transform 1 0 199548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2169
timestamp 1676037725
transform 1 0 200652 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_2181
timestamp 1676037725
transform 1 0 201756 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_2189
timestamp 1676037725
transform 1 0 202492 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2195
timestamp 1676037725
transform 1 0 203044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2207
timestamp 1676037725
transform 1 0 204148 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2211
timestamp 1676037725
transform 1 0 204516 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2213
timestamp 1676037725
transform 1 0 204700 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2225
timestamp 1676037725
transform 1 0 205804 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2237
timestamp 1676037725
transform 1 0 206908 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2249
timestamp 1676037725
transform 1 0 208012 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2261
timestamp 1676037725
transform 1 0 209116 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2267
timestamp 1676037725
transform 1 0 209668 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2269
timestamp 1676037725
transform 1 0 209852 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2281
timestamp 1676037725
transform 1 0 210956 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2293
timestamp 1676037725
transform 1 0 212060 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2305
timestamp 1676037725
transform 1 0 213164 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2317
timestamp 1676037725
transform 1 0 214268 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2323
timestamp 1676037725
transform 1 0 214820 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_2325
timestamp 1676037725
transform 1 0 215004 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2333
timestamp 1676037725
transform 1 0 215740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2350
timestamp 1676037725
transform 1 0 217304 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2360
timestamp 1676037725
transform 1 0 218224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2368
timestamp 1676037725
transform 1 0 218960 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2376
timestamp 1676037725
transform 1 0 219696 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2381
timestamp 1676037725
transform 1 0 220156 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2393
timestamp 1676037725
transform 1 0 221260 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2405
timestamp 1676037725
transform 1 0 222364 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2417
timestamp 1676037725
transform 1 0 223468 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2429
timestamp 1676037725
transform 1 0 224572 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2435
timestamp 1676037725
transform 1 0 225124 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2437
timestamp 1676037725
transform 1 0 225308 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2449
timestamp 1676037725
transform 1 0 226412 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2461
timestamp 1676037725
transform 1 0 227516 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2473
timestamp 1676037725
transform 1 0 228620 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2485
timestamp 1676037725
transform 1 0 229724 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2491
timestamp 1676037725
transform 1 0 230276 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_2493
timestamp 1676037725
transform 1 0 230460 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2499
timestamp 1676037725
transform 1 0 231012 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2511
timestamp 1676037725
transform 1 0 232116 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2523
timestamp 1676037725
transform 1 0 233220 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2535
timestamp 1676037725
transform 1 0 234324 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2547
timestamp 1676037725
transform 1 0 235428 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_2549
timestamp 1676037725
transform 1 0 235612 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_2554
timestamp 1676037725
transform 1 0 236072 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2562
timestamp 1676037725
transform 1 0 236808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2568
timestamp 1676037725
transform 1 0 237360 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2577
timestamp 1676037725
transform 1 0 238188 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2589
timestamp 1676037725
transform 1 0 239292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_2601
timestamp 1676037725
transform 1 0 240396 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2605
timestamp 1676037725
transform 1 0 240764 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2617
timestamp 1676037725
transform 1 0 241868 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2629
timestamp 1676037725
transform 1 0 242972 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2641
timestamp 1676037725
transform 1 0 244076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2653
timestamp 1676037725
transform 1 0 245180 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2659
timestamp 1676037725
transform 1 0 245732 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2661
timestamp 1676037725
transform 1 0 245916 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2673
timestamp 1676037725
transform 1 0 247020 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2685
timestamp 1676037725
transform 1 0 248124 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2697
timestamp 1676037725
transform 1 0 249228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2709
timestamp 1676037725
transform 1 0 250332 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2715
timestamp 1676037725
transform 1 0 250884 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2717
timestamp 1676037725
transform 1 0 251068 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2729
timestamp 1676037725
transform 1 0 252172 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2741
timestamp 1676037725
transform 1 0 253276 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2753
timestamp 1676037725
transform 1 0 254380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2765
timestamp 1676037725
transform 1 0 255484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2771
timestamp 1676037725
transform 1 0 256036 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_2773
timestamp 1676037725
transform 1 0 256220 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_2785
timestamp 1676037725
transform 1 0 257324 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2797
timestamp 1676037725
transform 1 0 258428 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2805
timestamp 1676037725
transform 1 0 259164 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2809
timestamp 1676037725
transform 1 0 259532 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2813
timestamp 1676037725
transform 1 0 259900 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2821
timestamp 1676037725
transform 1 0 260636 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2827
timestamp 1676037725
transform 1 0 261188 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2829
timestamp 1676037725
transform 1 0 261372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2838
timestamp 1676037725
transform 1 0 262200 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2847
timestamp 1676037725
transform 1 0 263028 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2856
timestamp 1676037725
transform 1 0 263856 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2863
timestamp 1676037725
transform 1 0 264500 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2872
timestamp 1676037725
transform 1 0 265328 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_2881
timestamp 1676037725
transform 1 0 266156 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_2885
timestamp 1676037725
transform 1 0 266524 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_2891
timestamp 1676037725
transform 1 0 267076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2898
timestamp 1676037725
transform 1 0 267720 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2909
timestamp 1676037725
transform 1 0 268732 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_2920
timestamp 1676037725
transform 1 0 269744 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_2934
timestamp 1676037725
transform 1 0 271032 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_237
timestamp 1676037725
transform 1 0 22908 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_245
timestamp 1676037725
transform 1 0 23644 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_252
timestamp 1676037725
transform 1 0 24288 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_256
timestamp 1676037725
transform 1 0 24656 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_263
timestamp 1676037725
transform 1 0 25300 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_278
timestamp 1676037725
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_289
timestamp 1676037725
transform 1 0 27692 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_295
timestamp 1676037725
transform 1 0 28244 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_301
timestamp 1676037725
transform 1 0 28796 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_307
timestamp 1676037725
transform 1 0 29348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_312
timestamp 1676037725
transform 1 0 29808 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_316
timestamp 1676037725
transform 1 0 30176 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_321
timestamp 1676037725
transform 1 0 30636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_325
timestamp 1676037725
transform 1 0 31004 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_330
timestamp 1676037725
transform 1 0 31464 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_344
timestamp 1676037725
transform 1 0 32752 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_351
timestamp 1676037725
transform 1 0 33396 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_363
timestamp 1676037725
transform 1 0 34500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_375
timestamp 1676037725
transform 1 0 35604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_387
timestamp 1676037725
transform 1 0 36708 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 1676037725
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_417
timestamp 1676037725
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_429
timestamp 1676037725
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_441
timestamp 1676037725
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_447
timestamp 1676037725
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_473
timestamp 1676037725
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_485
timestamp 1676037725
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_497
timestamp 1676037725
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_503
timestamp 1676037725
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_517
timestamp 1676037725
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_529
timestamp 1676037725
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_541
timestamp 1676037725
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_553
timestamp 1676037725
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_559
timestamp 1676037725
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_561
timestamp 1676037725
transform 1 0 52716 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_569
timestamp 1676037725
transform 1 0 53452 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_577
timestamp 1676037725
transform 1 0 54188 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_585
timestamp 1676037725
transform 1 0 54924 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_593
timestamp 1676037725
transform 1 0 55660 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_601
timestamp 1676037725
transform 1 0 56396 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_605
timestamp 1676037725
transform 1 0 56764 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_610
timestamp 1676037725
transform 1 0 57224 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_617
timestamp 1676037725
transform 1 0 57868 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_627
timestamp 1676037725
transform 1 0 58788 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_635
timestamp 1676037725
transform 1 0 59524 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_640
timestamp 1676037725
transform 1 0 59984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_649
timestamp 1676037725
transform 1 0 60812 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_659
timestamp 1676037725
transform 1 0 61732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_667
timestamp 1676037725
transform 1 0 62468 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_671
timestamp 1676037725
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_673
timestamp 1676037725
transform 1 0 63020 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_683
timestamp 1676037725
transform 1 0 63940 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_687
timestamp 1676037725
transform 1 0 64308 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_692
timestamp 1676037725
transform 1 0 64768 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_696
timestamp 1676037725
transform 1 0 65136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_701
timestamp 1676037725
transform 1 0 65596 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_709
timestamp 1676037725
transform 1 0 66332 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_717
timestamp 1676037725
transform 1 0 67068 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_724
timestamp 1676037725
transform 1 0 67712 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_729
timestamp 1676037725
transform 1 0 68172 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_741
timestamp 1676037725
transform 1 0 69276 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_753
timestamp 1676037725
transform 1 0 70380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_761
timestamp 1676037725
transform 1 0 71116 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_773
timestamp 1676037725
transform 1 0 72220 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_781
timestamp 1676037725
transform 1 0 72956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_785
timestamp 1676037725
transform 1 0 73324 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_793
timestamp 1676037725
transform 1 0 74060 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_805
timestamp 1676037725
transform 1 0 75164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_817
timestamp 1676037725
transform 1 0 76268 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_829
timestamp 1676037725
transform 1 0 77372 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_837
timestamp 1676037725
transform 1 0 78108 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_841
timestamp 1676037725
transform 1 0 78476 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_849
timestamp 1676037725
transform 1 0 79212 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_861
timestamp 1676037725
transform 1 0 80316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_873
timestamp 1676037725
transform 1 0 81420 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_885
timestamp 1676037725
transform 1 0 82524 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_893
timestamp 1676037725
transform 1 0 83260 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_897
timestamp 1676037725
transform 1 0 83628 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_909
timestamp 1676037725
transform 1 0 84732 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_921
timestamp 1676037725
transform 1 0 85836 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_933
timestamp 1676037725
transform 1 0 86940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_945
timestamp 1676037725
transform 1 0 88044 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_951
timestamp 1676037725
transform 1 0 88596 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_957
timestamp 1676037725
transform 1 0 89148 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_961
timestamp 1676037725
transform 1 0 89516 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_968
timestamp 1676037725
transform 1 0 90160 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_980
timestamp 1676037725
transform 1 0 91264 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_988
timestamp 1676037725
transform 1 0 92000 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_996
timestamp 1676037725
transform 1 0 92736 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_1005
timestamp 1676037725
transform 1 0 93564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1009
timestamp 1676037725
transform 1 0 93932 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1013
timestamp 1676037725
transform 1 0 94300 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1018
timestamp 1676037725
transform 1 0 94760 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_1026
timestamp 1676037725
transform 1 0 95496 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1034
timestamp 1676037725
transform 1 0 96232 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1041
timestamp 1676037725
transform 1 0 96876 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_1049
timestamp 1676037725
transform 1 0 97612 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1057
timestamp 1676037725
transform 1 0 98348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1062
timestamp 1676037725
transform 1 0 98808 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_1065
timestamp 1676037725
transform 1 0 99084 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1078
timestamp 1676037725
transform 1 0 100280 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1086
timestamp 1676037725
transform 1 0 101016 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1098
timestamp 1676037725
transform 1 0 102120 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_1110
timestamp 1676037725
transform 1 0 103224 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1118
timestamp 1676037725
transform 1 0 103960 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1121
timestamp 1676037725
transform 1 0 104236 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1133
timestamp 1676037725
transform 1 0 105340 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1145
timestamp 1676037725
transform 1 0 106444 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1157
timestamp 1676037725
transform 1 0 107548 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1169
timestamp 1676037725
transform 1 0 108652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1175
timestamp 1676037725
transform 1 0 109204 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1177
timestamp 1676037725
transform 1 0 109388 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1189
timestamp 1676037725
transform 1 0 110492 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1201
timestamp 1676037725
transform 1 0 111596 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1213
timestamp 1676037725
transform 1 0 112700 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1225
timestamp 1676037725
transform 1 0 113804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1231
timestamp 1676037725
transform 1 0 114356 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1233
timestamp 1676037725
transform 1 0 114540 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1245
timestamp 1676037725
transform 1 0 115644 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1257
timestamp 1676037725
transform 1 0 116748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1269
timestamp 1676037725
transform 1 0 117852 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1281
timestamp 1676037725
transform 1 0 118956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1287
timestamp 1676037725
transform 1 0 119508 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1289
timestamp 1676037725
transform 1 0 119692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1301
timestamp 1676037725
transform 1 0 120796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1307
timestamp 1676037725
transform 1 0 121348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_1314
timestamp 1676037725
transform 1 0 121992 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_1322
timestamp 1676037725
transform 1 0 122728 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1329
timestamp 1676037725
transform 1 0 123372 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1337
timestamp 1676037725
transform 1 0 124108 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1343
timestamp 1676037725
transform 1 0 124660 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1345
timestamp 1676037725
transform 1 0 124844 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1355
timestamp 1676037725
transform 1 0 125764 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1363
timestamp 1676037725
transform 1 0 126500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1371
timestamp 1676037725
transform 1 0 127236 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_1380
timestamp 1676037725
transform 1 0 128064 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_1388
timestamp 1676037725
transform 1 0 128800 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1396
timestamp 1676037725
transform 1 0 129536 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1401
timestamp 1676037725
transform 1 0 129996 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1412
timestamp 1676037725
transform 1 0 131008 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1420
timestamp 1676037725
transform 1 0 131744 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1428
timestamp 1676037725
transform 1 0 132480 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1432
timestamp 1676037725
transform 1 0 132848 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_1438
timestamp 1676037725
transform 1 0 133400 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1451
timestamp 1676037725
transform 1 0 134596 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1455
timestamp 1676037725
transform 1 0 134964 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1457
timestamp 1676037725
transform 1 0 135148 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1469
timestamp 1676037725
transform 1 0 136252 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1481
timestamp 1676037725
transform 1 0 137356 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1493
timestamp 1676037725
transform 1 0 138460 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1505
timestamp 1676037725
transform 1 0 139564 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1511
timestamp 1676037725
transform 1 0 140116 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1513
timestamp 1676037725
transform 1 0 140300 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1525
timestamp 1676037725
transform 1 0 141404 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1537
timestamp 1676037725
transform 1 0 142508 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1549
timestamp 1676037725
transform 1 0 143612 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1561
timestamp 1676037725
transform 1 0 144716 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1567
timestamp 1676037725
transform 1 0 145268 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1569
timestamp 1676037725
transform 1 0 145452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1581
timestamp 1676037725
transform 1 0 146556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1593
timestamp 1676037725
transform 1 0 147660 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1605
timestamp 1676037725
transform 1 0 148764 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1617
timestamp 1676037725
transform 1 0 149868 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1623
timestamp 1676037725
transform 1 0 150420 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1625
timestamp 1676037725
transform 1 0 150604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1637
timestamp 1676037725
transform 1 0 151708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1649
timestamp 1676037725
transform 1 0 152812 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1661
timestamp 1676037725
transform 1 0 153916 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1673
timestamp 1676037725
transform 1 0 155020 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1679
timestamp 1676037725
transform 1 0 155572 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_1681
timestamp 1676037725
transform 1 0 155756 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_1694
timestamp 1676037725
transform 1 0 156952 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_1702
timestamp 1676037725
transform 1 0 157688 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1710
timestamp 1676037725
transform 1 0 158424 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1721
timestamp 1676037725
transform 1 0 159436 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1730
timestamp 1676037725
transform 1 0 160264 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1737
timestamp 1676037725
transform 1 0 160908 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1748
timestamp 1676037725
transform 1 0 161920 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1757
timestamp 1676037725
transform 1 0 162748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1761
timestamp 1676037725
transform 1 0 163116 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_1764
timestamp 1676037725
transform 1 0 163392 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1775
timestamp 1676037725
transform 1 0 164404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_1784
timestamp 1676037725
transform 1 0 165232 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1793
timestamp 1676037725
transform 1 0 166060 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1811
timestamp 1676037725
transform 1 0 167716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_1827
timestamp 1676037725
transform 1 0 169188 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1836
timestamp 1676037725
transform 1 0 170016 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1849
timestamp 1676037725
transform 1 0 171212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1861
timestamp 1676037725
transform 1 0 172316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1873
timestamp 1676037725
transform 1 0 173420 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1885
timestamp 1676037725
transform 1 0 174524 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1897
timestamp 1676037725
transform 1 0 175628 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1903
timestamp 1676037725
transform 1 0 176180 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1905
timestamp 1676037725
transform 1 0 176364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1917
timestamp 1676037725
transform 1 0 177468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1929
timestamp 1676037725
transform 1 0 178572 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1941
timestamp 1676037725
transform 1 0 179676 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1953
timestamp 1676037725
transform 1 0 180780 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1959
timestamp 1676037725
transform 1 0 181332 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1961
timestamp 1676037725
transform 1 0 181516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_1973
timestamp 1676037725
transform 1 0 182620 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_1979
timestamp 1676037725
transform 1 0 183172 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_1990
timestamp 1676037725
transform 1 0 184184 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2002
timestamp 1676037725
transform 1 0 185288 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2014
timestamp 1676037725
transform 1 0 186392 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_2017
timestamp 1676037725
transform 1 0 186668 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2030
timestamp 1676037725
transform 1 0 187864 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_2046
timestamp 1676037725
transform 1 0 189336 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_2054
timestamp 1676037725
transform 1 0 190072 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2061
timestamp 1676037725
transform 1 0 190716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_2069
timestamp 1676037725
transform 1 0 191452 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2073
timestamp 1676037725
transform 1 0 191820 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_2079
timestamp 1676037725
transform 1 0 192372 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2087
timestamp 1676037725
transform 1 0 193108 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2093
timestamp 1676037725
transform 1 0 193660 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_2101
timestamp 1676037725
transform 1 0 194396 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_2109
timestamp 1676037725
transform 1 0 195132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2116
timestamp 1676037725
transform 1 0 195776 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2120
timestamp 1676037725
transform 1 0 196144 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2126
timestamp 1676037725
transform 1 0 196696 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2129
timestamp 1676037725
transform 1 0 196972 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2136
timestamp 1676037725
transform 1 0 197616 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2140
timestamp 1676037725
transform 1 0 197984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2144
timestamp 1676037725
transform 1 0 198352 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2150
timestamp 1676037725
transform 1 0 198904 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_2158
timestamp 1676037725
transform 1 0 199640 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_2166
timestamp 1676037725
transform 1 0 200376 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2173
timestamp 1676037725
transform 1 0 201020 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_2181
timestamp 1676037725
transform 1 0 201756 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2185
timestamp 1676037725
transform 1 0 202124 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2192
timestamp 1676037725
transform 1 0 202768 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2201
timestamp 1676037725
transform 1 0 203596 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2213
timestamp 1676037725
transform 1 0 204700 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2225
timestamp 1676037725
transform 1 0 205804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_2237
timestamp 1676037725
transform 1 0 206908 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2241
timestamp 1676037725
transform 1 0 207276 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2253
timestamp 1676037725
transform 1 0 208380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2265
timestamp 1676037725
transform 1 0 209484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2277
timestamp 1676037725
transform 1 0 210588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2289
timestamp 1676037725
transform 1 0 211692 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2295
timestamp 1676037725
transform 1 0 212244 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2297
timestamp 1676037725
transform 1 0 212428 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2309
timestamp 1676037725
transform 1 0 213532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2321
timestamp 1676037725
transform 1 0 214636 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2333
timestamp 1676037725
transform 1 0 215740 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2345
timestamp 1676037725
transform 1 0 216844 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2351
timestamp 1676037725
transform 1 0 217396 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2353
timestamp 1676037725
transform 1 0 217580 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2365
timestamp 1676037725
transform 1 0 218684 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2377
timestamp 1676037725
transform 1 0 219788 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2389
timestamp 1676037725
transform 1 0 220892 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2401
timestamp 1676037725
transform 1 0 221996 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2407
timestamp 1676037725
transform 1 0 222548 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2409
timestamp 1676037725
transform 1 0 222732 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2423
timestamp 1676037725
transform 1 0 224020 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2430
timestamp 1676037725
transform 1 0 224664 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2438
timestamp 1676037725
transform 1 0 225400 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2446
timestamp 1676037725
transform 1 0 226136 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_2454
timestamp 1676037725
transform 1 0 226872 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2462
timestamp 1676037725
transform 1 0 227608 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2465
timestamp 1676037725
transform 1 0 227884 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2471
timestamp 1676037725
transform 1 0 228436 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2475
timestamp 1676037725
transform 1 0 228804 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2480
timestamp 1676037725
transform 1 0 229264 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2491
timestamp 1676037725
transform 1 0 230276 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2500
timestamp 1676037725
transform 1 0 231104 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2506
timestamp 1676037725
transform 1 0 231656 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_2511
timestamp 1676037725
transform 1 0 232116 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2519
timestamp 1676037725
transform 1 0 232852 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2521
timestamp 1676037725
transform 1 0 233036 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_2527
timestamp 1676037725
transform 1 0 233588 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2535
timestamp 1676037725
transform 1 0 234324 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2542
timestamp 1676037725
transform 1 0 234968 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2548
timestamp 1676037725
transform 1 0 235520 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2554
timestamp 1676037725
transform 1 0 236072 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2562
timestamp 1676037725
transform 1 0 236808 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2574
timestamp 1676037725
transform 1 0 237912 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2577
timestamp 1676037725
transform 1 0 238188 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2589
timestamp 1676037725
transform 1 0 239292 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2601
timestamp 1676037725
transform 1 0 240396 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2613
timestamp 1676037725
transform 1 0 241500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2625
timestamp 1676037725
transform 1 0 242604 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2631
timestamp 1676037725
transform 1 0 243156 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2633
timestamp 1676037725
transform 1 0 243340 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2645
timestamp 1676037725
transform 1 0 244444 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_2657
timestamp 1676037725
transform 1 0 245548 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2665
timestamp 1676037725
transform 1 0 246284 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2676
timestamp 1676037725
transform 1 0 247296 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_2689
timestamp 1676037725
transform 1 0 248492 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2697
timestamp 1676037725
transform 1 0 249228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2708
timestamp 1676037725
transform 1 0 250240 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2720
timestamp 1676037725
transform 1 0 251344 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2732
timestamp 1676037725
transform 1 0 252448 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_2745
timestamp 1676037725
transform 1 0 253644 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2753
timestamp 1676037725
transform 1 0 254380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_2764
timestamp 1676037725
transform 1 0 255392 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2776
timestamp 1676037725
transform 1 0 256496 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2788
timestamp 1676037725
transform 1 0 257600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2792
timestamp 1676037725
transform 1 0 257968 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_2797
timestamp 1676037725
transform 1 0 258428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2801
timestamp 1676037725
transform 1 0 258796 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2808
timestamp 1676037725
transform 1 0 259440 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_2819
timestamp 1676037725
transform 1 0 260452 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_2833
timestamp 1676037725
transform 1 0 261740 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_2839
timestamp 1676037725
transform 1 0 262292 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2846
timestamp 1676037725
transform 1 0 262936 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2850
timestamp 1676037725
transform 1 0 263304 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2854
timestamp 1676037725
transform 1 0 263672 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2857
timestamp 1676037725
transform 1 0 263948 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2865
timestamp 1676037725
transform 1 0 264684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2875
timestamp 1676037725
transform 1 0 265604 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2885
timestamp 1676037725
transform 1 0 266524 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_2889
timestamp 1676037725
transform 1 0 266892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2899
timestamp 1676037725
transform 1 0 267812 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2910
timestamp 1676037725
transform 1 0 268824 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2913
timestamp 1676037725
transform 1 0 269100 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_2920
timestamp 1676037725
transform 1 0 269744 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_2934
timestamp 1676037725
transform 1 0 271032 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_8
timestamp 1676037725
transform 1 0 1840 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_20
timestamp 1676037725
transform 1 0 2944 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_25
timestamp 1676037725
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 1676037725
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_105
timestamp 1676037725
transform 1 0 10764 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_113
timestamp 1676037725
transform 1 0 11500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_125
timestamp 1676037725
transform 1 0 12604 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_137
timestamp 1676037725
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1676037725
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_233
timestamp 1676037725
transform 1 0 22540 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_241
timestamp 1676037725
transform 1 0 23276 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_259
timestamp 1676037725
transform 1 0 24932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_266
timestamp 1676037725
transform 1 0 25576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_276
timestamp 1676037725
transform 1 0 26496 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_290
timestamp 1676037725
transform 1 0 27784 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_298
timestamp 1676037725
transform 1 0 28520 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_306
timestamp 1676037725
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_313
timestamp 1676037725
transform 1 0 29900 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_319
timestamp 1676037725
transform 1 0 30452 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_330
timestamp 1676037725
transform 1 0 31464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_339
timestamp 1676037725
transform 1 0 32292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_347
timestamp 1676037725
transform 1 0 33028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_355
timestamp 1676037725
transform 1 0 33764 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 1676037725
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_371
timestamp 1676037725
transform 1 0 35236 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_383
timestamp 1676037725
transform 1 0 36340 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_395
timestamp 1676037725
transform 1 0 37444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_407
timestamp 1676037725
transform 1 0 38548 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_419
timestamp 1676037725
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_427
timestamp 1676037725
transform 1 0 40388 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_439
timestamp 1676037725
transform 1 0 41492 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_451
timestamp 1676037725
transform 1 0 42596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_463
timestamp 1676037725
transform 1 0 43700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_475
timestamp 1676037725
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_483
timestamp 1676037725
transform 1 0 45540 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_495
timestamp 1676037725
transform 1 0 46644 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_507
timestamp 1676037725
transform 1 0 47748 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_519
timestamp 1676037725
transform 1 0 48852 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_531
timestamp 1676037725
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_533
timestamp 1676037725
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_545
timestamp 1676037725
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_557
timestamp 1676037725
transform 1 0 52348 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_563
timestamp 1676037725
transform 1 0 52900 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_568
timestamp 1676037725
transform 1 0 53360 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_577
timestamp 1676037725
transform 1 0 54188 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_586
timestamp 1676037725
transform 1 0 55016 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_589
timestamp 1676037725
transform 1 0 55292 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_596
timestamp 1676037725
transform 1 0 55936 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_605
timestamp 1676037725
transform 1 0 56764 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_614
timestamp 1676037725
transform 1 0 57592 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_623
timestamp 1676037725
transform 1 0 58420 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_632
timestamp 1676037725
transform 1 0 59248 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_641
timestamp 1676037725
transform 1 0 60076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_645
timestamp 1676037725
transform 1 0 60444 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_653
timestamp 1676037725
transform 1 0 61180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_662
timestamp 1676037725
transform 1 0 62008 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_671
timestamp 1676037725
transform 1 0 62836 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_680
timestamp 1676037725
transform 1 0 63664 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_689
timestamp 1676037725
transform 1 0 64492 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_698
timestamp 1676037725
transform 1 0 65320 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_701
timestamp 1676037725
transform 1 0 65596 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_710
timestamp 1676037725
transform 1 0 66424 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_724
timestamp 1676037725
transform 1 0 67712 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_736
timestamp 1676037725
transform 1 0 68816 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_754
timestamp 1676037725
transform 1 0 70472 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_757
timestamp 1676037725
transform 1 0 70748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_769
timestamp 1676037725
transform 1 0 71852 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_781
timestamp 1676037725
transform 1 0 72956 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_785
timestamp 1676037725
transform 1 0 73324 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_796
timestamp 1676037725
transform 1 0 74336 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_810
timestamp 1676037725
transform 1 0 75624 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_813
timestamp 1676037725
transform 1 0 75900 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_825
timestamp 1676037725
transform 1 0 77004 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_837
timestamp 1676037725
transform 1 0 78108 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_841
timestamp 1676037725
transform 1 0 78476 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_852
timestamp 1676037725
transform 1 0 79488 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_866
timestamp 1676037725
transform 1 0 80776 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_869
timestamp 1676037725
transform 1 0 81052 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_881
timestamp 1676037725
transform 1 0 82156 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_893
timestamp 1676037725
transform 1 0 83260 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_909
timestamp 1676037725
transform 1 0 84732 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_919
timestamp 1676037725
transform 1 0 85652 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_923
timestamp 1676037725
transform 1 0 86020 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_925
timestamp 1676037725
transform 1 0 86204 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_931
timestamp 1676037725
transform 1 0 86756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_943
timestamp 1676037725
transform 1 0 87860 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_951
timestamp 1676037725
transform 1 0 88596 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_960
timestamp 1676037725
transform 1 0 89424 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_969
timestamp 1676037725
transform 1 0 90252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_978
timestamp 1676037725
transform 1 0 91080 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_981
timestamp 1676037725
transform 1 0 91356 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_989
timestamp 1676037725
transform 1 0 92092 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_998
timestamp 1676037725
transform 1 0 92920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1007
timestamp 1676037725
transform 1 0 93748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1016
timestamp 1676037725
transform 1 0 94576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1025
timestamp 1676037725
transform 1 0 95404 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1034
timestamp 1676037725
transform 1 0 96232 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_1037
timestamp 1676037725
transform 1 0 96508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1045
timestamp 1676037725
transform 1 0 97244 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1054
timestamp 1676037725
transform 1 0 98072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1063
timestamp 1676037725
transform 1 0 98900 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1072
timestamp 1676037725
transform 1 0 99728 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_1086
timestamp 1676037725
transform 1 0 101016 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1093
timestamp 1676037725
transform 1 0 101660 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1105
timestamp 1676037725
transform 1 0 102764 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1117
timestamp 1676037725
transform 1 0 103868 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1129
timestamp 1676037725
transform 1 0 104972 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_1141
timestamp 1676037725
transform 1 0 106076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_1147
timestamp 1676037725
transform 1 0 106628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1149
timestamp 1676037725
transform 1 0 106812 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1154
timestamp 1676037725
transform 1 0 107272 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1166
timestamp 1676037725
transform 1 0 108376 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1178
timestamp 1676037725
transform 1 0 109480 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1190
timestamp 1676037725
transform 1 0 110584 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1202
timestamp 1676037725
transform 1 0 111688 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1205
timestamp 1676037725
transform 1 0 111964 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1210
timestamp 1676037725
transform 1 0 112424 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1222
timestamp 1676037725
transform 1 0 113528 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1234
timestamp 1676037725
transform 1 0 114632 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1246
timestamp 1676037725
transform 1 0 115736 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1258
timestamp 1676037725
transform 1 0 116840 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1261
timestamp 1676037725
transform 1 0 117116 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1266
timestamp 1676037725
transform 1 0 117576 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1278
timestamp 1676037725
transform 1 0 118680 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1290
timestamp 1676037725
transform 1 0 119784 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_1298
timestamp 1676037725
transform 1 0 120520 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1305
timestamp 1676037725
transform 1 0 121164 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1314
timestamp 1676037725
transform 1 0 121992 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_1317
timestamp 1676037725
transform 1 0 122268 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1325
timestamp 1676037725
transform 1 0 123004 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1334
timestamp 1676037725
transform 1 0 123832 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1343
timestamp 1676037725
transform 1 0 124660 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1352
timestamp 1676037725
transform 1 0 125488 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1361
timestamp 1676037725
transform 1 0 126316 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1370
timestamp 1676037725
transform 1 0 127144 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1373
timestamp 1676037725
transform 1 0 127420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1379
timestamp 1676037725
transform 1 0 127972 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1388
timestamp 1676037725
transform 1 0 128800 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_1392
timestamp 1676037725
transform 1 0 129168 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1403
timestamp 1676037725
transform 1 0 130180 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_1411
timestamp 1676037725
transform 1 0 130916 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1417
timestamp 1676037725
transform 1 0 131468 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1426
timestamp 1676037725
transform 1 0 132296 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1429
timestamp 1676037725
transform 1 0 132572 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_1433
timestamp 1676037725
transform 1 0 132940 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1439
timestamp 1676037725
transform 1 0 133492 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1448
timestamp 1676037725
transform 1 0 134320 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1456
timestamp 1676037725
transform 1 0 135056 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1463
timestamp 1676037725
transform 1 0 135700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1475
timestamp 1676037725
transform 1 0 136804 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_1483
timestamp 1676037725
transform 1 0 137540 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1485
timestamp 1676037725
transform 1 0 137724 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1497
timestamp 1676037725
transform 1 0 138828 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1508
timestamp 1676037725
transform 1 0 139840 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1520
timestamp 1676037725
transform 1 0 140944 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1532
timestamp 1676037725
transform 1 0 142048 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1541
timestamp 1676037725
transform 1 0 142876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1553
timestamp 1676037725
transform 1 0 143980 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1564
timestamp 1676037725
transform 1 0 144992 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1576
timestamp 1676037725
transform 1 0 146096 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1588
timestamp 1676037725
transform 1 0 147200 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1597
timestamp 1676037725
transform 1 0 148028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1609
timestamp 1676037725
transform 1 0 149132 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1620
timestamp 1676037725
transform 1 0 150144 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1632
timestamp 1676037725
transform 1 0 151248 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1644
timestamp 1676037725
transform 1 0 152352 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1653
timestamp 1676037725
transform 1 0 153180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_1665
timestamp 1676037725
transform 1 0 154284 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_1671
timestamp 1676037725
transform 1 0 154836 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1675
timestamp 1676037725
transform 1 0 155204 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1679
timestamp 1676037725
transform 1 0 155572 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1686
timestamp 1676037725
transform 1 0 156216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1695
timestamp 1676037725
transform 1 0 157044 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1704
timestamp 1676037725
transform 1 0 157872 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1709
timestamp 1676037725
transform 1 0 158332 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1720
timestamp 1676037725
transform 1 0 159344 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1733
timestamp 1676037725
transform 1 0 160540 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1744
timestamp 1676037725
transform 1 0 161552 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1748
timestamp 1676037725
transform 1 0 161920 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1759
timestamp 1676037725
transform 1 0 162932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_1763
timestamp 1676037725
transform 1 0 163300 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1765
timestamp 1676037725
transform 1 0 163484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1776
timestamp 1676037725
transform 1 0 164496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_1780
timestamp 1676037725
transform 1 0 164864 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1793
timestamp 1676037725
transform 1 0 166060 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1809
timestamp 1676037725
transform 1 0 167532 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1818
timestamp 1676037725
transform 1 0 168360 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1821
timestamp 1676037725
transform 1 0 168636 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1835
timestamp 1676037725
transform 1 0 169924 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1843
timestamp 1676037725
transform 1 0 170660 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1855
timestamp 1676037725
transform 1 0 171764 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1867
timestamp 1676037725
transform 1 0 172868 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_1875
timestamp 1676037725
transform 1 0 173604 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1877
timestamp 1676037725
transform 1 0 173788 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1883
timestamp 1676037725
transform 1 0 174340 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1895
timestamp 1676037725
transform 1 0 175444 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_1907
timestamp 1676037725
transform 1 0 176548 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1912
timestamp 1676037725
transform 1 0 177008 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_1920
timestamp 1676037725
transform 1 0 177744 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_1933
timestamp 1676037725
transform 1 0 178940 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_1939
timestamp 1676037725
transform 1 0 179492 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1950
timestamp 1676037725
transform 1 0 180504 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_1964
timestamp 1676037725
transform 1 0 181792 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_1978
timestamp 1676037725
transform 1 0 183080 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1986
timestamp 1676037725
transform 1 0 183816 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_1989
timestamp 1676037725
transform 1 0 184092 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2001
timestamp 1676037725
transform 1 0 185196 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2015
timestamp 1676037725
transform 1 0 186484 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2029
timestamp 1676037725
transform 1 0 187772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_2041
timestamp 1676037725
transform 1 0 188876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2045
timestamp 1676037725
transform 1 0 189244 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2057
timestamp 1676037725
transform 1 0 190348 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2064
timestamp 1676037725
transform 1 0 190992 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2068
timestamp 1676037725
transform 1 0 191360 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2075
timestamp 1676037725
transform 1 0 192004 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2084
timestamp 1676037725
transform 1 0 192832 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2093
timestamp 1676037725
transform 1 0 193660 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_2099
timestamp 1676037725
transform 1 0 194212 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2101
timestamp 1676037725
transform 1 0 194396 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2108
timestamp 1676037725
transform 1 0 195040 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2117
timestamp 1676037725
transform 1 0 195868 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2126
timestamp 1676037725
transform 1 0 196696 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2142
timestamp 1676037725
transform 1 0 198168 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2151
timestamp 1676037725
transform 1 0 198996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_2155
timestamp 1676037725
transform 1 0 199364 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2157
timestamp 1676037725
transform 1 0 199548 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2164
timestamp 1676037725
transform 1 0 200192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2173
timestamp 1676037725
transform 1 0 201020 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2182
timestamp 1676037725
transform 1 0 201848 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2189
timestamp 1676037725
transform 1 0 202492 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2193
timestamp 1676037725
transform 1 0 202860 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2200
timestamp 1676037725
transform 1 0 203504 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2208
timestamp 1676037725
transform 1 0 204240 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2213
timestamp 1676037725
transform 1 0 204700 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2225
timestamp 1676037725
transform 1 0 205804 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2237
timestamp 1676037725
transform 1 0 206908 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2249
timestamp 1676037725
transform 1 0 208012 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2261
timestamp 1676037725
transform 1 0 209116 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_2267
timestamp 1676037725
transform 1 0 209668 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2269
timestamp 1676037725
transform 1 0 209852 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2281
timestamp 1676037725
transform 1 0 210956 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2290
timestamp 1676037725
transform 1 0 211784 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2302
timestamp 1676037725
transform 1 0 212888 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_2314
timestamp 1676037725
transform 1 0 213992 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2322
timestamp 1676037725
transform 1 0 214728 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2325
timestamp 1676037725
transform 1 0 215004 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2337
timestamp 1676037725
transform 1 0 216108 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2346
timestamp 1676037725
transform 1 0 216936 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2358
timestamp 1676037725
transform 1 0 218040 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_2370
timestamp 1676037725
transform 1 0 219144 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2378
timestamp 1676037725
transform 1 0 219880 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2381
timestamp 1676037725
transform 1 0 220156 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2393
timestamp 1676037725
transform 1 0 221260 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2402
timestamp 1676037725
transform 1 0 222088 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2418
timestamp 1676037725
transform 1 0 223560 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_2427
timestamp 1676037725
transform 1 0 224388 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_2435
timestamp 1676037725
transform 1 0 225124 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2437
timestamp 1676037725
transform 1 0 225308 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2444
timestamp 1676037725
transform 1 0 225952 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2453
timestamp 1676037725
transform 1 0 226780 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2462
timestamp 1676037725
transform 1 0 227608 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2471
timestamp 1676037725
transform 1 0 228436 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2480
timestamp 1676037725
transform 1 0 229264 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_2489
timestamp 1676037725
transform 1 0 230092 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_2493
timestamp 1676037725
transform 1 0 230460 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2506
timestamp 1676037725
transform 1 0 231656 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2515
timestamp 1676037725
transform 1 0 232484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2524
timestamp 1676037725
transform 1 0 233312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2533
timestamp 1676037725
transform 1 0 234140 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2542
timestamp 1676037725
transform 1 0 234968 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2549
timestamp 1676037725
transform 1 0 235612 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2556
timestamp 1676037725
transform 1 0 236256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2564
timestamp 1676037725
transform 1 0 236992 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2572
timestamp 1676037725
transform 1 0 237728 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2584
timestamp 1676037725
transform 1 0 238832 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_2596
timestamp 1676037725
transform 1 0 239936 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2605
timestamp 1676037725
transform 1 0 240764 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_2617
timestamp 1676037725
transform 1 0 241868 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2628
timestamp 1676037725
transform 1 0 242880 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2644
timestamp 1676037725
transform 1 0 244352 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2658
timestamp 1676037725
transform 1 0 245640 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2661
timestamp 1676037725
transform 1 0 245916 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2673
timestamp 1676037725
transform 1 0 247020 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2687
timestamp 1676037725
transform 1 0 248308 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2701
timestamp 1676037725
transform 1 0 249596 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_2713
timestamp 1676037725
transform 1 0 250700 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2717
timestamp 1676037725
transform 1 0 251068 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2729
timestamp 1676037725
transform 1 0 252172 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2743
timestamp 1676037725
transform 1 0 253460 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_2757
timestamp 1676037725
transform 1 0 254748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_2769
timestamp 1676037725
transform 1 0 255852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2773
timestamp 1676037725
transform 1 0 256220 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2785
timestamp 1676037725
transform 1 0 257324 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2799
timestamp 1676037725
transform 1 0 258612 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2809
timestamp 1676037725
transform 1 0 259532 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_2813
timestamp 1676037725
transform 1 0 259900 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_2820
timestamp 1676037725
transform 1 0 260544 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2829
timestamp 1676037725
transform 1 0 261372 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2837
timestamp 1676037725
transform 1 0 262108 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2847
timestamp 1676037725
transform 1 0 263028 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_2853
timestamp 1676037725
transform 1 0 263580 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2864
timestamp 1676037725
transform 1 0 264592 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2868
timestamp 1676037725
transform 1 0 264960 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_2876
timestamp 1676037725
transform 1 0 265696 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2885
timestamp 1676037725
transform 1 0 266524 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_2893
timestamp 1676037725
transform 1 0 267260 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2906
timestamp 1676037725
transform 1 0 268456 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_2920
timestamp 1676037725
transform 1 0 269744 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_2934
timestamp 1676037725
transform 1 0 271032 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_9
timestamp 1676037725
transform 1 0 1932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_17
timestamp 1676037725
transform 1 0 2668 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_21
timestamp 1676037725
transform 1 0 3036 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_26
timestamp 1676037725
transform 1 0 3496 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_29
timestamp 1676037725
transform 1 0 3772 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_33
timestamp 1676037725
transform 1 0 4140 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_38
timestamp 1676037725
transform 1 0 4600 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_46
timestamp 1676037725
transform 1 0 5336 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_65
timestamp 1676037725
transform 1 0 7084 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_73
timestamp 1676037725
transform 1 0 7820 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_77
timestamp 1676037725
transform 1 0 8188 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_82
timestamp 1676037725
transform 1 0 8648 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_85
timestamp 1676037725
transform 1 0 8924 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_103
timestamp 1676037725
transform 1 0 10580 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_121
timestamp 1676037725
transform 1 0 12236 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_129
timestamp 1676037725
transform 1 0 12972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_133
timestamp 1676037725
transform 1 0 13340 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_138
timestamp 1676037725
transform 1 0 13800 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_141
timestamp 1676037725
transform 1 0 14076 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_145
timestamp 1676037725
transform 1 0 14444 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_150
timestamp 1676037725
transform 1 0 14904 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_158
timestamp 1676037725
transform 1 0 15640 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_177
timestamp 1676037725
transform 1 0 17388 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_185
timestamp 1676037725
transform 1 0 18124 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_193
timestamp 1676037725
transform 1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_197
timestamp 1676037725
transform 1 0 19228 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_209
timestamp 1676037725
transform 1 0 20332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_221
timestamp 1676037725
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_237
timestamp 1676037725
transform 1 0 22908 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_250
timestamp 1676037725
transform 1 0 24104 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_253
timestamp 1676037725
transform 1 0 24380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_259
timestamp 1676037725
transform 1 0 24932 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_266
timestamp 1676037725
transform 1 0 25576 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_272
timestamp 1676037725
transform 1 0 26128 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_278
timestamp 1676037725
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_289
timestamp 1676037725
transform 1 0 27692 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_295
timestamp 1676037725
transform 1 0 28244 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_303
timestamp 1676037725
transform 1 0 28980 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_307
timestamp 1676037725
transform 1 0 29348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_309
timestamp 1676037725
transform 1 0 29532 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_315
timestamp 1676037725
transform 1 0 30084 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_327
timestamp 1676037725
transform 1 0 31188 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 1676037725
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_344
timestamp 1676037725
transform 1 0 32752 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_356
timestamp 1676037725
transform 1 0 33856 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_365
timestamp 1676037725
transform 1 0 34684 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_376
timestamp 1676037725
transform 1 0 35696 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_383
timestamp 1676037725
transform 1 0 36340 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_390
timestamp 1676037725
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_399
timestamp 1676037725
transform 1 0 37812 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_403
timestamp 1676037725
transform 1 0 38180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_407
timestamp 1676037725
transform 1 0 38548 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_411
timestamp 1676037725
transform 1 0 38916 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_418
timestamp 1676037725
transform 1 0 39560 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_421
timestamp 1676037725
transform 1 0 39836 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_432
timestamp 1676037725
transform 1 0 40848 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_439
timestamp 1676037725
transform 1 0 41492 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_446
timestamp 1676037725
transform 1 0 42136 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_455
timestamp 1676037725
transform 1 0 42964 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_459
timestamp 1676037725
transform 1 0 43332 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_463
timestamp 1676037725
transform 1 0 43700 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_467
timestamp 1676037725
transform 1 0 44068 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_474
timestamp 1676037725
transform 1 0 44712 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_477
timestamp 1676037725
transform 1 0 44988 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_488
timestamp 1676037725
transform 1 0 46000 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_495
timestamp 1676037725
transform 1 0 46644 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_502
timestamp 1676037725
transform 1 0 47288 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_511
timestamp 1676037725
transform 1 0 48116 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_515
timestamp 1676037725
transform 1 0 48484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_519
timestamp 1676037725
transform 1 0 48852 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_523
timestamp 1676037725
transform 1 0 49220 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_530
timestamp 1676037725
transform 1 0 49864 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_533
timestamp 1676037725
transform 1 0 50140 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_539
timestamp 1676037725
transform 1 0 50692 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_543
timestamp 1676037725
transform 1 0 51060 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_547
timestamp 1676037725
transform 1 0 51428 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_551
timestamp 1676037725
transform 1 0 51796 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_555
timestamp 1676037725
transform 1 0 52164 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_559
timestamp 1676037725
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_561
timestamp 1676037725
transform 1 0 52716 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_565
timestamp 1676037725
transform 1 0 53084 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_569
timestamp 1676037725
transform 1 0 53452 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_576
timestamp 1676037725
transform 1 0 54096 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_584
timestamp 1676037725
transform 1 0 54832 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_589
timestamp 1676037725
transform 1 0 55292 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_601
timestamp 1676037725
transform 1 0 56396 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_613
timestamp 1676037725
transform 1 0 57500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_617
timestamp 1676037725
transform 1 0 57868 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_623
timestamp 1676037725
transform 1 0 58420 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_629
timestamp 1676037725
transform 1 0 58972 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_634
timestamp 1676037725
transform 1 0 59432 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_642
timestamp 1676037725
transform 1 0 60168 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_645
timestamp 1676037725
transform 1 0 60444 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_651
timestamp 1676037725
transform 1 0 60996 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_663
timestamp 1676037725
transform 1 0 62100 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_671
timestamp 1676037725
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_673
timestamp 1676037725
transform 1 0 63020 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_679
timestamp 1676037725
transform 1 0 63572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_691
timestamp 1676037725
transform 1 0 64676 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_699
timestamp 1676037725
transform 1 0 65412 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_701
timestamp 1676037725
transform 1 0 65596 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_709
timestamp 1676037725
transform 1 0 66332 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_717
timestamp 1676037725
transform 1 0 67068 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_725
timestamp 1676037725
transform 1 0 67804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_729
timestamp 1676037725
transform 1 0 68172 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_740
timestamp 1676037725
transform 1 0 69184 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_754
timestamp 1676037725
transform 1 0 70472 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_757
timestamp 1676037725
transform 1 0 70748 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_769
timestamp 1676037725
transform 1 0 71852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_782
timestamp 1676037725
transform 1 0 73048 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_785
timestamp 1676037725
transform 1 0 73324 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_797
timestamp 1676037725
transform 1 0 74428 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_810
timestamp 1676037725
transform 1 0 75624 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_813
timestamp 1676037725
transform 1 0 75900 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_825
timestamp 1676037725
transform 1 0 77004 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_838
timestamp 1676037725
transform 1 0 78200 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_841
timestamp 1676037725
transform 1 0 78476 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_853
timestamp 1676037725
transform 1 0 79580 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_866
timestamp 1676037725
transform 1 0 80776 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_869
timestamp 1676037725
transform 1 0 81052 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_881
timestamp 1676037725
transform 1 0 82156 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_894
timestamp 1676037725
transform 1 0 83352 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_897
timestamp 1676037725
transform 1 0 83628 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_905
timestamp 1676037725
transform 1 0 84364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_917
timestamp 1676037725
transform 1 0 85468 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_923
timestamp 1676037725
transform 1 0 86020 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_925
timestamp 1676037725
transform 1 0 86204 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_941
timestamp 1676037725
transform 1 0 87676 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_949
timestamp 1676037725
transform 1 0 88412 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_953
timestamp 1676037725
transform 1 0 88780 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_961
timestamp 1676037725
transform 1 0 89516 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_965
timestamp 1676037725
transform 1 0 89884 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_972
timestamp 1676037725
transform 1 0 90528 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_981
timestamp 1676037725
transform 1 0 91356 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_993
timestamp 1676037725
transform 1 0 92460 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1001
timestamp 1676037725
transform 1 0 93196 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1006
timestamp 1676037725
transform 1 0 93656 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1009
timestamp 1676037725
transform 1 0 93932 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1021
timestamp 1676037725
transform 1 0 95036 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_1033
timestamp 1676037725
transform 1 0 96140 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1037
timestamp 1676037725
transform 1 0 96508 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1043
timestamp 1676037725
transform 1 0 97060 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1051
timestamp 1676037725
transform 1 0 97796 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_1057
timestamp 1676037725
transform 1 0 98348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1063
timestamp 1676037725
transform 1 0 98900 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1065
timestamp 1676037725
transform 1 0 99084 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1072
timestamp 1676037725
transform 1 0 99728 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1084
timestamp 1676037725
transform 1 0 100832 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_1093
timestamp 1676037725
transform 1 0 101660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_1105
timestamp 1676037725
transform 1 0 102764 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1111
timestamp 1676037725
transform 1 0 103316 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1118
timestamp 1676037725
transform 1 0 103960 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1121
timestamp 1676037725
transform 1 0 104236 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1125
timestamp 1676037725
transform 1 0 104604 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1129
timestamp 1676037725
transform 1 0 104972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1133
timestamp 1676037725
transform 1 0 105340 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1137
timestamp 1676037725
transform 1 0 105708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1141
timestamp 1676037725
transform 1 0 106076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_1145
timestamp 1676037725
transform 1 0 106444 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1149
timestamp 1676037725
transform 1 0 106812 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1160
timestamp 1676037725
transform 1 0 107824 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1167
timestamp 1676037725
transform 1 0 108468 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1174
timestamp 1676037725
transform 1 0 109112 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1177
timestamp 1676037725
transform 1 0 109388 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1181
timestamp 1676037725
transform 1 0 109756 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1185
timestamp 1676037725
transform 1 0 110124 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1189
timestamp 1676037725
transform 1 0 110492 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1193
timestamp 1676037725
transform 1 0 110860 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1197
timestamp 1676037725
transform 1 0 111228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_1201
timestamp 1676037725
transform 1 0 111596 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1205
timestamp 1676037725
transform 1 0 111964 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1216
timestamp 1676037725
transform 1 0 112976 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1223
timestamp 1676037725
transform 1 0 113620 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1230
timestamp 1676037725
transform 1 0 114264 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1233
timestamp 1676037725
transform 1 0 114540 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1237
timestamp 1676037725
transform 1 0 114908 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1241
timestamp 1676037725
transform 1 0 115276 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1245
timestamp 1676037725
transform 1 0 115644 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1249
timestamp 1676037725
transform 1 0 116012 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1253
timestamp 1676037725
transform 1 0 116380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_1257
timestamp 1676037725
transform 1 0 116748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1261
timestamp 1676037725
transform 1 0 117116 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1272
timestamp 1676037725
transform 1 0 118128 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1279
timestamp 1676037725
transform 1 0 118772 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1286
timestamp 1676037725
transform 1 0 119416 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1289
timestamp 1676037725
transform 1 0 119692 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1293
timestamp 1676037725
transform 1 0 120060 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1297
timestamp 1676037725
transform 1 0 120428 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1301
timestamp 1676037725
transform 1 0 120796 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1305
timestamp 1676037725
transform 1 0 121164 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1309
timestamp 1676037725
transform 1 0 121532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1314
timestamp 1676037725
transform 1 0 121992 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1317
timestamp 1676037725
transform 1 0 122268 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_1323
timestamp 1676037725
transform 1 0 122820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1335
timestamp 1676037725
transform 1 0 123924 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1343
timestamp 1676037725
transform 1 0 124660 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1345
timestamp 1676037725
transform 1 0 124844 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_1351
timestamp 1676037725
transform 1 0 125396 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1363
timestamp 1676037725
transform 1 0 126500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1371
timestamp 1676037725
transform 1 0 127236 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_1373
timestamp 1676037725
transform 1 0 127420 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_1380
timestamp 1676037725
transform 1 0 128064 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1390
timestamp 1676037725
transform 1 0 128984 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1398
timestamp 1676037725
transform 1 0 129720 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1401
timestamp 1676037725
transform 1 0 129996 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_1408
timestamp 1676037725
transform 1 0 130640 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1414
timestamp 1676037725
transform 1 0 131192 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1419
timestamp 1676037725
transform 1 0 131652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1427
timestamp 1676037725
transform 1 0 132388 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1429
timestamp 1676037725
transform 1 0 132572 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1441
timestamp 1676037725
transform 1 0 133676 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_1449
timestamp 1676037725
transform 1 0 134412 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1455
timestamp 1676037725
transform 1 0 134964 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_1457
timestamp 1676037725
transform 1 0 135148 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_1469
timestamp 1676037725
transform 1 0 136252 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_1481
timestamp 1676037725
transform 1 0 137356 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1485
timestamp 1676037725
transform 1 0 137724 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1490
timestamp 1676037725
transform 1 0 138184 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1497
timestamp 1676037725
transform 1 0 138828 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1504
timestamp 1676037725
transform 1 0 139472 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1513
timestamp 1676037725
transform 1 0 140300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1518
timestamp 1676037725
transform 1 0 140760 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1525
timestamp 1676037725
transform 1 0 141404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1532
timestamp 1676037725
transform 1 0 142048 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1541
timestamp 1676037725
transform 1 0 142876 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1546
timestamp 1676037725
transform 1 0 143336 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1553
timestamp 1676037725
transform 1 0 143980 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1560
timestamp 1676037725
transform 1 0 144624 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1569
timestamp 1676037725
transform 1 0 145452 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1574
timestamp 1676037725
transform 1 0 145912 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1581
timestamp 1676037725
transform 1 0 146556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1588
timestamp 1676037725
transform 1 0 147200 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1597
timestamp 1676037725
transform 1 0 148028 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1602
timestamp 1676037725
transform 1 0 148488 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1609
timestamp 1676037725
transform 1 0 149132 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1616
timestamp 1676037725
transform 1 0 149776 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1625
timestamp 1676037725
transform 1 0 150604 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1630
timestamp 1676037725
transform 1 0 151064 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1637
timestamp 1676037725
transform 1 0 151708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1644
timestamp 1676037725
transform 1 0 152352 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1653
timestamp 1676037725
transform 1 0 153180 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1658
timestamp 1676037725
transform 1 0 153640 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1665
timestamp 1676037725
transform 1 0 154284 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1672
timestamp 1676037725
transform 1 0 154928 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1681
timestamp 1676037725
transform 1 0 155756 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1687
timestamp 1676037725
transform 1 0 156308 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1695
timestamp 1676037725
transform 1 0 157044 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1703
timestamp 1676037725
transform 1 0 157780 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1707
timestamp 1676037725
transform 1 0 158148 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1709
timestamp 1676037725
transform 1 0 158332 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1715
timestamp 1676037725
transform 1 0 158884 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1723
timestamp 1676037725
transform 1 0 159620 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1731
timestamp 1676037725
transform 1 0 160356 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1735
timestamp 1676037725
transform 1 0 160724 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1737
timestamp 1676037725
transform 1 0 160908 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_1744
timestamp 1676037725
transform 1 0 161552 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1749
timestamp 1676037725
transform 1 0 162012 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1760
timestamp 1676037725
transform 1 0 163024 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1765
timestamp 1676037725
transform 1 0 163484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1771
timestamp 1676037725
transform 1 0 164036 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1782
timestamp 1676037725
transform 1 0 165048 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1790
timestamp 1676037725
transform 1 0 165784 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1793
timestamp 1676037725
transform 1 0 166060 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1800
timestamp 1676037725
transform 1 0 166704 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1809
timestamp 1676037725
transform 1 0 167532 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1818
timestamp 1676037725
transform 1 0 168360 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1821
timestamp 1676037725
transform 1 0 168636 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1825
timestamp 1676037725
transform 1 0 169004 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_1836
timestamp 1676037725
transform 1 0 170016 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_1849
timestamp 1676037725
transform 1 0 171212 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1855
timestamp 1676037725
transform 1 0 171764 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1859
timestamp 1676037725
transform 1 0 172132 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1864
timestamp 1676037725
transform 1 0 172592 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1872
timestamp 1676037725
transform 1 0 173328 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_1877
timestamp 1676037725
transform 1 0 173788 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1883
timestamp 1676037725
transform 1 0 174340 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_1894
timestamp 1676037725
transform 1 0 175352 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1902
timestamp 1676037725
transform 1 0 176088 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1905
timestamp 1676037725
transform 1 0 176364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_1911
timestamp 1676037725
transform 1 0 176916 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_1919
timestamp 1676037725
transform 1 0 177652 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1930
timestamp 1676037725
transform 1 0 178664 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1933
timestamp 1676037725
transform 1 0 178940 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_1945
timestamp 1676037725
transform 1 0 180044 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_1957
timestamp 1676037725
transform 1 0 181148 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1961
timestamp 1676037725
transform 1 0 181516 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_1973
timestamp 1676037725
transform 1 0 182620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_1985
timestamp 1676037725
transform 1 0 183724 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_1989
timestamp 1676037725
transform 1 0 184092 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2001
timestamp 1676037725
transform 1 0 185196 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_2013
timestamp 1676037725
transform 1 0 186300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2017
timestamp 1676037725
transform 1 0 186668 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2029
timestamp 1676037725
transform 1 0 187772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_2041
timestamp 1676037725
transform 1 0 188876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2045
timestamp 1676037725
transform 1 0 189244 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2057
timestamp 1676037725
transform 1 0 190348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_2065
timestamp 1676037725
transform 1 0 191084 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2071
timestamp 1676037725
transform 1 0 191636 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_2073
timestamp 1676037725
transform 1 0 191820 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2083
timestamp 1676037725
transform 1 0 192740 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2087
timestamp 1676037725
transform 1 0 193108 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2092
timestamp 1676037725
transform 1 0 193568 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_2101
timestamp 1676037725
transform 1 0 194396 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2108
timestamp 1676037725
transform 1 0 195040 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2124
timestamp 1676037725
transform 1 0 196512 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2129
timestamp 1676037725
transform 1 0 196972 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2135
timestamp 1676037725
transform 1 0 197524 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2143
timestamp 1676037725
transform 1 0 198260 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2151
timestamp 1676037725
transform 1 0 198996 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2155
timestamp 1676037725
transform 1 0 199364 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_2157
timestamp 1676037725
transform 1 0 199548 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2164
timestamp 1676037725
transform 1 0 200192 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2176
timestamp 1676037725
transform 1 0 201296 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2185
timestamp 1676037725
transform 1 0 202124 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2191
timestamp 1676037725
transform 1 0 202676 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2199
timestamp 1676037725
transform 1 0 203412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2211
timestamp 1676037725
transform 1 0 204516 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2213
timestamp 1676037725
transform 1 0 204700 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2221
timestamp 1676037725
transform 1 0 205436 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2226
timestamp 1676037725
transform 1 0 205896 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2230
timestamp 1676037725
transform 1 0 206264 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_2234
timestamp 1676037725
transform 1 0 206632 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2241
timestamp 1676037725
transform 1 0 207276 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2246
timestamp 1676037725
transform 1 0 207736 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2253
timestamp 1676037725
transform 1 0 208380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2260
timestamp 1676037725
transform 1 0 209024 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2269
timestamp 1676037725
transform 1 0 209852 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2274
timestamp 1676037725
transform 1 0 210312 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2281
timestamp 1676037725
transform 1 0 210956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2288
timestamp 1676037725
transform 1 0 211600 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2297
timestamp 1676037725
transform 1 0 212428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2302
timestamp 1676037725
transform 1 0 212888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2309
timestamp 1676037725
transform 1 0 213532 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2316
timestamp 1676037725
transform 1 0 214176 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2325
timestamp 1676037725
transform 1 0 215004 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2330
timestamp 1676037725
transform 1 0 215464 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2337
timestamp 1676037725
transform 1 0 216108 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2344
timestamp 1676037725
transform 1 0 216752 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2353
timestamp 1676037725
transform 1 0 217580 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2358
timestamp 1676037725
transform 1 0 218040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2365
timestamp 1676037725
transform 1 0 218684 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2372
timestamp 1676037725
transform 1 0 219328 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2381
timestamp 1676037725
transform 1 0 220156 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2386
timestamp 1676037725
transform 1 0 220616 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2393
timestamp 1676037725
transform 1 0 221260 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2400
timestamp 1676037725
transform 1 0 221904 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2409
timestamp 1676037725
transform 1 0 222732 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2414
timestamp 1676037725
transform 1 0 223192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2421
timestamp 1676037725
transform 1 0 223836 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2434
timestamp 1676037725
transform 1 0 225032 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2437
timestamp 1676037725
transform 1 0 225308 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2443
timestamp 1676037725
transform 1 0 225860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2455
timestamp 1676037725
transform 1 0 226964 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2463
timestamp 1676037725
transform 1 0 227700 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_2465
timestamp 1676037725
transform 1 0 227884 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2472
timestamp 1676037725
transform 1 0 228528 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2488
timestamp 1676037725
transform 1 0 230000 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2493
timestamp 1676037725
transform 1 0 230460 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2499
timestamp 1676037725
transform 1 0 231012 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2507
timestamp 1676037725
transform 1 0 231748 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2519
timestamp 1676037725
transform 1 0 232852 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_2521
timestamp 1676037725
transform 1 0 233036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2528
timestamp 1676037725
transform 1 0 233680 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2532
timestamp 1676037725
transform 1 0 234048 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2537
timestamp 1676037725
transform 1 0 234508 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_2545
timestamp 1676037725
transform 1 0 235244 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2549
timestamp 1676037725
transform 1 0 235612 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2556
timestamp 1676037725
transform 1 0 236256 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2560
timestamp 1676037725
transform 1 0 236624 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2572
timestamp 1676037725
transform 1 0 237728 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2577
timestamp 1676037725
transform 1 0 238188 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2589
timestamp 1676037725
transform 1 0 239292 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2594
timestamp 1676037725
transform 1 0 239752 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2602
timestamp 1676037725
transform 1 0 240488 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2605
timestamp 1676037725
transform 1 0 240764 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2609
timestamp 1676037725
transform 1 0 241132 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2620
timestamp 1676037725
transform 1 0 242144 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2633
timestamp 1676037725
transform 1 0 243340 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2645
timestamp 1676037725
transform 1 0 244444 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_2657
timestamp 1676037725
transform 1 0 245548 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2661
timestamp 1676037725
transform 1 0 245916 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2673
timestamp 1676037725
transform 1 0 247020 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_2685
timestamp 1676037725
transform 1 0 248124 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2689
timestamp 1676037725
transform 1 0 248492 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2701
timestamp 1676037725
transform 1 0 249596 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_2713
timestamp 1676037725
transform 1 0 250700 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2717
timestamp 1676037725
transform 1 0 251068 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_2729
timestamp 1676037725
transform 1 0 252172 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_2741
timestamp 1676037725
transform 1 0 253276 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2745
timestamp 1676037725
transform 1 0 253644 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_2757
timestamp 1676037725
transform 1 0 254748 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2765
timestamp 1676037725
transform 1 0 255484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2770
timestamp 1676037725
transform 1 0 255944 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2773
timestamp 1676037725
transform 1 0 256220 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2785
timestamp 1676037725
transform 1 0 257324 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2789
timestamp 1676037725
transform 1 0 257692 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2795
timestamp 1676037725
transform 1 0 258244 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2799
timestamp 1676037725
transform 1 0 258612 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2801
timestamp 1676037725
transform 1 0 258796 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2808
timestamp 1676037725
transform 1 0 259440 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2816
timestamp 1676037725
transform 1 0 260176 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2820
timestamp 1676037725
transform 1 0 260544 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2826
timestamp 1676037725
transform 1 0 261096 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2829
timestamp 1676037725
transform 1 0 261372 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2836
timestamp 1676037725
transform 1 0 262016 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2842
timestamp 1676037725
transform 1 0 262568 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2846
timestamp 1676037725
transform 1 0 262936 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2854
timestamp 1676037725
transform 1 0 263672 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2857
timestamp 1676037725
transform 1 0 263948 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2864
timestamp 1676037725
transform 1 0 264592 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2873
timestamp 1676037725
transform 1 0 265420 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2882
timestamp 1676037725
transform 1 0 266248 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2885
timestamp 1676037725
transform 1 0 266524 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_2889
timestamp 1676037725
transform 1 0 266892 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2896
timestamp 1676037725
transform 1 0 267536 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2900
timestamp 1676037725
transform 1 0 267904 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2908
timestamp 1676037725
transform 1 0 268640 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2913
timestamp 1676037725
transform 1 0 269100 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_2920
timestamp 1676037725
transform 1 0 269744 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_2934
timestamp 1676037725
transform 1 0 271032 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 265328 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 264408 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 263028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1676037725
transform 1 0 255668 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 259624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 265696 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1676037725
transform 1 0 262016 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1676037725
transform 1 0 262660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 263396 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 268548 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1676037725
transform 1 0 270756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 268456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1676037725
transform 1 0 267812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1676037725
transform 1 0 266984 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1676037725
transform 1 0 267904 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1676037725
transform 1 0 268824 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1676037725
transform 1 0 267168 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1676037725
transform 1 0 266340 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform 1 0 265144 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1676037725
transform 1 0 268364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1676037725
transform 1 0 267260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1676037725
transform 1 0 267720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1676037725
transform 1 0 266616 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1676037725
transform 1 0 265972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1676037725
transform 1 0 265052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1676037725
transform 1 0 267076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1676037725
transform 1 0 270112 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1676037725
transform 1 0 270112 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1676037725
transform 1 0 270112 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 1676037725
transform 1 0 270112 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1676037725
transform 1 0 259624 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1676037725
transform 1 0 270112 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 260268 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1676037725
transform 1 0 260912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1676037725
transform 1 0 18492 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1676037725
transform 1 0 82432 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input37
timestamp 1676037725
transform 1 0 82064 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1676037725
transform 1 0 82064 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1676037725
transform 1 0 81144 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1676037725
transform 1 0 79856 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1676037725
transform 1 0 79856 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1676037725
transform 1 0 79396 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp 1676037725
transform 1 0 77280 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1676037725
transform 1 0 77924 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1676037725
transform 1 0 77188 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1676037725
transform 1 0 10856 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1676037725
transform 1 0 76452 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp 1676037725
transform 1 0 75716 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1676037725
transform 1 0 74704 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1676037725
transform 1 0 74244 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1676037725
transform 1 0 73508 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1676037725
transform 1 0 72128 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1676037725
transform 1 0 72036 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1676037725
transform 1 0 71300 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input55
timestamp 1676037725
transform 1 0 70564 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1676037725
transform 1 0 69552 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1676037725
transform 1 0 10120 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1676037725
transform 1 0 86756 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1676037725
transform 1 0 86388 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1676037725
transform 1 0 85284 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1676037725
transform 1 0 84548 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1676037725
transform 1 0 83812 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 1676037725
transform 1 0 82432 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1676037725
transform 1 0 82340 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1676037725
transform 1 0 81604 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1676037725
transform 1 0 79856 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1676037725
transform 1 0 79856 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1676037725
transform 1 0 9384 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input69
timestamp 1676037725
transform 1 0 79396 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input70
timestamp 1676037725
transform 1 0 78568 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input71
timestamp 1676037725
transform 1 0 77280 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input72
timestamp 1676037725
transform 1 0 77188 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 1676037725
transform 1 0 76452 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1676037725
transform 1 0 74704 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1676037725
transform 1 0 74704 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1676037725
transform 1 0 74244 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1676037725
transform 1 0 73416 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input78
timestamp 1676037725
transform 1 0 72128 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1676037725
transform 1 0 8924 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input80
timestamp 1676037725
transform 1 0 72036 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input81
timestamp 1676037725
transform 1 0 71300 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input82
timestamp 1676037725
transform 1 0 69552 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input83
timestamp 1676037725
transform 1 0 69552 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1676037725
transform 1 0 120888 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1676037725
transform 1 0 120152 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1676037725
transform 1 0 119140 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1676037725
transform 1 0 118496 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1676037725
transform 1 0 117852 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1676037725
transform 1 0 117208 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1676037725
transform 1 0 8188 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1676037725
transform 1 0 116472 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1676037725
transform 1 0 115736 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1676037725
transform 1 0 115000 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1676037725
transform 1 0 113988 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1676037725
transform 1 0 113344 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1676037725
transform 1 0 112700 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 1676037725
transform 1 0 112056 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1676037725
transform 1 0 111320 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input99
timestamp 1676037725
transform 1 0 110584 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1676037725
transform 1 0 109848 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1676037725
transform 1 0 7452 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input102
timestamp 1676037725
transform 1 0 108836 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input103
timestamp 1676037725
transform 1 0 108192 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 1676037725
transform 1 0 107548 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 1676037725
transform 1 0 106904 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input106
timestamp 1676037725
transform 1 0 106168 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 1676037725
transform 1 0 105432 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input108
timestamp 1676037725
transform 1 0 104696 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1676037725
transform 1 0 103684 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 1676037725
transform 1 0 120888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input111
timestamp 1676037725
transform 1 0 120152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input112
timestamp 1676037725
transform 1 0 6716 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input113
timestamp 1676037725
transform 1 0 119140 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input114
timestamp 1676037725
transform 1 0 118496 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input115
timestamp 1676037725
transform 1 0 117852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input116
timestamp 1676037725
transform 1 0 117300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input117
timestamp 1676037725
transform 1 0 116472 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input118
timestamp 1676037725
transform 1 0 115736 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input119
timestamp 1676037725
transform 1 0 115000 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input120
timestamp 1676037725
transform 1 0 113988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input121
timestamp 1676037725
transform 1 0 113344 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input122
timestamp 1676037725
transform 1 0 112700 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input123
timestamp 1676037725
transform 1 0 6532 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input124
timestamp 1676037725
transform 1 0 112148 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input125
timestamp 1676037725
transform 1 0 111320 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input126
timestamp 1676037725
transform 1 0 110584 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input127
timestamp 1676037725
transform 1 0 109848 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input128
timestamp 1676037725
transform 1 0 108836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input129
timestamp 1676037725
transform 1 0 108192 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input130
timestamp 1676037725
transform 1 0 107548 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input131
timestamp 1676037725
transform 1 0 106996 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input132
timestamp 1676037725
transform 1 0 106168 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input133
timestamp 1676037725
transform 1 0 105432 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input134
timestamp 1676037725
transform 1 0 5152 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input135
timestamp 1676037725
transform 1 0 104696 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input136
timestamp 1676037725
transform 1 0 103684 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input137
timestamp 1676037725
transform 1 0 155020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input138
timestamp 1676037725
transform 1 0 154652 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input139
timestamp 1676037725
transform 1 0 154008 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input140
timestamp 1676037725
transform 1 0 153364 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input141
timestamp 1676037725
transform 1 0 152076 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input142
timestamp 1676037725
transform 1 0 151432 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input143
timestamp 1676037725
transform 1 0 150788 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input144
timestamp 1676037725
transform 1 0 149868 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input145
timestamp 1676037725
transform 1 0 4508 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input146
timestamp 1676037725
transform 1 0 17756 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input147
timestamp 1676037725
transform 1 0 149500 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input148
timestamp 1676037725
transform 1 0 148856 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input149
timestamp 1676037725
transform 1 0 148212 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input150
timestamp 1676037725
transform 1 0 146924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input151
timestamp 1676037725
transform 1 0 146280 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input152
timestamp 1676037725
transform 1 0 145636 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input153
timestamp 1676037725
transform 1 0 144716 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input154
timestamp 1676037725
transform 1 0 144348 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input155
timestamp 1676037725
transform 1 0 143704 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input156
timestamp 1676037725
transform 1 0 142784 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input157
timestamp 1676037725
transform 1 0 3956 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input158
timestamp 1676037725
transform 1 0 143060 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input159
timestamp 1676037725
transform 1 0 141772 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input160
timestamp 1676037725
transform 1 0 141128 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input161
timestamp 1676037725
transform 1 0 140484 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input162
timestamp 1676037725
transform 1 0 139196 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input163
timestamp 1676037725
transform 1 0 138552 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input164
timestamp 1676037725
transform 1 0 154928 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input165
timestamp 1676037725
transform 1 0 154652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input166
timestamp 1676037725
transform 1 0 154008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input167
timestamp 1676037725
transform 1 0 153364 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input168
timestamp 1676037725
transform 1 0 2576 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input169
timestamp 1676037725
transform 1 0 152076 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input170
timestamp 1676037725
transform 1 0 151432 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input171
timestamp 1676037725
transform 1 0 150788 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input172
timestamp 1676037725
transform 1 0 149868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input173
timestamp 1676037725
transform 1 0 149500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input174
timestamp 1676037725
transform 1 0 148856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input175
timestamp 1676037725
transform 1 0 148212 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input176
timestamp 1676037725
transform 1 0 146924 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input177
timestamp 1676037725
transform 1 0 146280 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input178
timestamp 1676037725
transform 1 0 145636 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input179
timestamp 1676037725
transform 1 0 2300 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input180
timestamp 1676037725
transform 1 0 144716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input181
timestamp 1676037725
transform 1 0 144348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input182
timestamp 1676037725
transform 1 0 143704 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input183
timestamp 1676037725
transform 1 0 143060 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input184
timestamp 1676037725
transform 1 0 141772 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input185
timestamp 1676037725
transform 1 0 141128 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input186
timestamp 1676037725
transform 1 0 140484 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input187
timestamp 1676037725
transform 1 0 139564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input188
timestamp 1676037725
transform 1 0 139196 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input189
timestamp 1676037725
transform 1 0 138552 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input190
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input191
timestamp 1676037725
transform 1 0 189428 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input192
timestamp 1676037725
transform 1 0 189428 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input193
timestamp 1676037725
transform 1 0 188140 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input194
timestamp 1676037725
transform 1 0 186944 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input195
timestamp 1676037725
transform 1 0 186852 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input196
timestamp 1676037725
transform 1 0 186852 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input197
timestamp 1676037725
transform 1 0 184736 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input198
timestamp 1676037725
transform 1 0 184276 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input199
timestamp 1676037725
transform 1 0 183264 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input200
timestamp 1676037725
transform 1 0 182528 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input201
timestamp 1676037725
transform 1 0 18492 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input202
timestamp 1676037725
transform 1 0 181792 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input203
timestamp 1676037725
transform 1 0 181700 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input204
timestamp 1676037725
transform 1 0 180412 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input205
timestamp 1676037725
transform 1 0 179584 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input206
timestamp 1676037725
transform 1 0 179124 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input207
timestamp 1676037725
transform 1 0 179124 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input208
timestamp 1676037725
transform 1 0 177836 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input209
timestamp 1676037725
transform 1 0 176640 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input210
timestamp 1676037725
transform 1 0 176548 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input211
timestamp 1676037725
transform 1 0 176548 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input212
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input213
timestamp 1676037725
transform 1 0 174432 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input214
timestamp 1676037725
transform 1 0 173972 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input215
timestamp 1676037725
transform 1 0 172960 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input216
timestamp 1676037725
transform 1 0 172224 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input217
timestamp 1676037725
transform 1 0 189428 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input218
timestamp 1676037725
transform 1 0 188416 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input219
timestamp 1676037725
transform 1 0 189428 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input220
timestamp 1676037725
transform 1 0 186944 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input221
timestamp 1676037725
transform 1 0 186852 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input222
timestamp 1676037725
transform 1 0 186852 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input223
timestamp 1676037725
transform 1 0 17020 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input224
timestamp 1676037725
transform 1 0 185564 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input225
timestamp 1676037725
transform 1 0 184276 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input226
timestamp 1676037725
transform 1 0 183264 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input227
timestamp 1676037725
transform 1 0 184276 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input228
timestamp 1676037725
transform 1 0 182160 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input229
timestamp 1676037725
transform 1 0 181700 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input230
timestamp 1676037725
transform 1 0 180872 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input231
timestamp 1676037725
transform 1 0 179584 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input232
timestamp 1676037725
transform 1 0 179124 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input233
timestamp 1676037725
transform 1 0 177744 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input234
timestamp 1676037725
transform 1 0 16008 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input235
timestamp 1676037725
transform 1 0 177376 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input236
timestamp 1676037725
transform 1 0 176640 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input237
timestamp 1676037725
transform 1 0 176548 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input238
timestamp 1676037725
transform 1 0 175720 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input239
timestamp 1676037725
transform 1 0 174432 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input240
timestamp 1676037725
transform 1 0 173972 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input241
timestamp 1676037725
transform 1 0 172960 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input242
timestamp 1676037725
transform 1 0 172224 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input243
timestamp 1676037725
transform 1 0 223836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input244
timestamp 1676037725
transform 1 0 222548 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input245
timestamp 1676037725
transform 1 0 15272 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input246
timestamp 1676037725
transform 1 0 224664 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input247
timestamp 1676037725
transform 1 0 222916 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input248
timestamp 1676037725
transform 1 0 221628 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input249
timestamp 1676037725
transform 1 0 221628 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input250
timestamp 1676037725
transform 1 0 220984 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input251
timestamp 1676037725
transform 1 0 220340 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input252
timestamp 1676037725
transform 1 0 219604 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input253
timestamp 1676037725
transform 1 0 216108 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input254
timestamp 1676037725
transform 1 0 216476 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input255
timestamp 1676037725
transform 1 0 215832 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input256
timestamp 1676037725
transform 1 0 14536 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input257
timestamp 1676037725
transform 1 0 17020 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input258
timestamp 1676037725
transform 1 0 215188 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input259
timestamp 1676037725
transform 1 0 213900 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input260
timestamp 1676037725
transform 1 0 213256 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input261
timestamp 1676037725
transform 1 0 212612 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input262
timestamp 1676037725
transform 1 0 211508 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input263
timestamp 1676037725
transform 1 0 211324 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input264
timestamp 1676037725
transform 1 0 210680 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input265
timestamp 1676037725
transform 1 0 210036 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input266
timestamp 1676037725
transform 1 0 208748 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input267
timestamp 1676037725
transform 1 0 208104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input268
timestamp 1676037725
transform 1 0 13432 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input269
timestamp 1676037725
transform 1 0 207460 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input270
timestamp 1676037725
transform 1 0 206356 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input271
timestamp 1676037725
transform 1 0 223560 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input272
timestamp 1676037725
transform 1 0 222916 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input273
timestamp 1676037725
transform 1 0 221812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input274
timestamp 1676037725
transform 1 0 221628 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input275
timestamp 1676037725
transform 1 0 220984 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input276
timestamp 1676037725
transform 1 0 220340 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input277
timestamp 1676037725
transform 1 0 219052 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input278
timestamp 1676037725
transform 1 0 218408 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input279
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input280
timestamp 1676037725
transform 1 0 217764 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input281
timestamp 1676037725
transform 1 0 216660 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input282
timestamp 1676037725
transform 1 0 216476 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input283
timestamp 1676037725
transform 1 0 215832 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input284
timestamp 1676037725
transform 1 0 215188 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input285
timestamp 1676037725
transform 1 0 213900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input286
timestamp 1676037725
transform 1 0 213256 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input287
timestamp 1676037725
transform 1 0 212612 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input288
timestamp 1676037725
transform 1 0 211508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input289
timestamp 1676037725
transform 1 0 211324 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input290
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input291
timestamp 1676037725
transform 1 0 210680 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input292
timestamp 1676037725
transform 1 0 210036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input293
timestamp 1676037725
transform 1 0 208748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input294
timestamp 1676037725
transform 1 0 208104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input295
timestamp 1676037725
transform 1 0 207460 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input296
timestamp 1676037725
transform 1 0 206356 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input297
timestamp 1676037725
transform 1 0 258980 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input298
timestamp 1676037725
transform 1 0 256680 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input299
timestamp 1676037725
transform 1 0 256404 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input300
timestamp 1676037725
transform 1 0 256404 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input301
timestamp 1676037725
transform 1 0 11868 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input302
timestamp 1676037725
transform 1 0 255116 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input303
timestamp 1676037725
transform 1 0 253828 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input304
timestamp 1676037725
transform 1 0 253828 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input305
timestamp 1676037725
transform 1 0 252264 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input306
timestamp 1676037725
transform 1 0 251528 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input307
timestamp 1676037725
transform 1 0 251252 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input308
timestamp 1676037725
transform 1 0 250056 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input309
timestamp 1676037725
transform 1 0 249964 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input310
timestamp 1676037725
transform 1 0 247848 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input311
timestamp 1676037725
transform 1 0 248676 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input312
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input313
timestamp 1676037725
transform 1 0 248676 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input314
timestamp 1676037725
transform 1 0 246376 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input315
timestamp 1676037725
transform 1 0 246100 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input316
timestamp 1676037725
transform 1 0 246100 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input317
timestamp 1676037725
transform 1 0 244812 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input318
timestamp 1676037725
transform 1 0 243432 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input319
timestamp 1676037725
transform 1 0 243524 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input320
timestamp 1676037725
transform 1 0 243524 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input321
timestamp 1676037725
transform 1 0 241224 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input322
timestamp 1676037725
transform 1 0 240948 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input323
timestamp 1676037725
transform 1 0 10396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input324
timestamp 1676037725
transform 1 0 257692 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input325
timestamp 1676037725
transform 1 0 256680 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input326
timestamp 1676037725
transform 1 0 256404 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input327
timestamp 1676037725
transform 1 0 256404 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input328
timestamp 1676037725
transform 1 0 254472 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input329
timestamp 1676037725
transform 1 0 253828 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input330
timestamp 1676037725
transform 1 0 253828 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input331
timestamp 1676037725
transform 1 0 252540 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input332
timestamp 1676037725
transform 1 0 251528 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input333
timestamp 1676037725
transform 1 0 251252 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input334
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input335
timestamp 1676037725
transform 1 0 251252 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input336
timestamp 1676037725
transform 1 0 249320 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input337
timestamp 1676037725
transform 1 0 248676 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input338
timestamp 1676037725
transform 1 0 248676 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input339
timestamp 1676037725
transform 1 0 247388 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input340
timestamp 1676037725
transform 1 0 246376 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input341
timestamp 1676037725
transform 1 0 246100 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input342
timestamp 1676037725
transform 1 0 246100 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input343
timestamp 1676037725
transform 1 0 244720 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input344
timestamp 1676037725
transform 1 0 243432 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input345
timestamp 1676037725
transform 1 0 8280 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input346
timestamp 1676037725
transform 1 0 243524 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input347
timestamp 1676037725
transform 1 0 241960 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input348
timestamp 1676037725
transform 1 0 241224 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input349
timestamp 1676037725
transform 1 0 240120 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input350
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input351
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input352
timestamp 1676037725
transform 1 0 16836 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input353
timestamp 1676037725
transform 1 0 6716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input354
timestamp 1676037725
transform 1 0 5704 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input355
timestamp 1676037725
transform 1 0 4968 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input356
timestamp 1676037725
transform 1 0 4232 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input357
timestamp 1676037725
transform 1 0 3128 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input358
timestamp 1676037725
transform 1 0 3036 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input359
timestamp 1676037725
transform 1 0 2300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input360
timestamp 1676037725
transform 1 0 1564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input361
timestamp 1676037725
transform 1 0 52164 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input362
timestamp 1676037725
transform 1 0 51520 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input363
timestamp 1676037725
transform 1 0 15548 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input364
timestamp 1676037725
transform 1 0 50876 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input365
timestamp 1676037725
transform 1 0 50416 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input366
timestamp 1676037725
transform 1 0 49588 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input367
timestamp 1676037725
transform 1 0 48944 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input368
timestamp 1676037725
transform 1 0 48208 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input369
timestamp 1676037725
transform 1 0 47012 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input370
timestamp 1676037725
transform 1 0 46368 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input371
timestamp 1676037725
transform 1 0 45724 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input372
timestamp 1676037725
transform 1 0 45264 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input373
timestamp 1676037725
transform 1 0 44436 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input374
timestamp 1676037725
transform 1 0 14812 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input375
timestamp 1676037725
transform 1 0 43792 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input376
timestamp 1676037725
transform 1 0 43056 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input377
timestamp 1676037725
transform 1 0 41860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input378
timestamp 1676037725
transform 1 0 41216 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input379
timestamp 1676037725
transform 1 0 40572 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input380
timestamp 1676037725
transform 1 0 39284 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input381
timestamp 1676037725
transform 1 0 38640 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input382
timestamp 1676037725
transform 1 0 37996 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input383
timestamp 1676037725
transform 1 0 37904 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input384
timestamp 1676037725
transform 1 0 36708 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input385
timestamp 1676037725
transform 1 0 14076 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input386
timestamp 1676037725
transform 1 0 36064 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input387
timestamp 1676037725
transform 1 0 35420 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input388
timestamp 1676037725
transform 1 0 52808 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input389
timestamp 1676037725
transform 1 0 51888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input390
timestamp 1676037725
transform 1 0 51152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input391
timestamp 1676037725
transform 1 0 50416 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input392
timestamp 1676037725
transform 1 0 49588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input393
timestamp 1676037725
transform 1 0 48944 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input394
timestamp 1676037725
transform 1 0 48208 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input395
timestamp 1676037725
transform 1 0 47012 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input396
timestamp 1676037725
transform 1 0 13340 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input397
timestamp 1676037725
transform 1 0 46368 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input398
timestamp 1676037725
transform 1 0 45724 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input399
timestamp 1676037725
transform 1 0 45264 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input400
timestamp 1676037725
transform 1 0 44436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input401
timestamp 1676037725
transform 1 0 43792 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input402
timestamp 1676037725
transform 1 0 43056 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input403
timestamp 1676037725
transform 1 0 41860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input404
timestamp 1676037725
transform 1 0 41216 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input405
timestamp 1676037725
transform 1 0 40572 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input406
timestamp 1676037725
transform 1 0 40112 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input407
timestamp 1676037725
transform 1 0 12604 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input408
timestamp 1676037725
transform 1 0 39284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input409
timestamp 1676037725
transform 1 0 38640 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input410
timestamp 1676037725
transform 1 0 37904 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input411
timestamp 1676037725
transform 1 0 36708 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input412
timestamp 1676037725
transform 1 0 36064 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input413
timestamp 1676037725
transform 1 0 35420 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input414
timestamp 1676037725
transform 1 0 86756 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input415
timestamp 1676037725
transform 1 0 86112 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input416
timestamp 1676037725
transform 1 0 85008 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input417
timestamp 1676037725
transform 1 0 82432 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input418
timestamp 1676037725
transform 1 0 11868 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 271492 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 271492 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 271492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 271492 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 271492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 271492 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 271492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 271492 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 271492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 271492 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 271492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 271492 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 271492 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 271492 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 271492 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 271492 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32 openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1676037725
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1676037725
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1676037725
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1676037725
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1676037725
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1676037725
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1676037725
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1676037725
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1676037725
transform 1 0 26864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1676037725
transform 1 0 29440 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1676037725
transform 1 0 32016 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1676037725
transform 1 0 34592 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1676037725
transform 1 0 37168 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1676037725
transform 1 0 39744 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1676037725
transform 1 0 42320 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1676037725
transform 1 0 44896 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1676037725
transform 1 0 47472 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1676037725
transform 1 0 50048 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1676037725
transform 1 0 52624 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1676037725
transform 1 0 55200 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1676037725
transform 1 0 57776 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1676037725
transform 1 0 60352 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1676037725
transform 1 0 62928 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1676037725
transform 1 0 65504 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1676037725
transform 1 0 68080 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1676037725
transform 1 0 70656 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1676037725
transform 1 0 73232 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1676037725
transform 1 0 75808 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1676037725
transform 1 0 78384 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1676037725
transform 1 0 80960 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1676037725
transform 1 0 83536 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1676037725
transform 1 0 86112 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1676037725
transform 1 0 88688 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1676037725
transform 1 0 91264 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1676037725
transform 1 0 93840 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1676037725
transform 1 0 96416 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1676037725
transform 1 0 98992 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1676037725
transform 1 0 101568 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1676037725
transform 1 0 104144 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1676037725
transform 1 0 106720 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 109296 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 111872 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 114448 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 117024 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 119600 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 122176 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 124752 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 127328 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 129904 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 132480 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 135056 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 137632 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 140208 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 142784 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 145360 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 147936 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 150512 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 153088 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 155664 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 158240 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 160816 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 163392 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 165968 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 168544 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 171120 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 173696 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 176272 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 178848 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 181424 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 184000 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 186576 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 189152 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 191728 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 194304 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 196880 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 199456 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 202032 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 204608 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 207184 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 209760 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 212336 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 214912 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 217488 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 220064 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 222640 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 225216 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 227792 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 230368 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 232944 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 235520 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 238096 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 240672 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 243248 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 245824 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 248400 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 250976 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 253552 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 256128 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 258704 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 261280 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 263856 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 266432 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 269008 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 26864 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 32016 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 37168 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 42320 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 47472 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 52624 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 57776 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 62928 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 68080 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 73232 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 78384 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 83536 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 88688 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 93840 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 98992 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 104144 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 109296 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 114448 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 119600 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 124752 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 129904 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 135056 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 140208 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 145360 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 150512 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 155664 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 160816 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 165968 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 171120 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 176272 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 181424 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 186576 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 191728 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 196880 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 202032 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 207184 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 212336 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 217488 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 222640 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 227792 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 232944 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 238096 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 243248 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 248400 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 253552 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 258704 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 263856 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 269008 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 91264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 96416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 101568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 106720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 111872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 117024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 122176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 127328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 132480 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 137632 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 142784 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 147936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 153088 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 158240 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 163392 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 168544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 173696 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 178848 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 184000 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 189152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 194304 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 199456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 204608 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 209760 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 214912 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 220064 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 225216 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 230368 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 235520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 240672 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 245824 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 250976 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 256128 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 261280 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 266432 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 88688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 93840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 98992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 104144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 109296 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 114448 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 119600 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 124752 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 129904 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 135056 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 140208 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 145360 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 150512 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 155664 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 160816 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 165968 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 171120 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 176272 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 181424 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 186576 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 191728 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 196880 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 202032 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 207184 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 212336 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 217488 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 222640 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 227792 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 232944 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 238096 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 243248 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 248400 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 253552 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 258704 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 263856 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 269008 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 91264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 96416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 101568 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 106720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 111872 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 117024 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 122176 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 127328 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 132480 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 137632 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 142784 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 147936 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 153088 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 158240 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 163392 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 168544 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 173696 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 178848 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 184000 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 189152 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 194304 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 199456 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 204608 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 209760 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 214912 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 220064 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 225216 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 230368 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 235520 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 240672 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 245824 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 250976 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 256128 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 261280 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 266432 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 88688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 93840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 98992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 104144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 109296 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 114448 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 119600 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 124752 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 129904 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 135056 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 140208 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 145360 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 150512 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 155664 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 160816 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 165968 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 171120 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 176272 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 181424 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 186576 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 191728 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 196880 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 202032 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 207184 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 212336 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 217488 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 222640 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 227792 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 232944 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 238096 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 243248 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 248400 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 253552 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 258704 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 263856 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 269008 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 91264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 96416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 101568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 106720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 111872 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 117024 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 122176 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 127328 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 132480 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 137632 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 142784 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 147936 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 153088 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 158240 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 163392 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 168544 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 173696 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 178848 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 184000 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 189152 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 194304 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 199456 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 204608 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 209760 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 214912 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 220064 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 225216 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 230368 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 235520 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 240672 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 245824 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 250976 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 256128 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 261280 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 266432 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 88688 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 93840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 98992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 104144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 109296 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 114448 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 119600 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 124752 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 129904 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 135056 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 140208 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 145360 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 150512 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 155664 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 160816 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 165968 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 171120 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 176272 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 181424 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 186576 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 191728 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 196880 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 202032 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 207184 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 212336 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 217488 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 222640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 227792 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 232944 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 238096 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 243248 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 248400 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 253552 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 258704 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 263856 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 269008 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 91264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 96416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 101568 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 106720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 111872 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 117024 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 122176 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 127328 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 132480 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 137632 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 142784 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 147936 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 153088 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 158240 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 163392 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 168544 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 173696 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 178848 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 184000 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 189152 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 194304 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 199456 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 204608 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 209760 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 214912 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 220064 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 225216 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 230368 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 235520 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 240672 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 245824 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 250976 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 256128 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 261280 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 266432 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 83536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 88688 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 93840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 98992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 104144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 109296 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 114448 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 119600 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 124752 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 129904 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 135056 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 140208 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 145360 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 150512 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 155664 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 160816 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 165968 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 171120 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 176272 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 181424 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 186576 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 191728 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 196880 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 202032 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 207184 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 212336 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 217488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 222640 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 227792 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 232944 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 238096 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 243248 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 248400 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 253552 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 258704 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 263856 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 269008 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 86112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 91264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 96416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 101568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 106720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 111872 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 117024 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 122176 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 127328 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 132480 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 137632 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 142784 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 147936 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1676037725
transform 1 0 153088 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1676037725
transform 1 0 158240 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1676037725
transform 1 0 163392 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1676037725
transform 1 0 168544 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1676037725
transform 1 0 173696 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1676037725
transform 1 0 178848 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1676037725
transform 1 0 184000 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1676037725
transform 1 0 189152 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1676037725
transform 1 0 194304 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1676037725
transform 1 0 199456 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1676037725
transform 1 0 204608 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1676037725
transform 1 0 209760 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1676037725
transform 1 0 214912 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1676037725
transform 1 0 220064 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1676037725
transform 1 0 225216 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1676037725
transform 1 0 230368 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1676037725
transform 1 0 235520 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1676037725
transform 1 0 240672 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1676037725
transform 1 0 245824 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1676037725
transform 1 0 250976 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1676037725
transform 1 0 256128 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1676037725
transform 1 0 261280 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1676037725
transform 1 0 266432 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1676037725
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1676037725
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1676037725
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1676037725
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1676037725
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1676037725
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1676037725
transform 1 0 83536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1676037725
transform 1 0 88688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1676037725
transform 1 0 93840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1676037725
transform 1 0 98992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1676037725
transform 1 0 104144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1676037725
transform 1 0 109296 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1676037725
transform 1 0 114448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1676037725
transform 1 0 119600 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1676037725
transform 1 0 124752 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1676037725
transform 1 0 129904 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1676037725
transform 1 0 135056 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1676037725
transform 1 0 140208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1676037725
transform 1 0 145360 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1676037725
transform 1 0 150512 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1676037725
transform 1 0 155664 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1676037725
transform 1 0 160816 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1676037725
transform 1 0 165968 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1676037725
transform 1 0 171120 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1676037725
transform 1 0 176272 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1676037725
transform 1 0 181424 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1676037725
transform 1 0 186576 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1676037725
transform 1 0 191728 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1676037725
transform 1 0 196880 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1676037725
transform 1 0 202032 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1676037725
transform 1 0 207184 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1676037725
transform 1 0 212336 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1676037725
transform 1 0 217488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1676037725
transform 1 0 222640 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1676037725
transform 1 0 227792 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1676037725
transform 1 0 232944 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1676037725
transform 1 0 238096 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1676037725
transform 1 0 243248 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1676037725
transform 1 0 248400 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1676037725
transform 1 0 253552 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1676037725
transform 1 0 258704 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1676037725
transform 1 0 263856 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1676037725
transform 1 0 269008 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1676037725
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1676037725
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1676037725
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1676037725
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1676037725
transform 1 0 70656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1676037725
transform 1 0 75808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1676037725
transform 1 0 80960 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1676037725
transform 1 0 86112 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1676037725
transform 1 0 91264 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1676037725
transform 1 0 96416 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1676037725
transform 1 0 101568 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1676037725
transform 1 0 106720 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1676037725
transform 1 0 111872 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1676037725
transform 1 0 117024 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1676037725
transform 1 0 122176 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1676037725
transform 1 0 127328 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1676037725
transform 1 0 132480 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1676037725
transform 1 0 137632 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1676037725
transform 1 0 142784 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1676037725
transform 1 0 147936 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1676037725
transform 1 0 153088 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1676037725
transform 1 0 158240 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1676037725
transform 1 0 163392 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1676037725
transform 1 0 168544 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1676037725
transform 1 0 173696 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1676037725
transform 1 0 178848 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1676037725
transform 1 0 184000 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1676037725
transform 1 0 189152 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1676037725
transform 1 0 194304 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1676037725
transform 1 0 199456 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1676037725
transform 1 0 204608 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1676037725
transform 1 0 209760 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1676037725
transform 1 0 214912 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1676037725
transform 1 0 220064 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1676037725
transform 1 0 225216 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1676037725
transform 1 0 230368 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1676037725
transform 1 0 235520 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1676037725
transform 1 0 240672 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1676037725
transform 1 0 245824 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1676037725
transform 1 0 250976 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1676037725
transform 1 0 256128 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1676037725
transform 1 0 261280 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1676037725
transform 1 0 266432 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1676037725
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1676037725
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1676037725
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1676037725
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1676037725
transform 1 0 73232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1676037725
transform 1 0 78384 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1676037725
transform 1 0 83536 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1676037725
transform 1 0 88688 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1676037725
transform 1 0 93840 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1676037725
transform 1 0 98992 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1676037725
transform 1 0 104144 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1676037725
transform 1 0 109296 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1676037725
transform 1 0 114448 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1676037725
transform 1 0 119600 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1676037725
transform 1 0 124752 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1676037725
transform 1 0 129904 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1676037725
transform 1 0 135056 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1676037725
transform 1 0 140208 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1676037725
transform 1 0 145360 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1676037725
transform 1 0 150512 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1676037725
transform 1 0 155664 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1676037725
transform 1 0 160816 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1676037725
transform 1 0 165968 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1676037725
transform 1 0 171120 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1676037725
transform 1 0 176272 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1676037725
transform 1 0 181424 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1676037725
transform 1 0 186576 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1676037725
transform 1 0 191728 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1676037725
transform 1 0 196880 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1676037725
transform 1 0 202032 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1676037725
transform 1 0 207184 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1676037725
transform 1 0 212336 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1676037725
transform 1 0 217488 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1676037725
transform 1 0 222640 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1676037725
transform 1 0 227792 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1676037725
transform 1 0 232944 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1676037725
transform 1 0 238096 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1676037725
transform 1 0 243248 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1676037725
transform 1 0 248400 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1676037725
transform 1 0 253552 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1676037725
transform 1 0 258704 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1676037725
transform 1 0 263856 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1676037725
transform 1 0 269008 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1676037725
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1676037725
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1676037725
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1676037725
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1676037725
transform 1 0 70656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1676037725
transform 1 0 75808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1676037725
transform 1 0 80960 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1676037725
transform 1 0 86112 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1676037725
transform 1 0 91264 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1676037725
transform 1 0 96416 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1676037725
transform 1 0 101568 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1676037725
transform 1 0 106720 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1676037725
transform 1 0 111872 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1676037725
transform 1 0 117024 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1676037725
transform 1 0 122176 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1676037725
transform 1 0 127328 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1676037725
transform 1 0 132480 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1676037725
transform 1 0 137632 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1676037725
transform 1 0 142784 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1676037725
transform 1 0 147936 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1676037725
transform 1 0 153088 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1676037725
transform 1 0 158240 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1676037725
transform 1 0 163392 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1676037725
transform 1 0 168544 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1676037725
transform 1 0 173696 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1676037725
transform 1 0 178848 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1676037725
transform 1 0 184000 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1676037725
transform 1 0 189152 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1676037725
transform 1 0 194304 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1676037725
transform 1 0 199456 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1676037725
transform 1 0 204608 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1676037725
transform 1 0 209760 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1676037725
transform 1 0 214912 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1676037725
transform 1 0 220064 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1676037725
transform 1 0 225216 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1676037725
transform 1 0 230368 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1676037725
transform 1 0 235520 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1676037725
transform 1 0 240672 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1676037725
transform 1 0 245824 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1676037725
transform 1 0 250976 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1676037725
transform 1 0 256128 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1676037725
transform 1 0 261280 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1676037725
transform 1 0 266432 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1676037725
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1676037725
transform 1 0 8832 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1676037725
transform 1 0 13984 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1676037725
transform 1 0 19136 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1676037725
transform 1 0 24288 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1676037725
transform 1 0 29440 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1676037725
transform 1 0 34592 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1676037725
transform 1 0 39744 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1676037725
transform 1 0 44896 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1676037725
transform 1 0 50048 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1676037725
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1676037725
transform 1 0 55200 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1676037725
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1676037725
transform 1 0 60352 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1676037725
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1676037725
transform 1 0 65504 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1676037725
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1676037725
transform 1 0 70656 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1676037725
transform 1 0 73232 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1676037725
transform 1 0 75808 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1676037725
transform 1 0 78384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1676037725
transform 1 0 80960 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1676037725
transform 1 0 83536 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1676037725
transform 1 0 86112 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1676037725
transform 1 0 88688 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1676037725
transform 1 0 91264 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1676037725
transform 1 0 93840 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1676037725
transform 1 0 96416 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1676037725
transform 1 0 98992 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1676037725
transform 1 0 101568 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1676037725
transform 1 0 104144 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1676037725
transform 1 0 106720 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1676037725
transform 1 0 109296 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1676037725
transform 1 0 111872 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1676037725
transform 1 0 114448 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1676037725
transform 1 0 117024 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1676037725
transform 1 0 119600 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1676037725
transform 1 0 122176 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1676037725
transform 1 0 124752 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1676037725
transform 1 0 127328 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1676037725
transform 1 0 129904 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1676037725
transform 1 0 132480 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1676037725
transform 1 0 135056 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1676037725
transform 1 0 137632 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1676037725
transform 1 0 140208 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1676037725
transform 1 0 142784 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1676037725
transform 1 0 145360 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1676037725
transform 1 0 147936 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1676037725
transform 1 0 150512 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1676037725
transform 1 0 153088 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1676037725
transform 1 0 155664 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1676037725
transform 1 0 158240 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1676037725
transform 1 0 160816 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1676037725
transform 1 0 163392 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1676037725
transform 1 0 165968 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1676037725
transform 1 0 168544 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1676037725
transform 1 0 171120 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1676037725
transform 1 0 173696 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1676037725
transform 1 0 176272 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1676037725
transform 1 0 178848 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1676037725
transform 1 0 181424 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1676037725
transform 1 0 184000 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1676037725
transform 1 0 186576 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1676037725
transform 1 0 189152 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1676037725
transform 1 0 191728 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1676037725
transform 1 0 194304 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1676037725
transform 1 0 196880 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1676037725
transform 1 0 199456 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1676037725
transform 1 0 202032 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1676037725
transform 1 0 204608 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1676037725
transform 1 0 207184 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1676037725
transform 1 0 209760 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1676037725
transform 1 0 212336 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1676037725
transform 1 0 214912 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1676037725
transform 1 0 217488 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1676037725
transform 1 0 220064 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1676037725
transform 1 0 222640 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1676037725
transform 1 0 225216 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1676037725
transform 1 0 227792 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1676037725
transform 1 0 230368 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1676037725
transform 1 0 232944 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1676037725
transform 1 0 235520 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1676037725
transform 1 0 238096 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1676037725
transform 1 0 240672 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1676037725
transform 1 0 243248 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1676037725
transform 1 0 245824 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1676037725
transform 1 0 248400 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1676037725
transform 1 0 250976 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1676037725
transform 1 0 253552 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1676037725
transform 1 0 256128 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1676037725
transform 1 0 258704 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1676037725
transform 1 0 261280 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1676037725
transform 1 0 263856 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1676037725
transform 1 0 266432 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1676037725
transform 1 0 269008 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  tbuf_row_ena_I.cell0_I openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 238556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  tbuf_spine_ow_I\[0\].cell0_I openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 243892 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  tbuf_spine_ow_I\[1\].cell0_I
timestamp 1676037725
transform 1 0 242604 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  tbuf_spine_ow_I\[2\].cell0_I
timestamp 1676037725
transform 1 0 240948 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  tbuf_spine_ow_I\[3\].cell0_I
timestamp 1676037725
transform 1 0 239016 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  tbuf_spine_ow_I\[4\].cell0_I openmpw/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 251896 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  tbuf_spine_ow_I\[5\].cell0_I
timestamp 1676037725
transform 1 0 253828 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  tbuf_spine_ow_I\[6\].cell0_I
timestamp 1676037725
transform 1 0 254288 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  tbuf_spine_ow_I\[7\].cell0_I
timestamp 1676037725
transform 1 0 256496 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  tbuf_spine_ow_I\[8\].cell0_I
timestamp 1676037725
transform 1 0 257048 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  tbuf_spine_ow_I\[9\].cell0_I
timestamp 1676037725
transform 1 0 251252 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  tbuf_spine_ow_I\[10\].cell0_I
timestamp 1676037725
transform 1 0 259624 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  tbuf_spine_ow_I\[11\].cell0_I
timestamp 1676037725
transform 1 0 257600 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  tbuf_spine_ow_I\[12\].cell0_I
timestamp 1676037725
transform 1 0 258152 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  tbuf_spine_ow_I\[13\].cell0_I
timestamp 1676037725
transform 1 0 221536 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  tbuf_spine_ow_I\[14\].cell0_I
timestamp 1676037725
transform 1 0 218868 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  tbuf_spine_ow_I\[15\].cell0_I
timestamp 1676037725
transform 1 0 216016 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  tbuf_spine_ow_I\[16\].cell0_I
timestamp 1676037725
transform 1 0 217764 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  tbuf_spine_ow_I\[17\].cell0_I
timestamp 1676037725
transform 1 0 217304 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  tbuf_spine_ow_I\[18\].cell0_I
timestamp 1676037725
transform 1 0 217764 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  tbuf_spine_ow_I\[19\].cell0_I
timestamp 1676037725
transform 1 0 218592 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  tbuf_spine_ow_I\[20\].cell0_I
timestamp 1676037725
transform 1 0 225860 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  tbuf_spine_ow_I\[21\].cell0_I
timestamp 1676037725
transform 1 0 220800 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  tbuf_spine_ow_I\[22\].cell0_I
timestamp 1676037725
transform 1 0 221904 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  tbuf_spine_ow_I\[23\].cell0_I
timestamp 1676037725
transform 1 0 223008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  tt_mux_517
timestamp 1676037725
transform 1 0 260820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_518
timestamp 1676037725
transform 1 0 265972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_519
timestamp 1676037725
transform 1 0 265328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_520
timestamp 1676037725
transform 1 0 1564 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_521
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_522
timestamp 1676037725
transform 1 0 34132 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_523
timestamp 1676037725
transform 1 0 34960 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_524
timestamp 1676037725
transform 1 0 68908 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_525
timestamp 1676037725
transform 1 0 68908 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_526
timestamp 1676037725
transform 1 0 103040 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_527
timestamp 1676037725
transform 1 0 103040 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_528
timestamp 1676037725
transform 1 0 137908 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_529
timestamp 1676037725
transform 1 0 137908 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_530
timestamp 1676037725
transform 1 0 171488 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_531
timestamp 1676037725
transform 1 0 171488 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_532
timestamp 1676037725
transform 1 0 205620 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_533
timestamp 1676037725
transform 1 0 205620 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_534
timestamp 1676037725
transform 1 0 239752 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_535
timestamp 1676037725
transform 1 0 239476 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_mux_552
timestamp 1676037725
transform 1 0 260176 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_ena_I.genblk1.cell0_I
timestamp 1676037725
transform 1 0 238372 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_8  zbuf_bus_ena_I.genblk1.cell1_I
timestamp 1676037725
transform 1 0 230920 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 270480 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[0\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 267996 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 269284 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[1\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 269284 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 269284 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[2\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 268272 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 268272 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[3\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 267720 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 269468 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[4\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 266708 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[5\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 270480 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[5\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 266524 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[6\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 267168 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[6\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 265328 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[7\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 269284 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[7\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 264132 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[8\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 270112 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[8\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 263948 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[9\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 270296 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[9\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 262844 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[10\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 266708 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[10\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 262752 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[11\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 265144 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[11\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 261096 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[12\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 262292 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[12\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 261556 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[13\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 261464 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[13\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 260268 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[14\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 264500 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[14\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 260084 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[15\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 265880 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[15\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 258888 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[16\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 265788 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[16\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 263672 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_iw_I\[17\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 268364 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_iw_I\[17\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 268088 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_sel_I\[0\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 237728 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_sel_I\[0\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 231104 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_sel_I\[1\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 235244 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_sel_I\[1\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 231196 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_sel_I\[2\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 237268 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_sel_I\[2\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 235612 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_sel_I\[3\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 236992 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_sel_I\[3\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 236072 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  zbuf_bus_sel_I\[4\].genblk1.cell0_I
timestamp 1676037725
transform 1 0 236900 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  zbuf_bus_sel_I\[4\].genblk1.cell1_I
timestamp 1676037725
transform 1 0 236072 0 -1 7616
box -38 -48 866 592
<< labels >>
flabel metal3 s 272304 9558 272504 9618 0 FreeSans 480 0 0 0 addr[0]
port 0 nsew signal input
flabel metal3 s 272304 9422 272504 9482 0 FreeSans 480 0 0 0 addr[1]
port 1 nsew signal input
flabel metal3 s 272304 9286 272504 9346 0 FreeSans 480 0 0 0 addr[2]
port 2 nsew signal input
flabel metal3 s 272304 9150 272504 9210 0 FreeSans 480 0 0 0 addr[3]
port 3 nsew signal input
flabel metal3 s 272304 9014 272504 9074 0 FreeSans 480 0 0 0 addr[4]
port 4 nsew signal input
flabel metal3 s 272304 8878 272504 8938 0 FreeSans 480 0 0 0 k_one
port 5 nsew signal tristate
flabel metal3 s 272304 8742 272504 8802 0 FreeSans 480 0 0 0 k_zero
port 6 nsew signal tristate
flabel metal3 s 272304 8606 272504 8666 0 FreeSans 480 0 0 0 spine_iw[0]
port 7 nsew signal input
flabel metal3 s 272304 7246 272504 7306 0 FreeSans 480 0 0 0 spine_iw[10]
port 8 nsew signal input
flabel metal3 s 272304 7110 272504 7170 0 FreeSans 480 0 0 0 spine_iw[11]
port 9 nsew signal input
flabel metal3 s 272304 6974 272504 7034 0 FreeSans 480 0 0 0 spine_iw[12]
port 10 nsew signal input
flabel metal3 s 272304 6838 272504 6898 0 FreeSans 480 0 0 0 spine_iw[13]
port 11 nsew signal input
flabel metal3 s 272304 6702 272504 6762 0 FreeSans 480 0 0 0 spine_iw[14]
port 12 nsew signal input
flabel metal3 s 272304 6566 272504 6626 0 FreeSans 480 0 0 0 spine_iw[15]
port 13 nsew signal input
flabel metal3 s 272304 6430 272504 6490 0 FreeSans 480 0 0 0 spine_iw[16]
port 14 nsew signal input
flabel metal3 s 272304 6294 272504 6354 0 FreeSans 480 0 0 0 spine_iw[17]
port 15 nsew signal input
flabel metal3 s 272304 6158 272504 6218 0 FreeSans 480 0 0 0 spine_iw[18]
port 16 nsew signal input
flabel metal3 s 272304 6022 272504 6082 0 FreeSans 480 0 0 0 spine_iw[19]
port 17 nsew signal input
flabel metal3 s 272304 8470 272504 8530 0 FreeSans 480 0 0 0 spine_iw[1]
port 18 nsew signal input
flabel metal3 s 272304 5886 272504 5946 0 FreeSans 480 0 0 0 spine_iw[20]
port 19 nsew signal input
flabel metal3 s 272304 5750 272504 5810 0 FreeSans 480 0 0 0 spine_iw[21]
port 20 nsew signal input
flabel metal3 s 272304 5614 272504 5674 0 FreeSans 480 0 0 0 spine_iw[22]
port 21 nsew signal input
flabel metal3 s 272304 5478 272504 5538 0 FreeSans 480 0 0 0 spine_iw[23]
port 22 nsew signal input
flabel metal3 s 272304 5342 272504 5402 0 FreeSans 480 0 0 0 spine_iw[24]
port 23 nsew signal input
flabel metal3 s 272304 5206 272504 5266 0 FreeSans 480 0 0 0 spine_iw[25]
port 24 nsew signal input
flabel metal3 s 272304 5070 272504 5130 0 FreeSans 480 0 0 0 spine_iw[26]
port 25 nsew signal input
flabel metal3 s 272304 4934 272504 4994 0 FreeSans 480 0 0 0 spine_iw[27]
port 26 nsew signal input
flabel metal3 s 272304 4798 272504 4858 0 FreeSans 480 0 0 0 spine_iw[28]
port 27 nsew signal input
flabel metal3 s 272304 4662 272504 4722 0 FreeSans 480 0 0 0 spine_iw[29]
port 28 nsew signal input
flabel metal3 s 272304 8334 272504 8394 0 FreeSans 480 0 0 0 spine_iw[2]
port 29 nsew signal input
flabel metal3 s 272304 4526 272504 4586 0 FreeSans 480 0 0 0 spine_iw[30]
port 30 nsew signal input
flabel metal3 s 272304 8198 272504 8258 0 FreeSans 480 0 0 0 spine_iw[3]
port 31 nsew signal input
flabel metal3 s 272304 8062 272504 8122 0 FreeSans 480 0 0 0 spine_iw[4]
port 32 nsew signal input
flabel metal3 s 272304 7926 272504 7986 0 FreeSans 480 0 0 0 spine_iw[5]
port 33 nsew signal input
flabel metal3 s 272304 7790 272504 7850 0 FreeSans 480 0 0 0 spine_iw[6]
port 34 nsew signal input
flabel metal3 s 272304 7654 272504 7714 0 FreeSans 480 0 0 0 spine_iw[7]
port 35 nsew signal input
flabel metal3 s 272304 7518 272504 7578 0 FreeSans 480 0 0 0 spine_iw[8]
port 36 nsew signal input
flabel metal3 s 272304 7382 272504 7442 0 FreeSans 480 0 0 0 spine_iw[9]
port 37 nsew signal input
flabel metal3 s 272304 4390 272504 4450 0 FreeSans 480 0 0 0 spine_ow[0]
port 38 nsew signal tristate
flabel metal3 s 272304 3030 272504 3090 0 FreeSans 480 0 0 0 spine_ow[10]
port 39 nsew signal tristate
flabel metal3 s 272304 2894 272504 2954 0 FreeSans 480 0 0 0 spine_ow[11]
port 40 nsew signal tristate
flabel metal3 s 272304 2758 272504 2818 0 FreeSans 480 0 0 0 spine_ow[12]
port 41 nsew signal tristate
flabel metal3 s 272304 2622 272504 2682 0 FreeSans 480 0 0 0 spine_ow[13]
port 42 nsew signal tristate
flabel metal3 s 272304 2486 272504 2546 0 FreeSans 480 0 0 0 spine_ow[14]
port 43 nsew signal tristate
flabel metal3 s 272304 2350 272504 2410 0 FreeSans 480 0 0 0 spine_ow[15]
port 44 nsew signal tristate
flabel metal3 s 272304 2214 272504 2274 0 FreeSans 480 0 0 0 spine_ow[16]
port 45 nsew signal tristate
flabel metal3 s 272304 2078 272504 2138 0 FreeSans 480 0 0 0 spine_ow[17]
port 46 nsew signal tristate
flabel metal3 s 272304 1942 272504 2002 0 FreeSans 480 0 0 0 spine_ow[18]
port 47 nsew signal tristate
flabel metal3 s 272304 1806 272504 1866 0 FreeSans 480 0 0 0 spine_ow[19]
port 48 nsew signal tristate
flabel metal3 s 272304 4254 272504 4314 0 FreeSans 480 0 0 0 spine_ow[1]
port 49 nsew signal tristate
flabel metal3 s 272304 1670 272504 1730 0 FreeSans 480 0 0 0 spine_ow[20]
port 50 nsew signal tristate
flabel metal3 s 272304 1534 272504 1594 0 FreeSans 480 0 0 0 spine_ow[21]
port 51 nsew signal tristate
flabel metal3 s 272304 1398 272504 1458 0 FreeSans 480 0 0 0 spine_ow[22]
port 52 nsew signal tristate
flabel metal3 s 272304 1262 272504 1322 0 FreeSans 480 0 0 0 spine_ow[23]
port 53 nsew signal tristate
flabel metal3 s 272304 1126 272504 1186 0 FreeSans 480 0 0 0 spine_ow[24]
port 54 nsew signal tristate
flabel metal3 s 272304 990 272504 1050 0 FreeSans 480 0 0 0 spine_ow[25]
port 55 nsew signal tristate
flabel metal3 s 272304 4118 272504 4178 0 FreeSans 480 0 0 0 spine_ow[2]
port 56 nsew signal tristate
flabel metal3 s 272304 3982 272504 4042 0 FreeSans 480 0 0 0 spine_ow[3]
port 57 nsew signal tristate
flabel metal3 s 272304 3846 272504 3906 0 FreeSans 480 0 0 0 spine_ow[4]
port 58 nsew signal tristate
flabel metal3 s 272304 3710 272504 3770 0 FreeSans 480 0 0 0 spine_ow[5]
port 59 nsew signal tristate
flabel metal3 s 272304 3574 272504 3634 0 FreeSans 480 0 0 0 spine_ow[6]
port 60 nsew signal tristate
flabel metal3 s 272304 3438 272504 3498 0 FreeSans 480 0 0 0 spine_ow[7]
port 61 nsew signal tristate
flabel metal3 s 272304 3302 272504 3362 0 FreeSans 480 0 0 0 spine_ow[8]
port 62 nsew signal tristate
flabel metal3 s 272304 3166 272504 3226 0 FreeSans 480 0 0 0 spine_ow[9]
port 63 nsew signal tristate
flabel metal4 s 32446 0 32506 200 0 FreeSans 480 90 0 0 um_ena[0]
port 64 nsew signal tristate
flabel metal4 s 203106 0 203166 200 0 FreeSans 480 90 0 0 um_ena[10]
port 65 nsew signal tristate
flabel metal4 s 203106 10680 203166 10880 0 FreeSans 480 90 0 0 um_ena[11]
port 66 nsew signal tristate
flabel metal4 s 237238 0 237298 200 0 FreeSans 480 90 0 0 um_ena[12]
port 67 nsew signal tristate
flabel metal4 s 237238 10680 237298 10880 0 FreeSans 480 90 0 0 um_ena[13]
port 68 nsew signal tristate
flabel metal4 s 271370 0 271430 200 0 FreeSans 480 90 0 0 um_ena[14]
port 69 nsew signal tristate
flabel metal4 s 271370 10680 271430 10880 0 FreeSans 480 90 0 0 um_ena[15]
port 70 nsew signal tristate
flabel metal4 s 32446 10680 32506 10880 0 FreeSans 480 90 0 0 um_ena[1]
port 71 nsew signal tristate
flabel metal4 s 66578 0 66638 200 0 FreeSans 480 90 0 0 um_ena[2]
port 72 nsew signal tristate
flabel metal4 s 66578 10680 66638 10880 0 FreeSans 480 90 0 0 um_ena[3]
port 73 nsew signal tristate
flabel metal4 s 100710 0 100770 200 0 FreeSans 480 90 0 0 um_ena[4]
port 74 nsew signal tristate
flabel metal4 s 100710 10680 100770 10880 0 FreeSans 480 90 0 0 um_ena[5]
port 75 nsew signal tristate
flabel metal4 s 134842 0 134902 200 0 FreeSans 480 90 0 0 um_ena[6]
port 76 nsew signal tristate
flabel metal4 s 134842 10680 134902 10880 0 FreeSans 480 90 0 0 um_ena[7]
port 77 nsew signal tristate
flabel metal4 s 168974 0 169034 200 0 FreeSans 480 90 0 0 um_ena[8]
port 78 nsew signal tristate
flabel metal4 s 168974 10680 169034 10880 0 FreeSans 480 90 0 0 um_ena[9]
port 79 nsew signal tristate
flabel metal4 s 31710 0 31770 200 0 FreeSans 480 90 0 0 um_iw[0]
port 80 nsew signal tristate
flabel metal4 s 92614 10680 92674 10880 0 FreeSans 480 90 0 0 um_iw[100]
port 81 nsew signal tristate
flabel metal4 s 91878 10680 91938 10880 0 FreeSans 480 90 0 0 um_iw[101]
port 82 nsew signal tristate
flabel metal4 s 91142 10680 91202 10880 0 FreeSans 480 90 0 0 um_iw[102]
port 83 nsew signal tristate
flabel metal4 s 90406 10680 90466 10880 0 FreeSans 480 90 0 0 um_iw[103]
port 84 nsew signal tristate
flabel metal4 s 89670 10680 89730 10880 0 FreeSans 480 90 0 0 um_iw[104]
port 85 nsew signal tristate
flabel metal4 s 88934 10680 88994 10880 0 FreeSans 480 90 0 0 um_iw[105]
port 86 nsew signal tristate
flabel metal4 s 88198 10680 88258 10880 0 FreeSans 480 90 0 0 um_iw[106]
port 87 nsew signal tristate
flabel metal4 s 87462 10680 87522 10880 0 FreeSans 480 90 0 0 um_iw[107]
port 88 nsew signal tristate
flabel metal4 s 134106 0 134166 200 0 FreeSans 480 90 0 0 um_iw[108]
port 89 nsew signal tristate
flabel metal4 s 133370 0 133430 200 0 FreeSans 480 90 0 0 um_iw[109]
port 90 nsew signal tristate
flabel metal4 s 24350 0 24410 200 0 FreeSans 480 90 0 0 um_iw[10]
port 91 nsew signal tristate
flabel metal4 s 132634 0 132694 200 0 FreeSans 480 90 0 0 um_iw[110]
port 92 nsew signal tristate
flabel metal4 s 131898 0 131958 200 0 FreeSans 480 90 0 0 um_iw[111]
port 93 nsew signal tristate
flabel metal4 s 131162 0 131222 200 0 FreeSans 480 90 0 0 um_iw[112]
port 94 nsew signal tristate
flabel metal4 s 130426 0 130486 200 0 FreeSans 480 90 0 0 um_iw[113]
port 95 nsew signal tristate
flabel metal4 s 129690 0 129750 200 0 FreeSans 480 90 0 0 um_iw[114]
port 96 nsew signal tristate
flabel metal4 s 128954 0 129014 200 0 FreeSans 480 90 0 0 um_iw[115]
port 97 nsew signal tristate
flabel metal4 s 128218 0 128278 200 0 FreeSans 480 90 0 0 um_iw[116]
port 98 nsew signal tristate
flabel metal4 s 127482 0 127542 200 0 FreeSans 480 90 0 0 um_iw[117]
port 99 nsew signal tristate
flabel metal4 s 126746 0 126806 200 0 FreeSans 480 90 0 0 um_iw[118]
port 100 nsew signal tristate
flabel metal4 s 126010 0 126070 200 0 FreeSans 480 90 0 0 um_iw[119]
port 101 nsew signal tristate
flabel metal4 s 23614 0 23674 200 0 FreeSans 480 90 0 0 um_iw[11]
port 102 nsew signal tristate
flabel metal4 s 125274 0 125334 200 0 FreeSans 480 90 0 0 um_iw[120]
port 103 nsew signal tristate
flabel metal4 s 124538 0 124598 200 0 FreeSans 480 90 0 0 um_iw[121]
port 104 nsew signal tristate
flabel metal4 s 123802 0 123862 200 0 FreeSans 480 90 0 0 um_iw[122]
port 105 nsew signal tristate
flabel metal4 s 123066 0 123126 200 0 FreeSans 480 90 0 0 um_iw[123]
port 106 nsew signal tristate
flabel metal4 s 122330 0 122390 200 0 FreeSans 480 90 0 0 um_iw[124]
port 107 nsew signal tristate
flabel metal4 s 121594 0 121654 200 0 FreeSans 480 90 0 0 um_iw[125]
port 108 nsew signal tristate
flabel metal4 s 134106 10680 134166 10880 0 FreeSans 480 90 0 0 um_iw[126]
port 109 nsew signal tristate
flabel metal4 s 133370 10680 133430 10880 0 FreeSans 480 90 0 0 um_iw[127]
port 110 nsew signal tristate
flabel metal4 s 132634 10680 132694 10880 0 FreeSans 480 90 0 0 um_iw[128]
port 111 nsew signal tristate
flabel metal4 s 131898 10680 131958 10880 0 FreeSans 480 90 0 0 um_iw[129]
port 112 nsew signal tristate
flabel metal4 s 22878 0 22938 200 0 FreeSans 480 90 0 0 um_iw[12]
port 113 nsew signal tristate
flabel metal4 s 131162 10680 131222 10880 0 FreeSans 480 90 0 0 um_iw[130]
port 114 nsew signal tristate
flabel metal4 s 130426 10680 130486 10880 0 FreeSans 480 90 0 0 um_iw[131]
port 115 nsew signal tristate
flabel metal4 s 129690 10680 129750 10880 0 FreeSans 480 90 0 0 um_iw[132]
port 116 nsew signal tristate
flabel metal4 s 128954 10680 129014 10880 0 FreeSans 480 90 0 0 um_iw[133]
port 117 nsew signal tristate
flabel metal4 s 128218 10680 128278 10880 0 FreeSans 480 90 0 0 um_iw[134]
port 118 nsew signal tristate
flabel metal4 s 127482 10680 127542 10880 0 FreeSans 480 90 0 0 um_iw[135]
port 119 nsew signal tristate
flabel metal4 s 126746 10680 126806 10880 0 FreeSans 480 90 0 0 um_iw[136]
port 120 nsew signal tristate
flabel metal4 s 126010 10680 126070 10880 0 FreeSans 480 90 0 0 um_iw[137]
port 121 nsew signal tristate
flabel metal4 s 125274 10680 125334 10880 0 FreeSans 480 90 0 0 um_iw[138]
port 122 nsew signal tristate
flabel metal4 s 124538 10680 124598 10880 0 FreeSans 480 90 0 0 um_iw[139]
port 123 nsew signal tristate
flabel metal4 s 22142 0 22202 200 0 FreeSans 480 90 0 0 um_iw[13]
port 124 nsew signal tristate
flabel metal4 s 123802 10680 123862 10880 0 FreeSans 480 90 0 0 um_iw[140]
port 125 nsew signal tristate
flabel metal4 s 123066 10680 123126 10880 0 FreeSans 480 90 0 0 um_iw[141]
port 126 nsew signal tristate
flabel metal4 s 122330 10680 122390 10880 0 FreeSans 480 90 0 0 um_iw[142]
port 127 nsew signal tristate
flabel metal4 s 121594 10680 121654 10880 0 FreeSans 480 90 0 0 um_iw[143]
port 128 nsew signal tristate
flabel metal4 s 168238 0 168298 200 0 FreeSans 480 90 0 0 um_iw[144]
port 129 nsew signal tristate
flabel metal4 s 167502 0 167562 200 0 FreeSans 480 90 0 0 um_iw[145]
port 130 nsew signal tristate
flabel metal4 s 166766 0 166826 200 0 FreeSans 480 90 0 0 um_iw[146]
port 131 nsew signal tristate
flabel metal4 s 166030 0 166090 200 0 FreeSans 480 90 0 0 um_iw[147]
port 132 nsew signal tristate
flabel metal4 s 165294 0 165354 200 0 FreeSans 480 90 0 0 um_iw[148]
port 133 nsew signal tristate
flabel metal4 s 164558 0 164618 200 0 FreeSans 480 90 0 0 um_iw[149]
port 134 nsew signal tristate
flabel metal4 s 21406 0 21466 200 0 FreeSans 480 90 0 0 um_iw[14]
port 135 nsew signal tristate
flabel metal4 s 163822 0 163882 200 0 FreeSans 480 90 0 0 um_iw[150]
port 136 nsew signal tristate
flabel metal4 s 163086 0 163146 200 0 FreeSans 480 90 0 0 um_iw[151]
port 137 nsew signal tristate
flabel metal4 s 162350 0 162410 200 0 FreeSans 480 90 0 0 um_iw[152]
port 138 nsew signal tristate
flabel metal4 s 161614 0 161674 200 0 FreeSans 480 90 0 0 um_iw[153]
port 139 nsew signal tristate
flabel metal4 s 160878 0 160938 200 0 FreeSans 480 90 0 0 um_iw[154]
port 140 nsew signal tristate
flabel metal4 s 160142 0 160202 200 0 FreeSans 480 90 0 0 um_iw[155]
port 141 nsew signal tristate
flabel metal4 s 159406 0 159466 200 0 FreeSans 480 90 0 0 um_iw[156]
port 142 nsew signal tristate
flabel metal4 s 158670 0 158730 200 0 FreeSans 480 90 0 0 um_iw[157]
port 143 nsew signal tristate
flabel metal4 s 157934 0 157994 200 0 FreeSans 480 90 0 0 um_iw[158]
port 144 nsew signal tristate
flabel metal4 s 157198 0 157258 200 0 FreeSans 480 90 0 0 um_iw[159]
port 145 nsew signal tristate
flabel metal4 s 20670 0 20730 200 0 FreeSans 480 90 0 0 um_iw[15]
port 146 nsew signal tristate
flabel metal4 s 156462 0 156522 200 0 FreeSans 480 90 0 0 um_iw[160]
port 147 nsew signal tristate
flabel metal4 s 155726 0 155786 200 0 FreeSans 480 90 0 0 um_iw[161]
port 148 nsew signal tristate
flabel metal4 s 168238 10680 168298 10880 0 FreeSans 480 90 0 0 um_iw[162]
port 149 nsew signal tristate
flabel metal4 s 167502 10680 167562 10880 0 FreeSans 480 90 0 0 um_iw[163]
port 150 nsew signal tristate
flabel metal4 s 166766 10680 166826 10880 0 FreeSans 480 90 0 0 um_iw[164]
port 151 nsew signal tristate
flabel metal4 s 166030 10680 166090 10880 0 FreeSans 480 90 0 0 um_iw[165]
port 152 nsew signal tristate
flabel metal4 s 165294 10680 165354 10880 0 FreeSans 480 90 0 0 um_iw[166]
port 153 nsew signal tristate
flabel metal4 s 164558 10680 164618 10880 0 FreeSans 480 90 0 0 um_iw[167]
port 154 nsew signal tristate
flabel metal4 s 163822 10680 163882 10880 0 FreeSans 480 90 0 0 um_iw[168]
port 155 nsew signal tristate
flabel metal4 s 163086 10680 163146 10880 0 FreeSans 480 90 0 0 um_iw[169]
port 156 nsew signal tristate
flabel metal4 s 19934 0 19994 200 0 FreeSans 480 90 0 0 um_iw[16]
port 157 nsew signal tristate
flabel metal4 s 162350 10680 162410 10880 0 FreeSans 480 90 0 0 um_iw[170]
port 158 nsew signal tristate
flabel metal4 s 161614 10680 161674 10880 0 FreeSans 480 90 0 0 um_iw[171]
port 159 nsew signal tristate
flabel metal4 s 160878 10680 160938 10880 0 FreeSans 480 90 0 0 um_iw[172]
port 160 nsew signal tristate
flabel metal4 s 160142 10680 160202 10880 0 FreeSans 480 90 0 0 um_iw[173]
port 161 nsew signal tristate
flabel metal4 s 159406 10680 159466 10880 0 FreeSans 480 90 0 0 um_iw[174]
port 162 nsew signal tristate
flabel metal4 s 158670 10680 158730 10880 0 FreeSans 480 90 0 0 um_iw[175]
port 163 nsew signal tristate
flabel metal4 s 157934 10680 157994 10880 0 FreeSans 480 90 0 0 um_iw[176]
port 164 nsew signal tristate
flabel metal4 s 157198 10680 157258 10880 0 FreeSans 480 90 0 0 um_iw[177]
port 165 nsew signal tristate
flabel metal4 s 156462 10680 156522 10880 0 FreeSans 480 90 0 0 um_iw[178]
port 166 nsew signal tristate
flabel metal4 s 155726 10680 155786 10880 0 FreeSans 480 90 0 0 um_iw[179]
port 167 nsew signal tristate
flabel metal4 s 19198 0 19258 200 0 FreeSans 480 90 0 0 um_iw[17]
port 168 nsew signal tristate
flabel metal4 s 202370 0 202430 200 0 FreeSans 480 90 0 0 um_iw[180]
port 169 nsew signal tristate
flabel metal4 s 201634 0 201694 200 0 FreeSans 480 90 0 0 um_iw[181]
port 170 nsew signal tristate
flabel metal4 s 200898 0 200958 200 0 FreeSans 480 90 0 0 um_iw[182]
port 171 nsew signal tristate
flabel metal4 s 200162 0 200222 200 0 FreeSans 480 90 0 0 um_iw[183]
port 172 nsew signal tristate
flabel metal4 s 199426 0 199486 200 0 FreeSans 480 90 0 0 um_iw[184]
port 173 nsew signal tristate
flabel metal4 s 198690 0 198750 200 0 FreeSans 480 90 0 0 um_iw[185]
port 174 nsew signal tristate
flabel metal4 s 197954 0 198014 200 0 FreeSans 480 90 0 0 um_iw[186]
port 175 nsew signal tristate
flabel metal4 s 197218 0 197278 200 0 FreeSans 480 90 0 0 um_iw[187]
port 176 nsew signal tristate
flabel metal4 s 196482 0 196542 200 0 FreeSans 480 90 0 0 um_iw[188]
port 177 nsew signal tristate
flabel metal4 s 195746 0 195806 200 0 FreeSans 480 90 0 0 um_iw[189]
port 178 nsew signal tristate
flabel metal4 s 31710 10680 31770 10880 0 FreeSans 480 90 0 0 um_iw[18]
port 179 nsew signal tristate
flabel metal4 s 195010 0 195070 200 0 FreeSans 480 90 0 0 um_iw[190]
port 180 nsew signal tristate
flabel metal4 s 194274 0 194334 200 0 FreeSans 480 90 0 0 um_iw[191]
port 181 nsew signal tristate
flabel metal4 s 193538 0 193598 200 0 FreeSans 480 90 0 0 um_iw[192]
port 182 nsew signal tristate
flabel metal4 s 192802 0 192862 200 0 FreeSans 480 90 0 0 um_iw[193]
port 183 nsew signal tristate
flabel metal4 s 192066 0 192126 200 0 FreeSans 480 90 0 0 um_iw[194]
port 184 nsew signal tristate
flabel metal4 s 191330 0 191390 200 0 FreeSans 480 90 0 0 um_iw[195]
port 185 nsew signal tristate
flabel metal4 s 190594 0 190654 200 0 FreeSans 480 90 0 0 um_iw[196]
port 186 nsew signal tristate
flabel metal4 s 189858 0 189918 200 0 FreeSans 480 90 0 0 um_iw[197]
port 187 nsew signal tristate
flabel metal4 s 202370 10680 202430 10880 0 FreeSans 480 90 0 0 um_iw[198]
port 188 nsew signal tristate
flabel metal4 s 201634 10680 201694 10880 0 FreeSans 480 90 0 0 um_iw[199]
port 189 nsew signal tristate
flabel metal4 s 30974 10680 31034 10880 0 FreeSans 480 90 0 0 um_iw[19]
port 190 nsew signal tristate
flabel metal4 s 30974 0 31034 200 0 FreeSans 480 90 0 0 um_iw[1]
port 191 nsew signal tristate
flabel metal4 s 200898 10680 200958 10880 0 FreeSans 480 90 0 0 um_iw[200]
port 192 nsew signal tristate
flabel metal4 s 200162 10680 200222 10880 0 FreeSans 480 90 0 0 um_iw[201]
port 193 nsew signal tristate
flabel metal4 s 199426 10680 199486 10880 0 FreeSans 480 90 0 0 um_iw[202]
port 194 nsew signal tristate
flabel metal4 s 198690 10680 198750 10880 0 FreeSans 480 90 0 0 um_iw[203]
port 195 nsew signal tristate
flabel metal4 s 197954 10680 198014 10880 0 FreeSans 480 90 0 0 um_iw[204]
port 196 nsew signal tristate
flabel metal4 s 197218 10680 197278 10880 0 FreeSans 480 90 0 0 um_iw[205]
port 197 nsew signal tristate
flabel metal4 s 196482 10680 196542 10880 0 FreeSans 480 90 0 0 um_iw[206]
port 198 nsew signal tristate
flabel metal4 s 195746 10680 195806 10880 0 FreeSans 480 90 0 0 um_iw[207]
port 199 nsew signal tristate
flabel metal4 s 195010 10680 195070 10880 0 FreeSans 480 90 0 0 um_iw[208]
port 200 nsew signal tristate
flabel metal4 s 194274 10680 194334 10880 0 FreeSans 480 90 0 0 um_iw[209]
port 201 nsew signal tristate
flabel metal4 s 30238 10680 30298 10880 0 FreeSans 480 90 0 0 um_iw[20]
port 202 nsew signal tristate
flabel metal4 s 193538 10680 193598 10880 0 FreeSans 480 90 0 0 um_iw[210]
port 203 nsew signal tristate
flabel metal4 s 192802 10680 192862 10880 0 FreeSans 480 90 0 0 um_iw[211]
port 204 nsew signal tristate
flabel metal4 s 192066 10680 192126 10880 0 FreeSans 480 90 0 0 um_iw[212]
port 205 nsew signal tristate
flabel metal4 s 191330 10680 191390 10880 0 FreeSans 480 90 0 0 um_iw[213]
port 206 nsew signal tristate
flabel metal4 s 190594 10680 190654 10880 0 FreeSans 480 90 0 0 um_iw[214]
port 207 nsew signal tristate
flabel metal4 s 189858 10680 189918 10880 0 FreeSans 480 90 0 0 um_iw[215]
port 208 nsew signal tristate
flabel metal4 s 236502 0 236562 200 0 FreeSans 480 90 0 0 um_iw[216]
port 209 nsew signal tristate
flabel metal4 s 235766 0 235826 200 0 FreeSans 480 90 0 0 um_iw[217]
port 210 nsew signal tristate
flabel metal4 s 235030 0 235090 200 0 FreeSans 480 90 0 0 um_iw[218]
port 211 nsew signal tristate
flabel metal4 s 234294 0 234354 200 0 FreeSans 480 90 0 0 um_iw[219]
port 212 nsew signal tristate
flabel metal4 s 29502 10680 29562 10880 0 FreeSans 480 90 0 0 um_iw[21]
port 213 nsew signal tristate
flabel metal4 s 233558 0 233618 200 0 FreeSans 480 90 0 0 um_iw[220]
port 214 nsew signal tristate
flabel metal4 s 232822 0 232882 200 0 FreeSans 480 90 0 0 um_iw[221]
port 215 nsew signal tristate
flabel metal4 s 232086 0 232146 200 0 FreeSans 480 90 0 0 um_iw[222]
port 216 nsew signal tristate
flabel metal4 s 231350 0 231410 200 0 FreeSans 480 90 0 0 um_iw[223]
port 217 nsew signal tristate
flabel metal4 s 230614 0 230674 200 0 FreeSans 480 90 0 0 um_iw[224]
port 218 nsew signal tristate
flabel metal4 s 229878 0 229938 200 0 FreeSans 480 90 0 0 um_iw[225]
port 219 nsew signal tristate
flabel metal4 s 229142 0 229202 200 0 FreeSans 480 90 0 0 um_iw[226]
port 220 nsew signal tristate
flabel metal4 s 228406 0 228466 200 0 FreeSans 480 90 0 0 um_iw[227]
port 221 nsew signal tristate
flabel metal4 s 227670 0 227730 200 0 FreeSans 480 90 0 0 um_iw[228]
port 222 nsew signal tristate
flabel metal4 s 226934 0 226994 200 0 FreeSans 480 90 0 0 um_iw[229]
port 223 nsew signal tristate
flabel metal4 s 28766 10680 28826 10880 0 FreeSans 480 90 0 0 um_iw[22]
port 224 nsew signal tristate
flabel metal4 s 226198 0 226258 200 0 FreeSans 480 90 0 0 um_iw[230]
port 225 nsew signal tristate
flabel metal4 s 225462 0 225522 200 0 FreeSans 480 90 0 0 um_iw[231]
port 226 nsew signal tristate
flabel metal4 s 224726 0 224786 200 0 FreeSans 480 90 0 0 um_iw[232]
port 227 nsew signal tristate
flabel metal4 s 223990 0 224050 200 0 FreeSans 480 90 0 0 um_iw[233]
port 228 nsew signal tristate
flabel metal4 s 236502 10680 236562 10880 0 FreeSans 480 90 0 0 um_iw[234]
port 229 nsew signal tristate
flabel metal4 s 235766 10680 235826 10880 0 FreeSans 480 90 0 0 um_iw[235]
port 230 nsew signal tristate
flabel metal4 s 235030 10680 235090 10880 0 FreeSans 480 90 0 0 um_iw[236]
port 231 nsew signal tristate
flabel metal4 s 234294 10680 234354 10880 0 FreeSans 480 90 0 0 um_iw[237]
port 232 nsew signal tristate
flabel metal4 s 233558 10680 233618 10880 0 FreeSans 480 90 0 0 um_iw[238]
port 233 nsew signal tristate
flabel metal4 s 232822 10680 232882 10880 0 FreeSans 480 90 0 0 um_iw[239]
port 234 nsew signal tristate
flabel metal4 s 28030 10680 28090 10880 0 FreeSans 480 90 0 0 um_iw[23]
port 235 nsew signal tristate
flabel metal4 s 232086 10680 232146 10880 0 FreeSans 480 90 0 0 um_iw[240]
port 236 nsew signal tristate
flabel metal4 s 231350 10680 231410 10880 0 FreeSans 480 90 0 0 um_iw[241]
port 237 nsew signal tristate
flabel metal4 s 230614 10680 230674 10880 0 FreeSans 480 90 0 0 um_iw[242]
port 238 nsew signal tristate
flabel metal4 s 229878 10680 229938 10880 0 FreeSans 480 90 0 0 um_iw[243]
port 239 nsew signal tristate
flabel metal4 s 229142 10680 229202 10880 0 FreeSans 480 90 0 0 um_iw[244]
port 240 nsew signal tristate
flabel metal4 s 228406 10680 228466 10880 0 FreeSans 480 90 0 0 um_iw[245]
port 241 nsew signal tristate
flabel metal4 s 227670 10680 227730 10880 0 FreeSans 480 90 0 0 um_iw[246]
port 242 nsew signal tristate
flabel metal4 s 226934 10680 226994 10880 0 FreeSans 480 90 0 0 um_iw[247]
port 243 nsew signal tristate
flabel metal4 s 226198 10680 226258 10880 0 FreeSans 480 90 0 0 um_iw[248]
port 244 nsew signal tristate
flabel metal4 s 225462 10680 225522 10880 0 FreeSans 480 90 0 0 um_iw[249]
port 245 nsew signal tristate
flabel metal4 s 27294 10680 27354 10880 0 FreeSans 480 90 0 0 um_iw[24]
port 246 nsew signal tristate
flabel metal4 s 224726 10680 224786 10880 0 FreeSans 480 90 0 0 um_iw[250]
port 247 nsew signal tristate
flabel metal4 s 223990 10680 224050 10880 0 FreeSans 480 90 0 0 um_iw[251]
port 248 nsew signal tristate
flabel metal4 s 270634 0 270694 200 0 FreeSans 480 90 0 0 um_iw[252]
port 249 nsew signal tristate
flabel metal4 s 269898 0 269958 200 0 FreeSans 480 90 0 0 um_iw[253]
port 250 nsew signal tristate
flabel metal4 s 269162 0 269222 200 0 FreeSans 480 90 0 0 um_iw[254]
port 251 nsew signal tristate
flabel metal4 s 268426 0 268486 200 0 FreeSans 480 90 0 0 um_iw[255]
port 252 nsew signal tristate
flabel metal4 s 267690 0 267750 200 0 FreeSans 480 90 0 0 um_iw[256]
port 253 nsew signal tristate
flabel metal4 s 266954 0 267014 200 0 FreeSans 480 90 0 0 um_iw[257]
port 254 nsew signal tristate
flabel metal4 s 266218 0 266278 200 0 FreeSans 480 90 0 0 um_iw[258]
port 255 nsew signal tristate
flabel metal4 s 265482 0 265542 200 0 FreeSans 480 90 0 0 um_iw[259]
port 256 nsew signal tristate
flabel metal4 s 26558 10680 26618 10880 0 FreeSans 480 90 0 0 um_iw[25]
port 257 nsew signal tristate
flabel metal4 s 264746 0 264806 200 0 FreeSans 480 90 0 0 um_iw[260]
port 258 nsew signal tristate
flabel metal4 s 264010 0 264070 200 0 FreeSans 480 90 0 0 um_iw[261]
port 259 nsew signal tristate
flabel metal4 s 263274 0 263334 200 0 FreeSans 480 90 0 0 um_iw[262]
port 260 nsew signal tristate
flabel metal4 s 262538 0 262598 200 0 FreeSans 480 90 0 0 um_iw[263]
port 261 nsew signal tristate
flabel metal4 s 261802 0 261862 200 0 FreeSans 480 90 0 0 um_iw[264]
port 262 nsew signal tristate
flabel metal4 s 261066 0 261126 200 0 FreeSans 480 90 0 0 um_iw[265]
port 263 nsew signal tristate
flabel metal4 s 260330 0 260390 200 0 FreeSans 480 90 0 0 um_iw[266]
port 264 nsew signal tristate
flabel metal4 s 259594 0 259654 200 0 FreeSans 480 90 0 0 um_iw[267]
port 265 nsew signal tristate
flabel metal4 s 258858 0 258918 200 0 FreeSans 480 90 0 0 um_iw[268]
port 266 nsew signal tristate
flabel metal4 s 258122 0 258182 200 0 FreeSans 480 90 0 0 um_iw[269]
port 267 nsew signal tristate
flabel metal4 s 25822 10680 25882 10880 0 FreeSans 480 90 0 0 um_iw[26]
port 268 nsew signal tristate
flabel metal4 s 270634 10680 270694 10880 0 FreeSans 480 90 0 0 um_iw[270]
port 269 nsew signal tristate
flabel metal4 s 269898 10680 269958 10880 0 FreeSans 480 90 0 0 um_iw[271]
port 270 nsew signal tristate
flabel metal4 s 269162 10680 269222 10880 0 FreeSans 480 90 0 0 um_iw[272]
port 271 nsew signal tristate
flabel metal4 s 268426 10680 268486 10880 0 FreeSans 480 90 0 0 um_iw[273]
port 272 nsew signal tristate
flabel metal4 s 267690 10680 267750 10880 0 FreeSans 480 90 0 0 um_iw[274]
port 273 nsew signal tristate
flabel metal4 s 266954 10680 267014 10880 0 FreeSans 480 90 0 0 um_iw[275]
port 274 nsew signal tristate
flabel metal4 s 266218 10680 266278 10880 0 FreeSans 480 90 0 0 um_iw[276]
port 275 nsew signal tristate
flabel metal4 s 265482 10680 265542 10880 0 FreeSans 480 90 0 0 um_iw[277]
port 276 nsew signal tristate
flabel metal4 s 264746 10680 264806 10880 0 FreeSans 480 90 0 0 um_iw[278]
port 277 nsew signal tristate
flabel metal4 s 264010 10680 264070 10880 0 FreeSans 480 90 0 0 um_iw[279]
port 278 nsew signal tristate
flabel metal4 s 25086 10680 25146 10880 0 FreeSans 480 90 0 0 um_iw[27]
port 279 nsew signal tristate
flabel metal4 s 263274 10680 263334 10880 0 FreeSans 480 90 0 0 um_iw[280]
port 280 nsew signal tristate
flabel metal4 s 262538 10680 262598 10880 0 FreeSans 480 90 0 0 um_iw[281]
port 281 nsew signal tristate
flabel metal4 s 261802 10680 261862 10880 0 FreeSans 480 90 0 0 um_iw[282]
port 282 nsew signal tristate
flabel metal4 s 261066 10680 261126 10880 0 FreeSans 480 90 0 0 um_iw[283]
port 283 nsew signal tristate
flabel metal4 s 260330 10680 260390 10880 0 FreeSans 480 90 0 0 um_iw[284]
port 284 nsew signal tristate
flabel metal4 s 259594 10680 259654 10880 0 FreeSans 480 90 0 0 um_iw[285]
port 285 nsew signal tristate
flabel metal4 s 258858 10680 258918 10880 0 FreeSans 480 90 0 0 um_iw[286]
port 286 nsew signal tristate
flabel metal4 s 258122 10680 258182 10880 0 FreeSans 480 90 0 0 um_iw[287]
port 287 nsew signal tristate
flabel metal4 s 24350 10680 24410 10880 0 FreeSans 480 90 0 0 um_iw[28]
port 288 nsew signal tristate
flabel metal4 s 23614 10680 23674 10880 0 FreeSans 480 90 0 0 um_iw[29]
port 289 nsew signal tristate
flabel metal4 s 30238 0 30298 200 0 FreeSans 480 90 0 0 um_iw[2]
port 290 nsew signal tristate
flabel metal4 s 22878 10680 22938 10880 0 FreeSans 480 90 0 0 um_iw[30]
port 291 nsew signal tristate
flabel metal4 s 22142 10680 22202 10880 0 FreeSans 480 90 0 0 um_iw[31]
port 292 nsew signal tristate
flabel metal4 s 21406 10680 21466 10880 0 FreeSans 480 90 0 0 um_iw[32]
port 293 nsew signal tristate
flabel metal4 s 20670 10680 20730 10880 0 FreeSans 480 90 0 0 um_iw[33]
port 294 nsew signal tristate
flabel metal4 s 19934 10680 19994 10880 0 FreeSans 480 90 0 0 um_iw[34]
port 295 nsew signal tristate
flabel metal4 s 19198 10680 19258 10880 0 FreeSans 480 90 0 0 um_iw[35]
port 296 nsew signal tristate
flabel metal4 s 65842 0 65902 200 0 FreeSans 480 90 0 0 um_iw[36]
port 297 nsew signal tristate
flabel metal4 s 65106 0 65166 200 0 FreeSans 480 90 0 0 um_iw[37]
port 298 nsew signal tristate
flabel metal4 s 64370 0 64430 200 0 FreeSans 480 90 0 0 um_iw[38]
port 299 nsew signal tristate
flabel metal4 s 63634 0 63694 200 0 FreeSans 480 90 0 0 um_iw[39]
port 300 nsew signal tristate
flabel metal4 s 29502 0 29562 200 0 FreeSans 480 90 0 0 um_iw[3]
port 301 nsew signal tristate
flabel metal4 s 62898 0 62958 200 0 FreeSans 480 90 0 0 um_iw[40]
port 302 nsew signal tristate
flabel metal4 s 62162 0 62222 200 0 FreeSans 480 90 0 0 um_iw[41]
port 303 nsew signal tristate
flabel metal4 s 61426 0 61486 200 0 FreeSans 480 90 0 0 um_iw[42]
port 304 nsew signal tristate
flabel metal4 s 60690 0 60750 200 0 FreeSans 480 90 0 0 um_iw[43]
port 305 nsew signal tristate
flabel metal4 s 59954 0 60014 200 0 FreeSans 480 90 0 0 um_iw[44]
port 306 nsew signal tristate
flabel metal4 s 59218 0 59278 200 0 FreeSans 480 90 0 0 um_iw[45]
port 307 nsew signal tristate
flabel metal4 s 58482 0 58542 200 0 FreeSans 480 90 0 0 um_iw[46]
port 308 nsew signal tristate
flabel metal4 s 57746 0 57806 200 0 FreeSans 480 90 0 0 um_iw[47]
port 309 nsew signal tristate
flabel metal4 s 57010 0 57070 200 0 FreeSans 480 90 0 0 um_iw[48]
port 310 nsew signal tristate
flabel metal4 s 56274 0 56334 200 0 FreeSans 480 90 0 0 um_iw[49]
port 311 nsew signal tristate
flabel metal4 s 28766 0 28826 200 0 FreeSans 480 90 0 0 um_iw[4]
port 312 nsew signal tristate
flabel metal4 s 55538 0 55598 200 0 FreeSans 480 90 0 0 um_iw[50]
port 313 nsew signal tristate
flabel metal4 s 54802 0 54862 200 0 FreeSans 480 90 0 0 um_iw[51]
port 314 nsew signal tristate
flabel metal4 s 54066 0 54126 200 0 FreeSans 480 90 0 0 um_iw[52]
port 315 nsew signal tristate
flabel metal4 s 53330 0 53390 200 0 FreeSans 480 90 0 0 um_iw[53]
port 316 nsew signal tristate
flabel metal4 s 65842 10680 65902 10880 0 FreeSans 480 90 0 0 um_iw[54]
port 317 nsew signal tristate
flabel metal4 s 65106 10680 65166 10880 0 FreeSans 480 90 0 0 um_iw[55]
port 318 nsew signal tristate
flabel metal4 s 64370 10680 64430 10880 0 FreeSans 480 90 0 0 um_iw[56]
port 319 nsew signal tristate
flabel metal4 s 63634 10680 63694 10880 0 FreeSans 480 90 0 0 um_iw[57]
port 320 nsew signal tristate
flabel metal4 s 62898 10680 62958 10880 0 FreeSans 480 90 0 0 um_iw[58]
port 321 nsew signal tristate
flabel metal4 s 62162 10680 62222 10880 0 FreeSans 480 90 0 0 um_iw[59]
port 322 nsew signal tristate
flabel metal4 s 28030 0 28090 200 0 FreeSans 480 90 0 0 um_iw[5]
port 323 nsew signal tristate
flabel metal4 s 61426 10680 61486 10880 0 FreeSans 480 90 0 0 um_iw[60]
port 324 nsew signal tristate
flabel metal4 s 60690 10680 60750 10880 0 FreeSans 480 90 0 0 um_iw[61]
port 325 nsew signal tristate
flabel metal4 s 59954 10680 60014 10880 0 FreeSans 480 90 0 0 um_iw[62]
port 326 nsew signal tristate
flabel metal4 s 59218 10680 59278 10880 0 FreeSans 480 90 0 0 um_iw[63]
port 327 nsew signal tristate
flabel metal4 s 58482 10680 58542 10880 0 FreeSans 480 90 0 0 um_iw[64]
port 328 nsew signal tristate
flabel metal4 s 57746 10680 57806 10880 0 FreeSans 480 90 0 0 um_iw[65]
port 329 nsew signal tristate
flabel metal4 s 57010 10680 57070 10880 0 FreeSans 480 90 0 0 um_iw[66]
port 330 nsew signal tristate
flabel metal4 s 56274 10680 56334 10880 0 FreeSans 480 90 0 0 um_iw[67]
port 331 nsew signal tristate
flabel metal4 s 55538 10680 55598 10880 0 FreeSans 480 90 0 0 um_iw[68]
port 332 nsew signal tristate
flabel metal4 s 54802 10680 54862 10880 0 FreeSans 480 90 0 0 um_iw[69]
port 333 nsew signal tristate
flabel metal4 s 27294 0 27354 200 0 FreeSans 480 90 0 0 um_iw[6]
port 334 nsew signal tristate
flabel metal4 s 54066 10680 54126 10880 0 FreeSans 480 90 0 0 um_iw[70]
port 335 nsew signal tristate
flabel metal4 s 53330 10680 53390 10880 0 FreeSans 480 90 0 0 um_iw[71]
port 336 nsew signal tristate
flabel metal4 s 99974 0 100034 200 0 FreeSans 480 90 0 0 um_iw[72]
port 337 nsew signal tristate
flabel metal4 s 99238 0 99298 200 0 FreeSans 480 90 0 0 um_iw[73]
port 338 nsew signal tristate
flabel metal4 s 98502 0 98562 200 0 FreeSans 480 90 0 0 um_iw[74]
port 339 nsew signal tristate
flabel metal4 s 97766 0 97826 200 0 FreeSans 480 90 0 0 um_iw[75]
port 340 nsew signal tristate
flabel metal4 s 97030 0 97090 200 0 FreeSans 480 90 0 0 um_iw[76]
port 341 nsew signal tristate
flabel metal4 s 96294 0 96354 200 0 FreeSans 480 90 0 0 um_iw[77]
port 342 nsew signal tristate
flabel metal4 s 95558 0 95618 200 0 FreeSans 480 90 0 0 um_iw[78]
port 343 nsew signal tristate
flabel metal4 s 94822 0 94882 200 0 FreeSans 480 90 0 0 um_iw[79]
port 344 nsew signal tristate
flabel metal4 s 26558 0 26618 200 0 FreeSans 480 90 0 0 um_iw[7]
port 345 nsew signal tristate
flabel metal4 s 94086 0 94146 200 0 FreeSans 480 90 0 0 um_iw[80]
port 346 nsew signal tristate
flabel metal4 s 93350 0 93410 200 0 FreeSans 480 90 0 0 um_iw[81]
port 347 nsew signal tristate
flabel metal4 s 92614 0 92674 200 0 FreeSans 480 90 0 0 um_iw[82]
port 348 nsew signal tristate
flabel metal4 s 91878 0 91938 200 0 FreeSans 480 90 0 0 um_iw[83]
port 349 nsew signal tristate
flabel metal4 s 91142 0 91202 200 0 FreeSans 480 90 0 0 um_iw[84]
port 350 nsew signal tristate
flabel metal4 s 90406 0 90466 200 0 FreeSans 480 90 0 0 um_iw[85]
port 351 nsew signal tristate
flabel metal4 s 89670 0 89730 200 0 FreeSans 480 90 0 0 um_iw[86]
port 352 nsew signal tristate
flabel metal4 s 88934 0 88994 200 0 FreeSans 480 90 0 0 um_iw[87]
port 353 nsew signal tristate
flabel metal4 s 88198 0 88258 200 0 FreeSans 480 90 0 0 um_iw[88]
port 354 nsew signal tristate
flabel metal4 s 87462 0 87522 200 0 FreeSans 480 90 0 0 um_iw[89]
port 355 nsew signal tristate
flabel metal4 s 25822 0 25882 200 0 FreeSans 480 90 0 0 um_iw[8]
port 356 nsew signal tristate
flabel metal4 s 99974 10680 100034 10880 0 FreeSans 480 90 0 0 um_iw[90]
port 357 nsew signal tristate
flabel metal4 s 99238 10680 99298 10880 0 FreeSans 480 90 0 0 um_iw[91]
port 358 nsew signal tristate
flabel metal4 s 98502 10680 98562 10880 0 FreeSans 480 90 0 0 um_iw[92]
port 359 nsew signal tristate
flabel metal4 s 97766 10680 97826 10880 0 FreeSans 480 90 0 0 um_iw[93]
port 360 nsew signal tristate
flabel metal4 s 97030 10680 97090 10880 0 FreeSans 480 90 0 0 um_iw[94]
port 361 nsew signal tristate
flabel metal4 s 96294 10680 96354 10880 0 FreeSans 480 90 0 0 um_iw[95]
port 362 nsew signal tristate
flabel metal4 s 95558 10680 95618 10880 0 FreeSans 480 90 0 0 um_iw[96]
port 363 nsew signal tristate
flabel metal4 s 94822 10680 94882 10880 0 FreeSans 480 90 0 0 um_iw[97]
port 364 nsew signal tristate
flabel metal4 s 94086 10680 94146 10880 0 FreeSans 480 90 0 0 um_iw[98]
port 365 nsew signal tristate
flabel metal4 s 93350 10680 93410 10880 0 FreeSans 480 90 0 0 um_iw[99]
port 366 nsew signal tristate
flabel metal4 s 25086 0 25146 200 0 FreeSans 480 90 0 0 um_iw[9]
port 367 nsew signal tristate
flabel metal4 s 798 0 858 200 0 FreeSans 480 90 0 0 um_k_zero[0]
port 368 nsew signal tristate
flabel metal4 s 171458 0 171518 200 0 FreeSans 480 90 0 0 um_k_zero[10]
port 369 nsew signal tristate
flabel metal4 s 171458 10680 171518 10880 0 FreeSans 480 90 0 0 um_k_zero[11]
port 370 nsew signal tristate
flabel metal4 s 205590 0 205650 200 0 FreeSans 480 90 0 0 um_k_zero[12]
port 371 nsew signal tristate
flabel metal4 s 205590 10680 205650 10880 0 FreeSans 480 90 0 0 um_k_zero[13]
port 372 nsew signal tristate
flabel metal4 s 239722 0 239782 200 0 FreeSans 480 90 0 0 um_k_zero[14]
port 373 nsew signal tristate
flabel metal4 s 239722 10680 239782 10880 0 FreeSans 480 90 0 0 um_k_zero[15]
port 374 nsew signal tristate
flabel metal4 s 798 10680 858 10880 0 FreeSans 480 90 0 0 um_k_zero[1]
port 375 nsew signal tristate
flabel metal4 s 34930 0 34990 200 0 FreeSans 480 90 0 0 um_k_zero[2]
port 376 nsew signal tristate
flabel metal4 s 34930 10680 34990 10880 0 FreeSans 480 90 0 0 um_k_zero[3]
port 377 nsew signal tristate
flabel metal4 s 69062 0 69122 200 0 FreeSans 480 90 0 0 um_k_zero[4]
port 378 nsew signal tristate
flabel metal4 s 69062 10680 69122 10880 0 FreeSans 480 90 0 0 um_k_zero[5]
port 379 nsew signal tristate
flabel metal4 s 103194 0 103254 200 0 FreeSans 480 90 0 0 um_k_zero[6]
port 380 nsew signal tristate
flabel metal4 s 103194 10680 103254 10880 0 FreeSans 480 90 0 0 um_k_zero[7]
port 381 nsew signal tristate
flabel metal4 s 137326 0 137386 200 0 FreeSans 480 90 0 0 um_k_zero[8]
port 382 nsew signal tristate
flabel metal4 s 137326 10680 137386 10880 0 FreeSans 480 90 0 0 um_k_zero[9]
port 383 nsew signal tristate
flabel metal4 s 18462 0 18522 200 0 FreeSans 480 90 0 0 um_ow[0]
port 384 nsew signal input
flabel metal4 s 83782 0 83842 200 0 FreeSans 480 90 0 0 um_ow[100]
port 385 nsew signal input
flabel metal4 s 83046 0 83106 200 0 FreeSans 480 90 0 0 um_ow[101]
port 386 nsew signal input
flabel metal4 s 82310 0 82370 200 0 FreeSans 480 90 0 0 um_ow[102]
port 387 nsew signal input
flabel metal4 s 81574 0 81634 200 0 FreeSans 480 90 0 0 um_ow[103]
port 388 nsew signal input
flabel metal4 s 80838 0 80898 200 0 FreeSans 480 90 0 0 um_ow[104]
port 389 nsew signal input
flabel metal4 s 80102 0 80162 200 0 FreeSans 480 90 0 0 um_ow[105]
port 390 nsew signal input
flabel metal4 s 79366 0 79426 200 0 FreeSans 480 90 0 0 um_ow[106]
port 391 nsew signal input
flabel metal4 s 78630 0 78690 200 0 FreeSans 480 90 0 0 um_ow[107]
port 392 nsew signal input
flabel metal4 s 77894 0 77954 200 0 FreeSans 480 90 0 0 um_ow[108]
port 393 nsew signal input
flabel metal4 s 77158 0 77218 200 0 FreeSans 480 90 0 0 um_ow[109]
port 394 nsew signal input
flabel metal4 s 11102 0 11162 200 0 FreeSans 480 90 0 0 um_ow[10]
port 395 nsew signal input
flabel metal4 s 76422 0 76482 200 0 FreeSans 480 90 0 0 um_ow[110]
port 396 nsew signal input
flabel metal4 s 75686 0 75746 200 0 FreeSans 480 90 0 0 um_ow[111]
port 397 nsew signal input
flabel metal4 s 74950 0 75010 200 0 FreeSans 480 90 0 0 um_ow[112]
port 398 nsew signal input
flabel metal4 s 74214 0 74274 200 0 FreeSans 480 90 0 0 um_ow[113]
port 399 nsew signal input
flabel metal4 s 73478 0 73538 200 0 FreeSans 480 90 0 0 um_ow[114]
port 400 nsew signal input
flabel metal4 s 72742 0 72802 200 0 FreeSans 480 90 0 0 um_ow[115]
port 401 nsew signal input
flabel metal4 s 72006 0 72066 200 0 FreeSans 480 90 0 0 um_ow[116]
port 402 nsew signal input
flabel metal4 s 71270 0 71330 200 0 FreeSans 480 90 0 0 um_ow[117]
port 403 nsew signal input
flabel metal4 s 70534 0 70594 200 0 FreeSans 480 90 0 0 um_ow[118]
port 404 nsew signal input
flabel metal4 s 69798 0 69858 200 0 FreeSans 480 90 0 0 um_ow[119]
port 405 nsew signal input
flabel metal4 s 10366 0 10426 200 0 FreeSans 480 90 0 0 um_ow[11]
port 406 nsew signal input
flabel metal4 s 86726 10680 86786 10880 0 FreeSans 480 90 0 0 um_ow[120]
port 407 nsew signal input
flabel metal4 s 85990 10680 86050 10880 0 FreeSans 480 90 0 0 um_ow[121]
port 408 nsew signal input
flabel metal4 s 85254 10680 85314 10880 0 FreeSans 480 90 0 0 um_ow[122]
port 409 nsew signal input
flabel metal4 s 84518 10680 84578 10880 0 FreeSans 480 90 0 0 um_ow[123]
port 410 nsew signal input
flabel metal4 s 83782 10680 83842 10880 0 FreeSans 480 90 0 0 um_ow[124]
port 411 nsew signal input
flabel metal4 s 83046 10680 83106 10880 0 FreeSans 480 90 0 0 um_ow[125]
port 412 nsew signal input
flabel metal4 s 82310 10680 82370 10880 0 FreeSans 480 90 0 0 um_ow[126]
port 413 nsew signal input
flabel metal4 s 81574 10680 81634 10880 0 FreeSans 480 90 0 0 um_ow[127]
port 414 nsew signal input
flabel metal4 s 80838 10680 80898 10880 0 FreeSans 480 90 0 0 um_ow[128]
port 415 nsew signal input
flabel metal4 s 80102 10680 80162 10880 0 FreeSans 480 90 0 0 um_ow[129]
port 416 nsew signal input
flabel metal4 s 9630 0 9690 200 0 FreeSans 480 90 0 0 um_ow[12]
port 417 nsew signal input
flabel metal4 s 79366 10680 79426 10880 0 FreeSans 480 90 0 0 um_ow[130]
port 418 nsew signal input
flabel metal4 s 78630 10680 78690 10880 0 FreeSans 480 90 0 0 um_ow[131]
port 419 nsew signal input
flabel metal4 s 77894 10680 77954 10880 0 FreeSans 480 90 0 0 um_ow[132]
port 420 nsew signal input
flabel metal4 s 77158 10680 77218 10880 0 FreeSans 480 90 0 0 um_ow[133]
port 421 nsew signal input
flabel metal4 s 76422 10680 76482 10880 0 FreeSans 480 90 0 0 um_ow[134]
port 422 nsew signal input
flabel metal4 s 75686 10680 75746 10880 0 FreeSans 480 90 0 0 um_ow[135]
port 423 nsew signal input
flabel metal4 s 74950 10680 75010 10880 0 FreeSans 480 90 0 0 um_ow[136]
port 424 nsew signal input
flabel metal4 s 74214 10680 74274 10880 0 FreeSans 480 90 0 0 um_ow[137]
port 425 nsew signal input
flabel metal4 s 73478 10680 73538 10880 0 FreeSans 480 90 0 0 um_ow[138]
port 426 nsew signal input
flabel metal4 s 72742 10680 72802 10880 0 FreeSans 480 90 0 0 um_ow[139]
port 427 nsew signal input
flabel metal4 s 8894 0 8954 200 0 FreeSans 480 90 0 0 um_ow[13]
port 428 nsew signal input
flabel metal4 s 72006 10680 72066 10880 0 FreeSans 480 90 0 0 um_ow[140]
port 429 nsew signal input
flabel metal4 s 71270 10680 71330 10880 0 FreeSans 480 90 0 0 um_ow[141]
port 430 nsew signal input
flabel metal4 s 70534 10680 70594 10880 0 FreeSans 480 90 0 0 um_ow[142]
port 431 nsew signal input
flabel metal4 s 69798 10680 69858 10880 0 FreeSans 480 90 0 0 um_ow[143]
port 432 nsew signal input
flabel metal4 s 120858 0 120918 200 0 FreeSans 480 90 0 0 um_ow[144]
port 433 nsew signal input
flabel metal4 s 120122 0 120182 200 0 FreeSans 480 90 0 0 um_ow[145]
port 434 nsew signal input
flabel metal4 s 119386 0 119446 200 0 FreeSans 480 90 0 0 um_ow[146]
port 435 nsew signal input
flabel metal4 s 118650 0 118710 200 0 FreeSans 480 90 0 0 um_ow[147]
port 436 nsew signal input
flabel metal4 s 117914 0 117974 200 0 FreeSans 480 90 0 0 um_ow[148]
port 437 nsew signal input
flabel metal4 s 117178 0 117238 200 0 FreeSans 480 90 0 0 um_ow[149]
port 438 nsew signal input
flabel metal4 s 8158 0 8218 200 0 FreeSans 480 90 0 0 um_ow[14]
port 439 nsew signal input
flabel metal4 s 116442 0 116502 200 0 FreeSans 480 90 0 0 um_ow[150]
port 440 nsew signal input
flabel metal4 s 115706 0 115766 200 0 FreeSans 480 90 0 0 um_ow[151]
port 441 nsew signal input
flabel metal4 s 114970 0 115030 200 0 FreeSans 480 90 0 0 um_ow[152]
port 442 nsew signal input
flabel metal4 s 114234 0 114294 200 0 FreeSans 480 90 0 0 um_ow[153]
port 443 nsew signal input
flabel metal4 s 113498 0 113558 200 0 FreeSans 480 90 0 0 um_ow[154]
port 444 nsew signal input
flabel metal4 s 112762 0 112822 200 0 FreeSans 480 90 0 0 um_ow[155]
port 445 nsew signal input
flabel metal4 s 112026 0 112086 200 0 FreeSans 480 90 0 0 um_ow[156]
port 446 nsew signal input
flabel metal4 s 111290 0 111350 200 0 FreeSans 480 90 0 0 um_ow[157]
port 447 nsew signal input
flabel metal4 s 110554 0 110614 200 0 FreeSans 480 90 0 0 um_ow[158]
port 448 nsew signal input
flabel metal4 s 109818 0 109878 200 0 FreeSans 480 90 0 0 um_ow[159]
port 449 nsew signal input
flabel metal4 s 7422 0 7482 200 0 FreeSans 480 90 0 0 um_ow[15]
port 450 nsew signal input
flabel metal4 s 109082 0 109142 200 0 FreeSans 480 90 0 0 um_ow[160]
port 451 nsew signal input
flabel metal4 s 108346 0 108406 200 0 FreeSans 480 90 0 0 um_ow[161]
port 452 nsew signal input
flabel metal4 s 107610 0 107670 200 0 FreeSans 480 90 0 0 um_ow[162]
port 453 nsew signal input
flabel metal4 s 106874 0 106934 200 0 FreeSans 480 90 0 0 um_ow[163]
port 454 nsew signal input
flabel metal4 s 106138 0 106198 200 0 FreeSans 480 90 0 0 um_ow[164]
port 455 nsew signal input
flabel metal4 s 105402 0 105462 200 0 FreeSans 480 90 0 0 um_ow[165]
port 456 nsew signal input
flabel metal4 s 104666 0 104726 200 0 FreeSans 480 90 0 0 um_ow[166]
port 457 nsew signal input
flabel metal4 s 103930 0 103990 200 0 FreeSans 480 90 0 0 um_ow[167]
port 458 nsew signal input
flabel metal4 s 120858 10680 120918 10880 0 FreeSans 480 90 0 0 um_ow[168]
port 459 nsew signal input
flabel metal4 s 120122 10680 120182 10880 0 FreeSans 480 90 0 0 um_ow[169]
port 460 nsew signal input
flabel metal4 s 6686 0 6746 200 0 FreeSans 480 90 0 0 um_ow[16]
port 461 nsew signal input
flabel metal4 s 119386 10680 119446 10880 0 FreeSans 480 90 0 0 um_ow[170]
port 462 nsew signal input
flabel metal4 s 118650 10680 118710 10880 0 FreeSans 480 90 0 0 um_ow[171]
port 463 nsew signal input
flabel metal4 s 117914 10680 117974 10880 0 FreeSans 480 90 0 0 um_ow[172]
port 464 nsew signal input
flabel metal4 s 117178 10680 117238 10880 0 FreeSans 480 90 0 0 um_ow[173]
port 465 nsew signal input
flabel metal4 s 116442 10680 116502 10880 0 FreeSans 480 90 0 0 um_ow[174]
port 466 nsew signal input
flabel metal4 s 115706 10680 115766 10880 0 FreeSans 480 90 0 0 um_ow[175]
port 467 nsew signal input
flabel metal4 s 114970 10680 115030 10880 0 FreeSans 480 90 0 0 um_ow[176]
port 468 nsew signal input
flabel metal4 s 114234 10680 114294 10880 0 FreeSans 480 90 0 0 um_ow[177]
port 469 nsew signal input
flabel metal4 s 113498 10680 113558 10880 0 FreeSans 480 90 0 0 um_ow[178]
port 470 nsew signal input
flabel metal4 s 112762 10680 112822 10880 0 FreeSans 480 90 0 0 um_ow[179]
port 471 nsew signal input
flabel metal4 s 5950 0 6010 200 0 FreeSans 480 90 0 0 um_ow[17]
port 472 nsew signal input
flabel metal4 s 112026 10680 112086 10880 0 FreeSans 480 90 0 0 um_ow[180]
port 473 nsew signal input
flabel metal4 s 111290 10680 111350 10880 0 FreeSans 480 90 0 0 um_ow[181]
port 474 nsew signal input
flabel metal4 s 110554 10680 110614 10880 0 FreeSans 480 90 0 0 um_ow[182]
port 475 nsew signal input
flabel metal4 s 109818 10680 109878 10880 0 FreeSans 480 90 0 0 um_ow[183]
port 476 nsew signal input
flabel metal4 s 109082 10680 109142 10880 0 FreeSans 480 90 0 0 um_ow[184]
port 477 nsew signal input
flabel metal4 s 108346 10680 108406 10880 0 FreeSans 480 90 0 0 um_ow[185]
port 478 nsew signal input
flabel metal4 s 107610 10680 107670 10880 0 FreeSans 480 90 0 0 um_ow[186]
port 479 nsew signal input
flabel metal4 s 106874 10680 106934 10880 0 FreeSans 480 90 0 0 um_ow[187]
port 480 nsew signal input
flabel metal4 s 106138 10680 106198 10880 0 FreeSans 480 90 0 0 um_ow[188]
port 481 nsew signal input
flabel metal4 s 105402 10680 105462 10880 0 FreeSans 480 90 0 0 um_ow[189]
port 482 nsew signal input
flabel metal4 s 5214 0 5274 200 0 FreeSans 480 90 0 0 um_ow[18]
port 483 nsew signal input
flabel metal4 s 104666 10680 104726 10880 0 FreeSans 480 90 0 0 um_ow[190]
port 484 nsew signal input
flabel metal4 s 103930 10680 103990 10880 0 FreeSans 480 90 0 0 um_ow[191]
port 485 nsew signal input
flabel metal4 s 154990 0 155050 200 0 FreeSans 480 90 0 0 um_ow[192]
port 486 nsew signal input
flabel metal4 s 154254 0 154314 200 0 FreeSans 480 90 0 0 um_ow[193]
port 487 nsew signal input
flabel metal4 s 153518 0 153578 200 0 FreeSans 480 90 0 0 um_ow[194]
port 488 nsew signal input
flabel metal4 s 152782 0 152842 200 0 FreeSans 480 90 0 0 um_ow[195]
port 489 nsew signal input
flabel metal4 s 152046 0 152106 200 0 FreeSans 480 90 0 0 um_ow[196]
port 490 nsew signal input
flabel metal4 s 151310 0 151370 200 0 FreeSans 480 90 0 0 um_ow[197]
port 491 nsew signal input
flabel metal4 s 150574 0 150634 200 0 FreeSans 480 90 0 0 um_ow[198]
port 492 nsew signal input
flabel metal4 s 149838 0 149898 200 0 FreeSans 480 90 0 0 um_ow[199]
port 493 nsew signal input
flabel metal4 s 4478 0 4538 200 0 FreeSans 480 90 0 0 um_ow[19]
port 494 nsew signal input
flabel metal4 s 17726 0 17786 200 0 FreeSans 480 90 0 0 um_ow[1]
port 495 nsew signal input
flabel metal4 s 149102 0 149162 200 0 FreeSans 480 90 0 0 um_ow[200]
port 496 nsew signal input
flabel metal4 s 148366 0 148426 200 0 FreeSans 480 90 0 0 um_ow[201]
port 497 nsew signal input
flabel metal4 s 147630 0 147690 200 0 FreeSans 480 90 0 0 um_ow[202]
port 498 nsew signal input
flabel metal4 s 146894 0 146954 200 0 FreeSans 480 90 0 0 um_ow[203]
port 499 nsew signal input
flabel metal4 s 146158 0 146218 200 0 FreeSans 480 90 0 0 um_ow[204]
port 500 nsew signal input
flabel metal4 s 145422 0 145482 200 0 FreeSans 480 90 0 0 um_ow[205]
port 501 nsew signal input
flabel metal4 s 144686 0 144746 200 0 FreeSans 480 90 0 0 um_ow[206]
port 502 nsew signal input
flabel metal4 s 143950 0 144010 200 0 FreeSans 480 90 0 0 um_ow[207]
port 503 nsew signal input
flabel metal4 s 143214 0 143274 200 0 FreeSans 480 90 0 0 um_ow[208]
port 504 nsew signal input
flabel metal4 s 142478 0 142538 200 0 FreeSans 480 90 0 0 um_ow[209]
port 505 nsew signal input
flabel metal4 s 3742 0 3802 200 0 FreeSans 480 90 0 0 um_ow[20]
port 506 nsew signal input
flabel metal4 s 141742 0 141802 200 0 FreeSans 480 90 0 0 um_ow[210]
port 507 nsew signal input
flabel metal4 s 141006 0 141066 200 0 FreeSans 480 90 0 0 um_ow[211]
port 508 nsew signal input
flabel metal4 s 140270 0 140330 200 0 FreeSans 480 90 0 0 um_ow[212]
port 509 nsew signal input
flabel metal4 s 139534 0 139594 200 0 FreeSans 480 90 0 0 um_ow[213]
port 510 nsew signal input
flabel metal4 s 138798 0 138858 200 0 FreeSans 480 90 0 0 um_ow[214]
port 511 nsew signal input
flabel metal4 s 138062 0 138122 200 0 FreeSans 480 90 0 0 um_ow[215]
port 512 nsew signal input
flabel metal4 s 154990 10680 155050 10880 0 FreeSans 480 90 0 0 um_ow[216]
port 513 nsew signal input
flabel metal4 s 154254 10680 154314 10880 0 FreeSans 480 90 0 0 um_ow[217]
port 514 nsew signal input
flabel metal4 s 153518 10680 153578 10880 0 FreeSans 480 90 0 0 um_ow[218]
port 515 nsew signal input
flabel metal4 s 152782 10680 152842 10880 0 FreeSans 480 90 0 0 um_ow[219]
port 516 nsew signal input
flabel metal4 s 3006 0 3066 200 0 FreeSans 480 90 0 0 um_ow[21]
port 517 nsew signal input
flabel metal4 s 152046 10680 152106 10880 0 FreeSans 480 90 0 0 um_ow[220]
port 518 nsew signal input
flabel metal4 s 151310 10680 151370 10880 0 FreeSans 480 90 0 0 um_ow[221]
port 519 nsew signal input
flabel metal4 s 150574 10680 150634 10880 0 FreeSans 480 90 0 0 um_ow[222]
port 520 nsew signal input
flabel metal4 s 149838 10680 149898 10880 0 FreeSans 480 90 0 0 um_ow[223]
port 521 nsew signal input
flabel metal4 s 149102 10680 149162 10880 0 FreeSans 480 90 0 0 um_ow[224]
port 522 nsew signal input
flabel metal4 s 148366 10680 148426 10880 0 FreeSans 480 90 0 0 um_ow[225]
port 523 nsew signal input
flabel metal4 s 147630 10680 147690 10880 0 FreeSans 480 90 0 0 um_ow[226]
port 524 nsew signal input
flabel metal4 s 146894 10680 146954 10880 0 FreeSans 480 90 0 0 um_ow[227]
port 525 nsew signal input
flabel metal4 s 146158 10680 146218 10880 0 FreeSans 480 90 0 0 um_ow[228]
port 526 nsew signal input
flabel metal4 s 145422 10680 145482 10880 0 FreeSans 480 90 0 0 um_ow[229]
port 527 nsew signal input
flabel metal4 s 2270 0 2330 200 0 FreeSans 480 90 0 0 um_ow[22]
port 528 nsew signal input
flabel metal4 s 144686 10680 144746 10880 0 FreeSans 480 90 0 0 um_ow[230]
port 529 nsew signal input
flabel metal4 s 143950 10680 144010 10880 0 FreeSans 480 90 0 0 um_ow[231]
port 530 nsew signal input
flabel metal4 s 143214 10680 143274 10880 0 FreeSans 480 90 0 0 um_ow[232]
port 531 nsew signal input
flabel metal4 s 142478 10680 142538 10880 0 FreeSans 480 90 0 0 um_ow[233]
port 532 nsew signal input
flabel metal4 s 141742 10680 141802 10880 0 FreeSans 480 90 0 0 um_ow[234]
port 533 nsew signal input
flabel metal4 s 141006 10680 141066 10880 0 FreeSans 480 90 0 0 um_ow[235]
port 534 nsew signal input
flabel metal4 s 140270 10680 140330 10880 0 FreeSans 480 90 0 0 um_ow[236]
port 535 nsew signal input
flabel metal4 s 139534 10680 139594 10880 0 FreeSans 480 90 0 0 um_ow[237]
port 536 nsew signal input
flabel metal4 s 138798 10680 138858 10880 0 FreeSans 480 90 0 0 um_ow[238]
port 537 nsew signal input
flabel metal4 s 138062 10680 138122 10880 0 FreeSans 480 90 0 0 um_ow[239]
port 538 nsew signal input
flabel metal4 s 1534 0 1594 200 0 FreeSans 480 90 0 0 um_ow[23]
port 539 nsew signal input
flabel metal4 s 189122 0 189182 200 0 FreeSans 480 90 0 0 um_ow[240]
port 540 nsew signal input
flabel metal4 s 188386 0 188446 200 0 FreeSans 480 90 0 0 um_ow[241]
port 541 nsew signal input
flabel metal4 s 187650 0 187710 200 0 FreeSans 480 90 0 0 um_ow[242]
port 542 nsew signal input
flabel metal4 s 186914 0 186974 200 0 FreeSans 480 90 0 0 um_ow[243]
port 543 nsew signal input
flabel metal4 s 186178 0 186238 200 0 FreeSans 480 90 0 0 um_ow[244]
port 544 nsew signal input
flabel metal4 s 185442 0 185502 200 0 FreeSans 480 90 0 0 um_ow[245]
port 545 nsew signal input
flabel metal4 s 184706 0 184766 200 0 FreeSans 480 90 0 0 um_ow[246]
port 546 nsew signal input
flabel metal4 s 183970 0 184030 200 0 FreeSans 480 90 0 0 um_ow[247]
port 547 nsew signal input
flabel metal4 s 183234 0 183294 200 0 FreeSans 480 90 0 0 um_ow[248]
port 548 nsew signal input
flabel metal4 s 182498 0 182558 200 0 FreeSans 480 90 0 0 um_ow[249]
port 549 nsew signal input
flabel metal4 s 18462 10680 18522 10880 0 FreeSans 480 90 0 0 um_ow[24]
port 550 nsew signal input
flabel metal4 s 181762 0 181822 200 0 FreeSans 480 90 0 0 um_ow[250]
port 551 nsew signal input
flabel metal4 s 181026 0 181086 200 0 FreeSans 480 90 0 0 um_ow[251]
port 552 nsew signal input
flabel metal4 s 180290 0 180350 200 0 FreeSans 480 90 0 0 um_ow[252]
port 553 nsew signal input
flabel metal4 s 179554 0 179614 200 0 FreeSans 480 90 0 0 um_ow[253]
port 554 nsew signal input
flabel metal4 s 178818 0 178878 200 0 FreeSans 480 90 0 0 um_ow[254]
port 555 nsew signal input
flabel metal4 s 178082 0 178142 200 0 FreeSans 480 90 0 0 um_ow[255]
port 556 nsew signal input
flabel metal4 s 177346 0 177406 200 0 FreeSans 480 90 0 0 um_ow[256]
port 557 nsew signal input
flabel metal4 s 176610 0 176670 200 0 FreeSans 480 90 0 0 um_ow[257]
port 558 nsew signal input
flabel metal4 s 175874 0 175934 200 0 FreeSans 480 90 0 0 um_ow[258]
port 559 nsew signal input
flabel metal4 s 175138 0 175198 200 0 FreeSans 480 90 0 0 um_ow[259]
port 560 nsew signal input
flabel metal4 s 17726 10680 17786 10880 0 FreeSans 480 90 0 0 um_ow[25]
port 561 nsew signal input
flabel metal4 s 174402 0 174462 200 0 FreeSans 480 90 0 0 um_ow[260]
port 562 nsew signal input
flabel metal4 s 173666 0 173726 200 0 FreeSans 480 90 0 0 um_ow[261]
port 563 nsew signal input
flabel metal4 s 172930 0 172990 200 0 FreeSans 480 90 0 0 um_ow[262]
port 564 nsew signal input
flabel metal4 s 172194 0 172254 200 0 FreeSans 480 90 0 0 um_ow[263]
port 565 nsew signal input
flabel metal4 s 189122 10680 189182 10880 0 FreeSans 480 90 0 0 um_ow[264]
port 566 nsew signal input
flabel metal4 s 188386 10680 188446 10880 0 FreeSans 480 90 0 0 um_ow[265]
port 567 nsew signal input
flabel metal4 s 187650 10680 187710 10880 0 FreeSans 480 90 0 0 um_ow[266]
port 568 nsew signal input
flabel metal4 s 186914 10680 186974 10880 0 FreeSans 480 90 0 0 um_ow[267]
port 569 nsew signal input
flabel metal4 s 186178 10680 186238 10880 0 FreeSans 480 90 0 0 um_ow[268]
port 570 nsew signal input
flabel metal4 s 185442 10680 185502 10880 0 FreeSans 480 90 0 0 um_ow[269]
port 571 nsew signal input
flabel metal4 s 16990 10680 17050 10880 0 FreeSans 480 90 0 0 um_ow[26]
port 572 nsew signal input
flabel metal4 s 184706 10680 184766 10880 0 FreeSans 480 90 0 0 um_ow[270]
port 573 nsew signal input
flabel metal4 s 183970 10680 184030 10880 0 FreeSans 480 90 0 0 um_ow[271]
port 574 nsew signal input
flabel metal4 s 183234 10680 183294 10880 0 FreeSans 480 90 0 0 um_ow[272]
port 575 nsew signal input
flabel metal4 s 182498 10680 182558 10880 0 FreeSans 480 90 0 0 um_ow[273]
port 576 nsew signal input
flabel metal4 s 181762 10680 181822 10880 0 FreeSans 480 90 0 0 um_ow[274]
port 577 nsew signal input
flabel metal4 s 181026 10680 181086 10880 0 FreeSans 480 90 0 0 um_ow[275]
port 578 nsew signal input
flabel metal4 s 180290 10680 180350 10880 0 FreeSans 480 90 0 0 um_ow[276]
port 579 nsew signal input
flabel metal4 s 179554 10680 179614 10880 0 FreeSans 480 90 0 0 um_ow[277]
port 580 nsew signal input
flabel metal4 s 178818 10680 178878 10880 0 FreeSans 480 90 0 0 um_ow[278]
port 581 nsew signal input
flabel metal4 s 178082 10680 178142 10880 0 FreeSans 480 90 0 0 um_ow[279]
port 582 nsew signal input
flabel metal4 s 16254 10680 16314 10880 0 FreeSans 480 90 0 0 um_ow[27]
port 583 nsew signal input
flabel metal4 s 177346 10680 177406 10880 0 FreeSans 480 90 0 0 um_ow[280]
port 584 nsew signal input
flabel metal4 s 176610 10680 176670 10880 0 FreeSans 480 90 0 0 um_ow[281]
port 585 nsew signal input
flabel metal4 s 175874 10680 175934 10880 0 FreeSans 480 90 0 0 um_ow[282]
port 586 nsew signal input
flabel metal4 s 175138 10680 175198 10880 0 FreeSans 480 90 0 0 um_ow[283]
port 587 nsew signal input
flabel metal4 s 174402 10680 174462 10880 0 FreeSans 480 90 0 0 um_ow[284]
port 588 nsew signal input
flabel metal4 s 173666 10680 173726 10880 0 FreeSans 480 90 0 0 um_ow[285]
port 589 nsew signal input
flabel metal4 s 172930 10680 172990 10880 0 FreeSans 480 90 0 0 um_ow[286]
port 590 nsew signal input
flabel metal4 s 172194 10680 172254 10880 0 FreeSans 480 90 0 0 um_ow[287]
port 591 nsew signal input
flabel metal4 s 223254 0 223314 200 0 FreeSans 480 90 0 0 um_ow[288]
port 592 nsew signal input
flabel metal4 s 222518 0 222578 200 0 FreeSans 480 90 0 0 um_ow[289]
port 593 nsew signal input
flabel metal4 s 15518 10680 15578 10880 0 FreeSans 480 90 0 0 um_ow[28]
port 594 nsew signal input
flabel metal4 s 221782 0 221842 200 0 FreeSans 480 90 0 0 um_ow[290]
port 595 nsew signal input
flabel metal4 s 221046 0 221106 200 0 FreeSans 480 90 0 0 um_ow[291]
port 596 nsew signal input
flabel metal4 s 220310 0 220370 200 0 FreeSans 480 90 0 0 um_ow[292]
port 597 nsew signal input
flabel metal4 s 219574 0 219634 200 0 FreeSans 480 90 0 0 um_ow[293]
port 598 nsew signal input
flabel metal4 s 218838 0 218898 200 0 FreeSans 480 90 0 0 um_ow[294]
port 599 nsew signal input
flabel metal4 s 218102 0 218162 200 0 FreeSans 480 90 0 0 um_ow[295]
port 600 nsew signal input
flabel metal4 s 217366 0 217426 200 0 FreeSans 480 90 0 0 um_ow[296]
port 601 nsew signal input
flabel metal4 s 216630 0 216690 200 0 FreeSans 480 90 0 0 um_ow[297]
port 602 nsew signal input
flabel metal4 s 215894 0 215954 200 0 FreeSans 480 90 0 0 um_ow[298]
port 603 nsew signal input
flabel metal4 s 215158 0 215218 200 0 FreeSans 480 90 0 0 um_ow[299]
port 604 nsew signal input
flabel metal4 s 14782 10680 14842 10880 0 FreeSans 480 90 0 0 um_ow[29]
port 605 nsew signal input
flabel metal4 s 16990 0 17050 200 0 FreeSans 480 90 0 0 um_ow[2]
port 606 nsew signal input
flabel metal4 s 214422 0 214482 200 0 FreeSans 480 90 0 0 um_ow[300]
port 607 nsew signal input
flabel metal4 s 213686 0 213746 200 0 FreeSans 480 90 0 0 um_ow[301]
port 608 nsew signal input
flabel metal4 s 212950 0 213010 200 0 FreeSans 480 90 0 0 um_ow[302]
port 609 nsew signal input
flabel metal4 s 212214 0 212274 200 0 FreeSans 480 90 0 0 um_ow[303]
port 610 nsew signal input
flabel metal4 s 211478 0 211538 200 0 FreeSans 480 90 0 0 um_ow[304]
port 611 nsew signal input
flabel metal4 s 210742 0 210802 200 0 FreeSans 480 90 0 0 um_ow[305]
port 612 nsew signal input
flabel metal4 s 210006 0 210066 200 0 FreeSans 480 90 0 0 um_ow[306]
port 613 nsew signal input
flabel metal4 s 209270 0 209330 200 0 FreeSans 480 90 0 0 um_ow[307]
port 614 nsew signal input
flabel metal4 s 208534 0 208594 200 0 FreeSans 480 90 0 0 um_ow[308]
port 615 nsew signal input
flabel metal4 s 207798 0 207858 200 0 FreeSans 480 90 0 0 um_ow[309]
port 616 nsew signal input
flabel metal4 s 14046 10680 14106 10880 0 FreeSans 480 90 0 0 um_ow[30]
port 617 nsew signal input
flabel metal4 s 207062 0 207122 200 0 FreeSans 480 90 0 0 um_ow[310]
port 618 nsew signal input
flabel metal4 s 206326 0 206386 200 0 FreeSans 480 90 0 0 um_ow[311]
port 619 nsew signal input
flabel metal4 s 223254 10680 223314 10880 0 FreeSans 480 90 0 0 um_ow[312]
port 620 nsew signal input
flabel metal4 s 222518 10680 222578 10880 0 FreeSans 480 90 0 0 um_ow[313]
port 621 nsew signal input
flabel metal4 s 221782 10680 221842 10880 0 FreeSans 480 90 0 0 um_ow[314]
port 622 nsew signal input
flabel metal4 s 221046 10680 221106 10880 0 FreeSans 480 90 0 0 um_ow[315]
port 623 nsew signal input
flabel metal4 s 220310 10680 220370 10880 0 FreeSans 480 90 0 0 um_ow[316]
port 624 nsew signal input
flabel metal4 s 219574 10680 219634 10880 0 FreeSans 480 90 0 0 um_ow[317]
port 625 nsew signal input
flabel metal4 s 218838 10680 218898 10880 0 FreeSans 480 90 0 0 um_ow[318]
port 626 nsew signal input
flabel metal4 s 218102 10680 218162 10880 0 FreeSans 480 90 0 0 um_ow[319]
port 627 nsew signal input
flabel metal4 s 13310 10680 13370 10880 0 FreeSans 480 90 0 0 um_ow[31]
port 628 nsew signal input
flabel metal4 s 217366 10680 217426 10880 0 FreeSans 480 90 0 0 um_ow[320]
port 629 nsew signal input
flabel metal4 s 216630 10680 216690 10880 0 FreeSans 480 90 0 0 um_ow[321]
port 630 nsew signal input
flabel metal4 s 215894 10680 215954 10880 0 FreeSans 480 90 0 0 um_ow[322]
port 631 nsew signal input
flabel metal4 s 215158 10680 215218 10880 0 FreeSans 480 90 0 0 um_ow[323]
port 632 nsew signal input
flabel metal4 s 214422 10680 214482 10880 0 FreeSans 480 90 0 0 um_ow[324]
port 633 nsew signal input
flabel metal4 s 213686 10680 213746 10880 0 FreeSans 480 90 0 0 um_ow[325]
port 634 nsew signal input
flabel metal4 s 212950 10680 213010 10880 0 FreeSans 480 90 0 0 um_ow[326]
port 635 nsew signal input
flabel metal4 s 212214 10680 212274 10880 0 FreeSans 480 90 0 0 um_ow[327]
port 636 nsew signal input
flabel metal4 s 211478 10680 211538 10880 0 FreeSans 480 90 0 0 um_ow[328]
port 637 nsew signal input
flabel metal4 s 210742 10680 210802 10880 0 FreeSans 480 90 0 0 um_ow[329]
port 638 nsew signal input
flabel metal4 s 12574 10680 12634 10880 0 FreeSans 480 90 0 0 um_ow[32]
port 639 nsew signal input
flabel metal4 s 210006 10680 210066 10880 0 FreeSans 480 90 0 0 um_ow[330]
port 640 nsew signal input
flabel metal4 s 209270 10680 209330 10880 0 FreeSans 480 90 0 0 um_ow[331]
port 641 nsew signal input
flabel metal4 s 208534 10680 208594 10880 0 FreeSans 480 90 0 0 um_ow[332]
port 642 nsew signal input
flabel metal4 s 207798 10680 207858 10880 0 FreeSans 480 90 0 0 um_ow[333]
port 643 nsew signal input
flabel metal4 s 207062 10680 207122 10880 0 FreeSans 480 90 0 0 um_ow[334]
port 644 nsew signal input
flabel metal4 s 206326 10680 206386 10880 0 FreeSans 480 90 0 0 um_ow[335]
port 645 nsew signal input
flabel metal4 s 257386 0 257446 200 0 FreeSans 480 90 0 0 um_ow[336]
port 646 nsew signal input
flabel metal4 s 256650 0 256710 200 0 FreeSans 480 90 0 0 um_ow[337]
port 647 nsew signal input
flabel metal4 s 255914 0 255974 200 0 FreeSans 480 90 0 0 um_ow[338]
port 648 nsew signal input
flabel metal4 s 255178 0 255238 200 0 FreeSans 480 90 0 0 um_ow[339]
port 649 nsew signal input
flabel metal4 s 11838 10680 11898 10880 0 FreeSans 480 90 0 0 um_ow[33]
port 650 nsew signal input
flabel metal4 s 254442 0 254502 200 0 FreeSans 480 90 0 0 um_ow[340]
port 651 nsew signal input
flabel metal4 s 253706 0 253766 200 0 FreeSans 480 90 0 0 um_ow[341]
port 652 nsew signal input
flabel metal4 s 252970 0 253030 200 0 FreeSans 480 90 0 0 um_ow[342]
port 653 nsew signal input
flabel metal4 s 252234 0 252294 200 0 FreeSans 480 90 0 0 um_ow[343]
port 654 nsew signal input
flabel metal4 s 251498 0 251558 200 0 FreeSans 480 90 0 0 um_ow[344]
port 655 nsew signal input
flabel metal4 s 250762 0 250822 200 0 FreeSans 480 90 0 0 um_ow[345]
port 656 nsew signal input
flabel metal4 s 250026 0 250086 200 0 FreeSans 480 90 0 0 um_ow[346]
port 657 nsew signal input
flabel metal4 s 249290 0 249350 200 0 FreeSans 480 90 0 0 um_ow[347]
port 658 nsew signal input
flabel metal4 s 248554 0 248614 200 0 FreeSans 480 90 0 0 um_ow[348]
port 659 nsew signal input
flabel metal4 s 247818 0 247878 200 0 FreeSans 480 90 0 0 um_ow[349]
port 660 nsew signal input
flabel metal4 s 11102 10680 11162 10880 0 FreeSans 480 90 0 0 um_ow[34]
port 661 nsew signal input
flabel metal4 s 247082 0 247142 200 0 FreeSans 480 90 0 0 um_ow[350]
port 662 nsew signal input
flabel metal4 s 246346 0 246406 200 0 FreeSans 480 90 0 0 um_ow[351]
port 663 nsew signal input
flabel metal4 s 245610 0 245670 200 0 FreeSans 480 90 0 0 um_ow[352]
port 664 nsew signal input
flabel metal4 s 244874 0 244934 200 0 FreeSans 480 90 0 0 um_ow[353]
port 665 nsew signal input
flabel metal4 s 244138 0 244198 200 0 FreeSans 480 90 0 0 um_ow[354]
port 666 nsew signal input
flabel metal4 s 243402 0 243462 200 0 FreeSans 480 90 0 0 um_ow[355]
port 667 nsew signal input
flabel metal4 s 242666 0 242726 200 0 FreeSans 480 90 0 0 um_ow[356]
port 668 nsew signal input
flabel metal4 s 241930 0 241990 200 0 FreeSans 480 90 0 0 um_ow[357]
port 669 nsew signal input
flabel metal4 s 241194 0 241254 200 0 FreeSans 480 90 0 0 um_ow[358]
port 670 nsew signal input
flabel metal4 s 240458 0 240518 200 0 FreeSans 480 90 0 0 um_ow[359]
port 671 nsew signal input
flabel metal4 s 10366 10680 10426 10880 0 FreeSans 480 90 0 0 um_ow[35]
port 672 nsew signal input
flabel metal4 s 257386 10680 257446 10880 0 FreeSans 480 90 0 0 um_ow[360]
port 673 nsew signal input
flabel metal4 s 256650 10680 256710 10880 0 FreeSans 480 90 0 0 um_ow[361]
port 674 nsew signal input
flabel metal4 s 255914 10680 255974 10880 0 FreeSans 480 90 0 0 um_ow[362]
port 675 nsew signal input
flabel metal4 s 255178 10680 255238 10880 0 FreeSans 480 90 0 0 um_ow[363]
port 676 nsew signal input
flabel metal4 s 254442 10680 254502 10880 0 FreeSans 480 90 0 0 um_ow[364]
port 677 nsew signal input
flabel metal4 s 253706 10680 253766 10880 0 FreeSans 480 90 0 0 um_ow[365]
port 678 nsew signal input
flabel metal4 s 252970 10680 253030 10880 0 FreeSans 480 90 0 0 um_ow[366]
port 679 nsew signal input
flabel metal4 s 252234 10680 252294 10880 0 FreeSans 480 90 0 0 um_ow[367]
port 680 nsew signal input
flabel metal4 s 251498 10680 251558 10880 0 FreeSans 480 90 0 0 um_ow[368]
port 681 nsew signal input
flabel metal4 s 250762 10680 250822 10880 0 FreeSans 480 90 0 0 um_ow[369]
port 682 nsew signal input
flabel metal4 s 9630 10680 9690 10880 0 FreeSans 480 90 0 0 um_ow[36]
port 683 nsew signal input
flabel metal4 s 250026 10680 250086 10880 0 FreeSans 480 90 0 0 um_ow[370]
port 684 nsew signal input
flabel metal4 s 249290 10680 249350 10880 0 FreeSans 480 90 0 0 um_ow[371]
port 685 nsew signal input
flabel metal4 s 248554 10680 248614 10880 0 FreeSans 480 90 0 0 um_ow[372]
port 686 nsew signal input
flabel metal4 s 247818 10680 247878 10880 0 FreeSans 480 90 0 0 um_ow[373]
port 687 nsew signal input
flabel metal4 s 247082 10680 247142 10880 0 FreeSans 480 90 0 0 um_ow[374]
port 688 nsew signal input
flabel metal4 s 246346 10680 246406 10880 0 FreeSans 480 90 0 0 um_ow[375]
port 689 nsew signal input
flabel metal4 s 245610 10680 245670 10880 0 FreeSans 480 90 0 0 um_ow[376]
port 690 nsew signal input
flabel metal4 s 244874 10680 244934 10880 0 FreeSans 480 90 0 0 um_ow[377]
port 691 nsew signal input
flabel metal4 s 244138 10680 244198 10880 0 FreeSans 480 90 0 0 um_ow[378]
port 692 nsew signal input
flabel metal4 s 243402 10680 243462 10880 0 FreeSans 480 90 0 0 um_ow[379]
port 693 nsew signal input
flabel metal4 s 8894 10680 8954 10880 0 FreeSans 480 90 0 0 um_ow[37]
port 694 nsew signal input
flabel metal4 s 242666 10680 242726 10880 0 FreeSans 480 90 0 0 um_ow[380]
port 695 nsew signal input
flabel metal4 s 241930 10680 241990 10880 0 FreeSans 480 90 0 0 um_ow[381]
port 696 nsew signal input
flabel metal4 s 241194 10680 241254 10880 0 FreeSans 480 90 0 0 um_ow[382]
port 697 nsew signal input
flabel metal4 s 240458 10680 240518 10880 0 FreeSans 480 90 0 0 um_ow[383]
port 698 nsew signal input
flabel metal4 s 8158 10680 8218 10880 0 FreeSans 480 90 0 0 um_ow[38]
port 699 nsew signal input
flabel metal4 s 7422 10680 7482 10880 0 FreeSans 480 90 0 0 um_ow[39]
port 700 nsew signal input
flabel metal4 s 16254 0 16314 200 0 FreeSans 480 90 0 0 um_ow[3]
port 701 nsew signal input
flabel metal4 s 6686 10680 6746 10880 0 FreeSans 480 90 0 0 um_ow[40]
port 702 nsew signal input
flabel metal4 s 5950 10680 6010 10880 0 FreeSans 480 90 0 0 um_ow[41]
port 703 nsew signal input
flabel metal4 s 5214 10680 5274 10880 0 FreeSans 480 90 0 0 um_ow[42]
port 704 nsew signal input
flabel metal4 s 4478 10680 4538 10880 0 FreeSans 480 90 0 0 um_ow[43]
port 705 nsew signal input
flabel metal4 s 3742 10680 3802 10880 0 FreeSans 480 90 0 0 um_ow[44]
port 706 nsew signal input
flabel metal4 s 3006 10680 3066 10880 0 FreeSans 480 90 0 0 um_ow[45]
port 707 nsew signal input
flabel metal4 s 2270 10680 2330 10880 0 FreeSans 480 90 0 0 um_ow[46]
port 708 nsew signal input
flabel metal4 s 1534 10680 1594 10880 0 FreeSans 480 90 0 0 um_ow[47]
port 709 nsew signal input
flabel metal4 s 52594 0 52654 200 0 FreeSans 480 90 0 0 um_ow[48]
port 710 nsew signal input
flabel metal4 s 51858 0 51918 200 0 FreeSans 480 90 0 0 um_ow[49]
port 711 nsew signal input
flabel metal4 s 15518 0 15578 200 0 FreeSans 480 90 0 0 um_ow[4]
port 712 nsew signal input
flabel metal4 s 51122 0 51182 200 0 FreeSans 480 90 0 0 um_ow[50]
port 713 nsew signal input
flabel metal4 s 50386 0 50446 200 0 FreeSans 480 90 0 0 um_ow[51]
port 714 nsew signal input
flabel metal4 s 49650 0 49710 200 0 FreeSans 480 90 0 0 um_ow[52]
port 715 nsew signal input
flabel metal4 s 48914 0 48974 200 0 FreeSans 480 90 0 0 um_ow[53]
port 716 nsew signal input
flabel metal4 s 48178 0 48238 200 0 FreeSans 480 90 0 0 um_ow[54]
port 717 nsew signal input
flabel metal4 s 47442 0 47502 200 0 FreeSans 480 90 0 0 um_ow[55]
port 718 nsew signal input
flabel metal4 s 46706 0 46766 200 0 FreeSans 480 90 0 0 um_ow[56]
port 719 nsew signal input
flabel metal4 s 45970 0 46030 200 0 FreeSans 480 90 0 0 um_ow[57]
port 720 nsew signal input
flabel metal4 s 45234 0 45294 200 0 FreeSans 480 90 0 0 um_ow[58]
port 721 nsew signal input
flabel metal4 s 44498 0 44558 200 0 FreeSans 480 90 0 0 um_ow[59]
port 722 nsew signal input
flabel metal4 s 14782 0 14842 200 0 FreeSans 480 90 0 0 um_ow[5]
port 723 nsew signal input
flabel metal4 s 43762 0 43822 200 0 FreeSans 480 90 0 0 um_ow[60]
port 724 nsew signal input
flabel metal4 s 43026 0 43086 200 0 FreeSans 480 90 0 0 um_ow[61]
port 725 nsew signal input
flabel metal4 s 42290 0 42350 200 0 FreeSans 480 90 0 0 um_ow[62]
port 726 nsew signal input
flabel metal4 s 41554 0 41614 200 0 FreeSans 480 90 0 0 um_ow[63]
port 727 nsew signal input
flabel metal4 s 40818 0 40878 200 0 FreeSans 480 90 0 0 um_ow[64]
port 728 nsew signal input
flabel metal4 s 40082 0 40142 200 0 FreeSans 480 90 0 0 um_ow[65]
port 729 nsew signal input
flabel metal4 s 39346 0 39406 200 0 FreeSans 480 90 0 0 um_ow[66]
port 730 nsew signal input
flabel metal4 s 38610 0 38670 200 0 FreeSans 480 90 0 0 um_ow[67]
port 731 nsew signal input
flabel metal4 s 37874 0 37934 200 0 FreeSans 480 90 0 0 um_ow[68]
port 732 nsew signal input
flabel metal4 s 37138 0 37198 200 0 FreeSans 480 90 0 0 um_ow[69]
port 733 nsew signal input
flabel metal4 s 14046 0 14106 200 0 FreeSans 480 90 0 0 um_ow[6]
port 734 nsew signal input
flabel metal4 s 36402 0 36462 200 0 FreeSans 480 90 0 0 um_ow[70]
port 735 nsew signal input
flabel metal4 s 35666 0 35726 200 0 FreeSans 480 90 0 0 um_ow[71]
port 736 nsew signal input
flabel metal4 s 52594 10680 52654 10880 0 FreeSans 480 90 0 0 um_ow[72]
port 737 nsew signal input
flabel metal4 s 51858 10680 51918 10880 0 FreeSans 480 90 0 0 um_ow[73]
port 738 nsew signal input
flabel metal4 s 51122 10680 51182 10880 0 FreeSans 480 90 0 0 um_ow[74]
port 739 nsew signal input
flabel metal4 s 50386 10680 50446 10880 0 FreeSans 480 90 0 0 um_ow[75]
port 740 nsew signal input
flabel metal4 s 49650 10680 49710 10880 0 FreeSans 480 90 0 0 um_ow[76]
port 741 nsew signal input
flabel metal4 s 48914 10680 48974 10880 0 FreeSans 480 90 0 0 um_ow[77]
port 742 nsew signal input
flabel metal4 s 48178 10680 48238 10880 0 FreeSans 480 90 0 0 um_ow[78]
port 743 nsew signal input
flabel metal4 s 47442 10680 47502 10880 0 FreeSans 480 90 0 0 um_ow[79]
port 744 nsew signal input
flabel metal4 s 13310 0 13370 200 0 FreeSans 480 90 0 0 um_ow[7]
port 745 nsew signal input
flabel metal4 s 46706 10680 46766 10880 0 FreeSans 480 90 0 0 um_ow[80]
port 746 nsew signal input
flabel metal4 s 45970 10680 46030 10880 0 FreeSans 480 90 0 0 um_ow[81]
port 747 nsew signal input
flabel metal4 s 45234 10680 45294 10880 0 FreeSans 480 90 0 0 um_ow[82]
port 748 nsew signal input
flabel metal4 s 44498 10680 44558 10880 0 FreeSans 480 90 0 0 um_ow[83]
port 749 nsew signal input
flabel metal4 s 43762 10680 43822 10880 0 FreeSans 480 90 0 0 um_ow[84]
port 750 nsew signal input
flabel metal4 s 43026 10680 43086 10880 0 FreeSans 480 90 0 0 um_ow[85]
port 751 nsew signal input
flabel metal4 s 42290 10680 42350 10880 0 FreeSans 480 90 0 0 um_ow[86]
port 752 nsew signal input
flabel metal4 s 41554 10680 41614 10880 0 FreeSans 480 90 0 0 um_ow[87]
port 753 nsew signal input
flabel metal4 s 40818 10680 40878 10880 0 FreeSans 480 90 0 0 um_ow[88]
port 754 nsew signal input
flabel metal4 s 40082 10680 40142 10880 0 FreeSans 480 90 0 0 um_ow[89]
port 755 nsew signal input
flabel metal4 s 12574 0 12634 200 0 FreeSans 480 90 0 0 um_ow[8]
port 756 nsew signal input
flabel metal4 s 39346 10680 39406 10880 0 FreeSans 480 90 0 0 um_ow[90]
port 757 nsew signal input
flabel metal4 s 38610 10680 38670 10880 0 FreeSans 480 90 0 0 um_ow[91]
port 758 nsew signal input
flabel metal4 s 37874 10680 37934 10880 0 FreeSans 480 90 0 0 um_ow[92]
port 759 nsew signal input
flabel metal4 s 37138 10680 37198 10880 0 FreeSans 480 90 0 0 um_ow[93]
port 760 nsew signal input
flabel metal4 s 36402 10680 36462 10880 0 FreeSans 480 90 0 0 um_ow[94]
port 761 nsew signal input
flabel metal4 s 35666 10680 35726 10880 0 FreeSans 480 90 0 0 um_ow[95]
port 762 nsew signal input
flabel metal4 s 86726 0 86786 200 0 FreeSans 480 90 0 0 um_ow[96]
port 763 nsew signal input
flabel metal4 s 85990 0 86050 200 0 FreeSans 480 90 0 0 um_ow[97]
port 764 nsew signal input
flabel metal4 s 85254 0 85314 200 0 FreeSans 480 90 0 0 um_ow[98]
port 765 nsew signal input
flabel metal4 s 84518 0 84578 200 0 FreeSans 480 90 0 0 um_ow[99]
port 766 nsew signal input
flabel metal4 s 11838 0 11898 200 0 FreeSans 480 90 0 0 um_ow[9]
port 767 nsew signal input
flabel metal4 s 34742 1040 35062 9840 0 FreeSans 1920 90 0 0 vccd1
port 768 nsew power bidirectional
flabel metal4 s 102339 1040 102659 9840 0 FreeSans 1920 90 0 0 vccd1
port 768 nsew power bidirectional
flabel metal4 s 169936 1040 170256 9840 0 FreeSans 1920 90 0 0 vccd1
port 768 nsew power bidirectional
flabel metal4 s 237533 1040 237853 9840 0 FreeSans 1920 90 0 0 vccd1
port 768 nsew power bidirectional
flabel metal4 s 68540 1040 68860 9840 0 FreeSans 1920 90 0 0 vssd1
port 769 nsew ground bidirectional
flabel metal4 s 136137 1040 136457 9840 0 FreeSans 1920 90 0 0 vssd1
port 769 nsew ground bidirectional
flabel metal4 s 203734 1040 204054 9840 0 FreeSans 1920 90 0 0 vssd1
port 769 nsew ground bidirectional
flabel metal4 s 271331 1040 271651 9840 0 FreeSans 1920 90 0 0 vssd1
port 769 nsew ground bidirectional
rlabel metal1 136298 9248 136298 9248 0 vccd1
rlabel via1 136377 9792 136377 9792 0 vssd1
rlabel metal1 229126 5780 229126 5780 0 _000_
rlabel metal1 267628 4590 267628 4590 0 _001_
rlabel metal1 267444 4590 267444 4590 0 _002_
rlabel metal1 269514 4522 269514 4522 0 _003_
rlabel metal2 270894 6290 270894 6290 0 _004_
rlabel metal2 270802 6290 270802 6290 0 _005_
rlabel metal1 269468 4794 269468 4794 0 _006_
rlabel metal1 268916 8058 268916 8058 0 _007_
rlabel metal1 270304 4522 270304 4522 0 _008_
rlabel metal1 270756 4794 270756 4794 0 _009_
rlabel via2 80362 5253 80362 5253 0 _010_
rlabel metal2 79074 6018 79074 6018 0 _011_
rlabel metal1 80500 5542 80500 5542 0 _012_
rlabel metal1 79396 6358 79396 6358 0 _013_
rlabel metal2 79626 6800 79626 6800 0 _014_
rlabel metal2 77326 4692 77326 4692 0 _015_
rlabel metal2 79442 7174 79442 7174 0 _016_
rlabel metal1 99866 2006 99866 2006 0 _017_
rlabel metal2 100142 5950 100142 5950 0 _018_
rlabel metal1 100280 6426 100280 6426 0 _019_
rlabel metal2 122590 4794 122590 4794 0 _020_
rlabel metal2 120290 6766 120290 6766 0 _021_
rlabel metal2 162978 4012 162978 4012 0 _022_
rlabel metal2 189198 5848 189198 5848 0 _023_
rlabel metal2 169786 7140 169786 7140 0 _024_
rlabel metal2 190026 4590 190026 4590 0 _025_
rlabel metal2 189382 6596 189382 6596 0 _026_
rlabel metal1 231104 3502 231104 3502 0 _027_
rlabel via1 230882 5610 230882 5610 0 _028_
rlabel metal2 230138 7174 230138 7174 0 _029_
rlabel metal2 235658 4590 235658 4590 0 _030_
rlabel metal1 231196 5882 231196 5882 0 _031_
rlabel metal3 272305 9588 272305 9588 0 addr[0]
rlabel metal3 272213 9452 272213 9452 0 addr[1]
rlabel metal3 270672 9316 270672 9316 0 addr[2]
rlabel metal3 270212 9180 270212 9180 0 addr[3]
rlabel metal3 270258 9044 270258 9044 0 addr[4]
rlabel metal1 84180 4182 84180 4182 0 col\[0\].genblk1.mux4_I\[0\].x
rlabel metal2 81926 5151 81926 5151 0 col\[0\].genblk1.mux4_I\[10\].x
rlabel via2 91770 5117 91770 5117 0 col\[0\].genblk1.mux4_I\[11\].x
rlabel metal2 92690 5933 92690 5933 0 col\[0\].genblk1.mux4_I\[12\].x
rlabel metal2 60766 3961 60766 3961 0 col\[0\].genblk1.mux4_I\[13\].x
rlabel metal2 94346 4335 94346 4335 0 col\[0\].genblk1.mux4_I\[14\].x
rlabel metal1 79350 3400 79350 3400 0 col\[0\].genblk1.mux4_I\[15\].x
rlabel metal2 86066 3230 86066 3230 0 col\[0\].genblk1.mux4_I\[16\].x
rlabel via2 41170 2907 41170 2907 0 col\[0\].genblk1.mux4_I\[17\].x
rlabel via2 40342 1819 40342 1819 0 col\[0\].genblk1.mux4_I\[18\].x
rlabel metal2 86618 3247 86618 3247 0 col\[0\].genblk1.mux4_I\[19\].x
rlabel metal2 81466 3604 81466 3604 0 col\[0\].genblk1.mux4_I\[1\].x
rlabel metal1 64860 4624 64860 4624 0 col\[0\].genblk1.mux4_I\[20\].x
rlabel metal2 38226 2329 38226 2329 0 col\[0\].genblk1.mux4_I\[21\].x
rlabel metal1 83122 2346 83122 2346 0 col\[0\].genblk1.mux4_I\[22\].x
rlabel via2 36846 1717 36846 1717 0 col\[0\].genblk1.mux4_I\[23\].x
rlabel via1 67022 3485 67022 3485 0 col\[0\].genblk1.mux4_I\[2\].x
rlabel metal1 83398 5644 83398 5644 0 col\[0\].genblk1.mux4_I\[3\].x
rlabel metal2 78154 4828 78154 4828 0 col\[0\].genblk1.mux4_I\[4\].x
rlabel metal1 81466 5270 81466 5270 0 col\[0\].genblk1.mux4_I\[5\].x
rlabel metal2 79258 3570 79258 3570 0 col\[0\].genblk1.mux4_I\[6\].x
rlabel metal2 87906 5678 87906 5678 0 col\[0\].genblk1.mux4_I\[7\].x
rlabel metal1 89470 5100 89470 5100 0 col\[0\].genblk1.mux4_I\[8\].x
rlabel metal1 79350 6120 79350 6120 0 col\[0\].genblk1.mux4_I\[9\].x
rlabel metal2 81466 5185 81466 5185 0 col\[0\].genblk1.tbuf_row_ena_I.t
rlabel metal1 94714 4590 94714 4590 0 col\[0\].genblk1.tbuf_row_ena_I.tx
rlabel metal1 86802 4114 86802 4114 0 col\[0\].genblk1.tbuf_spine_ow_I\[0\].z
rlabel metal2 95266 5491 95266 5491 0 col\[0\].genblk1.tbuf_spine_ow_I\[10\].z
rlabel metal2 214682 5610 214682 5610 0 col\[0\].genblk1.tbuf_spine_ow_I\[11\].z
rlabel metal1 214774 6834 214774 6834 0 col\[0\].genblk1.tbuf_spine_ow_I\[12\].z
rlabel metal1 214314 4556 214314 4556 0 col\[0\].genblk1.tbuf_spine_ow_I\[13\].z
rlabel metal3 166244 1768 166244 1768 0 col\[0\].genblk1.tbuf_spine_ow_I\[14\].z
rlabel metal1 214176 4522 214176 4522 0 col\[0\].genblk1.tbuf_spine_ow_I\[15\].z
rlabel metal2 212382 3723 212382 3723 0 col\[0\].genblk1.tbuf_spine_ow_I\[16\].z
rlabel metal1 213026 3910 213026 3910 0 col\[0\].genblk1.tbuf_spine_ow_I\[17\].z
rlabel metal2 210910 3349 210910 3349 0 col\[0\].genblk1.tbuf_spine_ow_I\[18\].z
rlabel metal2 210082 4318 210082 4318 0 col\[0\].genblk1.tbuf_spine_ow_I\[19\].z
rlabel metal2 83950 2193 83950 2193 0 col\[0\].genblk1.tbuf_spine_ow_I\[1\].z
rlabel metal2 86618 5933 86618 5933 0 col\[0\].genblk1.tbuf_spine_ow_I\[20\].z
rlabel metal1 132480 2992 132480 2992 0 col\[0\].genblk1.tbuf_spine_ow_I\[21\].z
rlabel metal2 133262 1904 133262 1904 0 col\[0\].genblk1.tbuf_spine_ow_I\[22\].z
rlabel metal2 86066 1598 86066 1598 0 col\[0\].genblk1.tbuf_spine_ow_I\[23\].z
rlabel metal1 83030 3570 83030 3570 0 col\[0\].genblk1.tbuf_spine_ow_I\[2\].z
rlabel metal1 82938 5542 82938 5542 0 col\[0\].genblk1.tbuf_spine_ow_I\[3\].z
rlabel metal1 83582 4488 83582 4488 0 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z
rlabel metal1 83582 5134 83582 5134 0 col\[0\].genblk1.tbuf_spine_ow_I\[5\].z
rlabel metal1 213118 5576 213118 5576 0 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z
rlabel metal2 214590 5576 214590 5576 0 col\[0\].genblk1.tbuf_spine_ow_I\[7\].z
rlabel metal1 88826 5270 88826 5270 0 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z
rlabel via2 250654 4675 250654 4675 0 col\[0\].genblk1.tbuf_spine_ow_I\[9\].z
rlabel metal2 32522 2176 32522 2176 0 col\[0\].zbuf_bot_ena_I.e
rlabel metal1 32936 1938 32936 1938 0 col\[0\].zbuf_bot_ena_I.z
rlabel metal1 170292 8806 170292 8806 0 col\[0\].zbuf_bot_iw_I\[0\].a
rlabel metal2 32338 1802 32338 1802 0 col\[0\].zbuf_bot_iw_I\[0\].z
rlabel metal2 226274 1088 226274 1088 0 col\[0\].zbuf_bot_iw_I\[10\].a
rlabel metal1 25530 2618 25530 2618 0 col\[0\].zbuf_bot_iw_I\[10\].z
rlabel metal2 187726 8313 187726 8313 0 col\[0\].zbuf_bot_iw_I\[11\].a
rlabel metal2 23782 1530 23782 1530 0 col\[0\].zbuf_bot_iw_I\[11\].z
rlabel metal2 224802 391 224802 391 0 col\[0\].zbuf_bot_iw_I\[12\].a
rlabel metal1 24104 3026 24104 3026 0 col\[0\].zbuf_bot_iw_I\[12\].z
rlabel metal2 175858 3298 175858 3298 0 col\[0\].zbuf_bot_iw_I\[13\].a
rlabel metal1 24564 3366 24564 3366 0 col\[0\].zbuf_bot_iw_I\[13\].z
rlabel metal2 158654 1445 158654 1445 0 col\[0\].zbuf_bot_iw_I\[14\].a
rlabel metal1 25438 2006 25438 2006 0 col\[0\].zbuf_bot_iw_I\[14\].z
rlabel metal2 158010 2006 158010 2006 0 col\[0\].zbuf_bot_iw_I\[15\].a
rlabel metal1 25622 1258 25622 1258 0 col\[0\].zbuf_bot_iw_I\[15\].z
rlabel metal3 249780 680 249780 680 0 col\[0\].zbuf_bot_iw_I\[16\].a
rlabel metal1 26358 2006 26358 2006 0 col\[0\].zbuf_bot_iw_I\[16\].z
rlabel metal2 169326 1020 169326 1020 0 col\[0\].zbuf_bot_iw_I\[17\].a
rlabel metal1 27508 2006 27508 2006 0 col\[0\].zbuf_bot_iw_I\[17\].z
rlabel metal1 192510 9588 192510 9588 0 col\[0\].zbuf_bot_iw_I\[1\].a
rlabel metal2 31786 1530 31786 1530 0 col\[0\].zbuf_bot_iw_I\[1\].z
rlabel metal2 167394 8670 167394 8670 0 col\[0\].zbuf_bot_iw_I\[2\].a
rlabel metal2 30590 1530 30590 1530 0 col\[0\].zbuf_bot_iw_I\[2\].z
rlabel metal2 212474 8364 212474 8364 0 col\[0\].zbuf_bot_iw_I\[3\].a
rlabel metal2 29762 1530 29762 1530 0 col\[0\].zbuf_bot_iw_I\[3\].z
rlabel metal2 266846 9758 266846 9758 0 col\[0\].zbuf_bot_iw_I\[4\].a
rlabel metal2 28934 1530 28934 1530 0 col\[0\].zbuf_bot_iw_I\[4\].z
rlabel metal1 266432 8534 266432 8534 0 col\[0\].zbuf_bot_iw_I\[5\].a
rlabel metal1 28474 1530 28474 1530 0 col\[0\].zbuf_bot_iw_I\[5\].z
rlabel metal2 265190 7344 265190 7344 0 col\[0\].zbuf_bot_iw_I\[6\].a
rlabel metal1 27416 3502 27416 3502 0 col\[0\].zbuf_bot_iw_I\[6\].z
rlabel metal2 264822 9894 264822 9894 0 col\[0\].zbuf_bot_iw_I\[7\].a
rlabel metal1 26818 2618 26818 2618 0 col\[0\].zbuf_bot_iw_I\[7\].z
rlabel metal1 264408 8466 264408 8466 0 col\[0\].zbuf_bot_iw_I\[8\].a
rlabel metal1 26036 3502 26036 3502 0 col\[0\].zbuf_bot_iw_I\[8\].z
rlabel metal2 162242 9554 162242 9554 0 col\[0\].zbuf_bot_iw_I\[9\].a
rlabel metal1 28060 2618 28060 2618 0 col\[0\].zbuf_bot_iw_I\[9\].z
rlabel metal2 37030 8058 37030 8058 0 col\[0\].zbuf_top_ena_I.e
rlabel metal2 32706 9078 32706 9078 0 col\[0\].zbuf_top_ena_I.z
rlabel metal1 32844 8942 32844 8942 0 col\[0\].zbuf_top_iw_I\[0\].z
rlabel metal2 25254 8194 25254 8194 0 col\[0\].zbuf_top_iw_I\[10\].z
rlabel metal1 24932 6766 24932 6766 0 col\[0\].zbuf_top_iw_I\[11\].z
rlabel metal2 24518 8364 24518 8364 0 col\[0\].zbuf_top_iw_I\[12\].z
rlabel metal1 24196 9146 24196 9146 0 col\[0\].zbuf_top_iw_I\[13\].z
rlabel metal1 25392 7514 25392 7514 0 col\[0\].zbuf_top_iw_I\[14\].z
rlabel metal1 25760 8534 25760 8534 0 col\[0\].zbuf_top_iw_I\[15\].z
rlabel metal2 26450 8194 26450 8194 0 col\[0\].zbuf_top_iw_I\[16\].z
rlabel metal1 27278 8568 27278 8568 0 col\[0\].zbuf_top_iw_I\[17\].z
rlabel metal2 31142 8636 31142 8636 0 col\[0\].zbuf_top_iw_I\[1\].z
rlabel metal2 30314 8636 30314 8636 0 col\[0\].zbuf_top_iw_I\[2\].z
rlabel metal2 29486 8636 29486 8636 0 col\[0\].zbuf_top_iw_I\[3\].z
rlabel metal2 28750 9078 28750 9078 0 col\[0\].zbuf_top_iw_I\[4\].z
rlabel metal2 28198 8602 28198 8602 0 col\[0\].zbuf_top_iw_I\[5\].z
rlabel metal2 28934 8738 28934 8738 0 col\[0\].zbuf_top_iw_I\[6\].z
rlabel metal2 26542 7242 26542 7242 0 col\[0\].zbuf_top_iw_I\[7\].z
rlabel metal1 27416 8466 27416 8466 0 col\[0\].zbuf_top_iw_I\[8\].z
rlabel metal2 27830 7548 27830 7548 0 col\[0\].zbuf_top_iw_I\[9\].z
rlabel metal1 63434 1904 63434 1904 0 col\[1\].zbuf_bot_ena_I.e
rlabel metal1 67160 1938 67160 1938 0 col\[1\].zbuf_bot_ena_I.z
rlabel metal2 66010 1530 66010 1530 0 col\[1\].zbuf_bot_iw_I\[0\].z
rlabel metal2 58466 1530 58466 1530 0 col\[1\].zbuf_bot_iw_I\[10\].z
rlabel metal2 57546 2244 57546 2244 0 col\[1\].zbuf_bot_iw_I\[11\].z
rlabel metal2 56902 1530 56902 1530 0 col\[1\].zbuf_bot_iw_I\[12\].z
rlabel metal2 56074 1530 56074 1530 0 col\[1\].zbuf_bot_iw_I\[13\].z
rlabel metal2 55062 2210 55062 2210 0 col\[1\].zbuf_bot_iw_I\[14\].z
rlabel metal2 54234 2210 54234 2210 0 col\[1\].zbuf_bot_iw_I\[15\].z
rlabel metal1 53636 1258 53636 1258 0 col\[1\].zbuf_bot_iw_I\[16\].z
rlabel metal1 53544 1326 53544 1326 0 col\[1\].zbuf_bot_iw_I\[17\].z
rlabel metal2 65274 2244 65274 2244 0 col\[1\].zbuf_bot_iw_I\[1\].z
rlabel metal2 64354 1530 64354 1530 0 col\[1\].zbuf_bot_iw_I\[2\].z
rlabel metal2 63618 1530 63618 1530 0 col\[1\].zbuf_bot_iw_I\[3\].z
rlabel metal2 62698 2244 62698 2244 0 col\[1\].zbuf_bot_iw_I\[4\].z
rlabel metal1 62008 1326 62008 1326 0 col\[1\].zbuf_bot_iw_I\[5\].z
rlabel metal2 61410 1530 61410 1530 0 col\[1\].zbuf_bot_iw_I\[6\].z
rlabel metal2 60674 1530 60674 1530 0 col\[1\].zbuf_bot_iw_I\[7\].z
rlabel metal2 60030 1972 60030 1972 0 col\[1\].zbuf_bot_iw_I\[8\].z
rlabel metal2 59294 2244 59294 2244 0 col\[1\].zbuf_bot_iw_I\[9\].z
rlabel metal1 66884 8942 66884 8942 0 col\[1\].zbuf_top_ena_I.e
rlabel metal2 67022 9044 67022 9044 0 col\[1\].zbuf_top_ena_I.z
rlabel metal2 66378 9350 66378 9350 0 col\[1\].zbuf_top_iw_I\[0\].z
rlabel metal2 58466 8636 58466 8636 0 col\[1\].zbuf_top_iw_I\[10\].z
rlabel metal2 57546 9350 57546 9350 0 col\[1\].zbuf_top_iw_I\[11\].z
rlabel metal2 56902 8636 56902 8636 0 col\[1\].zbuf_top_iw_I\[12\].z
rlabel metal2 56074 8636 56074 8636 0 col\[1\].zbuf_top_iw_I\[13\].z
rlabel metal2 55338 8636 55338 8636 0 col\[1\].zbuf_top_iw_I\[14\].z
rlabel metal2 54602 8636 54602 8636 0 col\[1\].zbuf_top_iw_I\[15\].z
rlabel metal2 54142 9078 54142 9078 0 col\[1\].zbuf_top_iw_I\[16\].z
rlabel metal1 53222 8942 53222 8942 0 col\[1\].zbuf_top_iw_I\[17\].z
rlabel metal2 65274 8636 65274 8636 0 col\[1\].zbuf_top_iw_I\[1\].z
rlabel metal2 64446 8636 64446 8636 0 col\[1\].zbuf_top_iw_I\[2\].z
rlabel metal2 63618 8636 63618 8636 0 col\[1\].zbuf_top_iw_I\[3\].z
rlabel metal2 62790 9350 62790 9350 0 col\[1\].zbuf_top_iw_I\[4\].z
rlabel metal2 62146 8636 62146 8636 0 col\[1\].zbuf_top_iw_I\[5\].z
rlabel metal2 61410 8636 61410 8636 0 col\[1\].zbuf_top_iw_I\[6\].z
rlabel metal2 60766 9078 60766 9078 0 col\[1\].zbuf_top_iw_I\[7\].z
rlabel metal2 60030 9350 60030 9350 0 col\[1\].zbuf_top_iw_I\[8\].z
rlabel metal2 59202 9350 59202 9350 0 col\[1\].zbuf_top_iw_I\[9\].z
rlabel metal1 122222 4658 122222 4658 0 col\[2\].genblk1.mux4_I\[0\].x
rlabel metal1 110446 6290 110446 6290 0 col\[2\].genblk1.mux4_I\[10\].x
rlabel metal2 109066 6086 109066 6086 0 col\[2\].genblk1.mux4_I\[11\].x
rlabel metal1 106674 6290 106674 6290 0 col\[2\].genblk1.mux4_I\[12\].x
rlabel metal2 110262 3468 110262 3468 0 col\[2\].genblk1.mux4_I\[13\].x
rlabel metal2 108882 4012 108882 4012 0 col\[2\].genblk1.mux4_I\[14\].x
rlabel metal1 108238 2482 108238 2482 0 col\[2\].genblk1.mux4_I\[15\].x
rlabel metal2 107134 3468 107134 3468 0 col\[2\].genblk1.mux4_I\[16\].x
rlabel metal1 104972 3570 104972 3570 0 col\[2\].genblk1.mux4_I\[17\].x
rlabel metal1 104006 2958 104006 2958 0 col\[2\].genblk1.mux4_I\[18\].x
rlabel metal2 101522 3332 101522 3332 0 col\[2\].genblk1.mux4_I\[19\].x
rlabel metal2 121026 3842 121026 3842 0 col\[2\].genblk1.mux4_I\[1\].x
rlabel metal2 101798 6460 101798 6460 0 col\[2\].genblk1.mux4_I\[20\].x
rlabel metal2 98762 3332 98762 3332 0 col\[2\].genblk1.mux4_I\[21\].x
rlabel metal2 98578 3332 98578 3332 0 col\[2\].genblk1.mux4_I\[22\].x
rlabel metal2 98486 2924 98486 2924 0 col\[2\].genblk1.mux4_I\[23\].x
rlabel metal1 120842 3026 120842 3026 0 col\[2\].genblk1.mux4_I\[2\].x
rlabel metal1 119692 5338 119692 5338 0 col\[2\].genblk1.mux4_I\[3\].x
rlabel metal2 116794 3876 116794 3876 0 col\[2\].genblk1.mux4_I\[4\].x
rlabel metal2 116518 3468 116518 3468 0 col\[2\].genblk1.mux4_I\[5\].x
rlabel metal2 114218 4624 114218 4624 0 col\[2\].genblk1.mux4_I\[6\].x
rlabel metal1 113896 4658 113896 4658 0 col\[2\].genblk1.mux4_I\[7\].x
rlabel metal1 111734 4726 111734 4726 0 col\[2\].genblk1.mux4_I\[8\].x
rlabel metal2 112470 7038 112470 7038 0 col\[2\].genblk1.mux4_I\[9\].x
rlabel metal2 150282 6511 150282 6511 0 col\[2\].genblk1.tbuf_row_ena_I.t
rlabel metal1 101246 5338 101246 5338 0 col\[2\].genblk1.tbuf_row_ena_I.tx
rlabel metal1 89286 1904 89286 1904 0 col\[2\].zbuf_bot_ena_I.e
rlabel metal1 100924 1938 100924 1938 0 col\[2\].zbuf_bot_ena_I.z
rlabel metal1 100556 1326 100556 1326 0 col\[2\].zbuf_bot_iw_I\[0\].z
rlabel metal2 92782 2244 92782 2244 0 col\[2\].zbuf_bot_iw_I\[10\].z
rlabel metal2 92046 1530 92046 1530 0 col\[2\].zbuf_bot_iw_I\[11\].z
rlabel metal2 91126 2244 91126 2244 0 col\[2\].zbuf_bot_iw_I\[12\].z
rlabel metal2 90482 1530 90482 1530 0 col\[2\].zbuf_bot_iw_I\[13\].z
rlabel metal2 89930 2176 89930 2176 0 col\[2\].zbuf_bot_iw_I\[14\].z
rlabel metal1 88826 1938 88826 1938 0 col\[2\].zbuf_bot_iw_I\[15\].z
rlabel metal1 89332 1326 89332 1326 0 col\[2\].zbuf_bot_iw_I\[16\].z
rlabel metal1 88412 1326 88412 1326 0 col\[2\].zbuf_bot_iw_I\[17\].z
rlabel metal1 101246 1870 101246 1870 0 col\[2\].zbuf_bot_iw_I\[1\].z
rlabel metal1 98072 1326 98072 1326 0 col\[2\].zbuf_bot_iw_I\[2\].z
rlabel metal1 97060 1326 97060 1326 0 col\[2\].zbuf_bot_iw_I\[3\].z
rlabel metal1 96278 1326 96278 1326 0 col\[2\].zbuf_bot_iw_I\[4\].z
rlabel metal2 96278 2244 96278 2244 0 col\[2\].zbuf_bot_iw_I\[5\].z
rlabel metal2 95450 2244 95450 2244 0 col\[2\].zbuf_bot_iw_I\[6\].z
rlabel metal1 94806 1530 94806 1530 0 col\[2\].zbuf_bot_iw_I\[7\].z
rlabel metal1 94116 2074 94116 2074 0 col\[2\].zbuf_bot_iw_I\[8\].z
rlabel metal2 93334 1530 93334 1530 0 col\[2\].zbuf_bot_iw_I\[9\].z
rlabel metal2 98118 9316 98118 9316 0 col\[2\].zbuf_top_ena_I.e
rlabel metal2 100234 9078 100234 9078 0 col\[2\].zbuf_top_ena_I.z
rlabel metal2 100694 8636 100694 8636 0 col\[2\].zbuf_top_iw_I\[0\].z
rlabel metal2 93150 8058 93150 8058 0 col\[2\].zbuf_top_iw_I\[10\].z
rlabel metal2 92414 8636 92414 8636 0 col\[2\].zbuf_top_iw_I\[11\].z
rlabel metal2 91678 8636 91678 8636 0 col\[2\].zbuf_top_iw_I\[12\].z
rlabel metal2 90942 8636 90942 8636 0 col\[2\].zbuf_top_iw_I\[13\].z
rlabel metal2 90206 9350 90206 9350 0 col\[2\].zbuf_top_iw_I\[14\].z
rlabel metal2 90114 8058 90114 8058 0 col\[2\].zbuf_top_iw_I\[15\].z
rlabel metal1 88274 8976 88274 8976 0 col\[2\].zbuf_top_iw_I\[16\].z
rlabel metal2 88826 8908 88826 8908 0 col\[2\].zbuf_top_iw_I\[17\].z
rlabel metal2 99406 8602 99406 8602 0 col\[2\].zbuf_top_iw_I\[1\].z
rlabel metal2 98486 8636 98486 8636 0 col\[2\].zbuf_top_iw_I\[2\].z
rlabel metal2 98026 9350 98026 9350 0 col\[2\].zbuf_top_iw_I\[3\].z
rlabel metal2 97290 8636 97290 8636 0 col\[2\].zbuf_top_iw_I\[4\].z
rlabel metal2 96830 9078 96830 9078 0 col\[2\].zbuf_top_iw_I\[5\].z
rlabel metal2 96186 9350 96186 9350 0 col\[2\].zbuf_top_iw_I\[6\].z
rlabel metal2 95174 8636 95174 8636 0 col\[2\].zbuf_top_iw_I\[7\].z
rlabel metal2 94438 8636 94438 8636 0 col\[2\].zbuf_top_iw_I\[8\].z
rlabel metal2 93702 9248 93702 9248 0 col\[2\].zbuf_top_iw_I\[9\].z
rlabel metal1 121440 1938 121440 1938 0 col\[3\].zbuf_bot_ena_I.e
rlabel metal1 134918 1938 134918 1938 0 col\[3\].zbuf_bot_ena_I.z
rlabel metal2 134366 1938 134366 1938 0 col\[3\].zbuf_bot_iw_I\[0\].z
rlabel metal1 126960 1326 126960 1326 0 col\[3\].zbuf_bot_iw_I\[10\].z
rlabel metal2 126270 2244 126270 2244 0 col\[3\].zbuf_bot_iw_I\[11\].z
rlabel metal2 125442 1530 125442 1530 0 col\[3\].zbuf_bot_iw_I\[12\].z
rlabel metal2 124522 2244 124522 2244 0 col\[3\].zbuf_bot_iw_I\[13\].z
rlabel metal2 123786 1530 123786 1530 0 col\[3\].zbuf_bot_iw_I\[14\].z
rlabel metal2 122958 1530 122958 1530 0 col\[3\].zbuf_bot_iw_I\[15\].z
rlabel metal2 122038 2244 122038 2244 0 col\[3\].zbuf_bot_iw_I\[16\].z
rlabel metal1 121440 1326 121440 1326 0 col\[3\].zbuf_bot_iw_I\[17\].z
rlabel metal2 133630 2210 133630 2210 0 col\[3\].zbuf_bot_iw_I\[1\].z
rlabel metal2 133354 1938 133354 1938 0 col\[3\].zbuf_bot_iw_I\[2\].z
rlabel metal2 132618 1530 132618 1530 0 col\[3\].zbuf_bot_iw_I\[3\].z
rlabel metal2 131698 2244 131698 2244 0 col\[3\].zbuf_bot_iw_I\[4\].z
rlabel metal2 130686 1530 130686 1530 0 col\[3\].zbuf_bot_iw_I\[5\].z
rlabel metal2 129674 2244 129674 2244 0 col\[3\].zbuf_bot_iw_I\[6\].z
rlabel metal2 129122 1530 129122 1530 0 col\[3\].zbuf_bot_iw_I\[7\].z
rlabel metal2 128662 1870 128662 1870 0 col\[3\].zbuf_bot_iw_I\[8\].z
rlabel metal2 127926 2244 127926 2244 0 col\[3\].zbuf_bot_iw_I\[9\].z
rlabel metal2 129306 9180 129306 9180 0 col\[3\].zbuf_top_ena_I.e
rlabel metal2 134550 8772 134550 8772 0 col\[3\].zbuf_top_ena_I.z
rlabel metal2 134274 9316 134274 9316 0 col\[3\].zbuf_top_iw_I\[0\].z
rlabel metal2 126914 8636 126914 8636 0 col\[3\].zbuf_top_iw_I\[10\].z
rlabel metal2 126178 8636 126178 8636 0 col\[3\].zbuf_top_iw_I\[11\].z
rlabel metal2 125442 8636 125442 8636 0 col\[3\].zbuf_top_iw_I\[12\].z
rlabel metal2 124614 9350 124614 9350 0 col\[3\].zbuf_top_iw_I\[13\].z
rlabel metal2 123786 8636 123786 8636 0 col\[3\].zbuf_top_iw_I\[14\].z
rlabel metal2 123050 8636 123050 8636 0 col\[3\].zbuf_top_iw_I\[15\].z
rlabel metal1 122222 9146 122222 9146 0 col\[3\].zbuf_top_iw_I\[16\].z
rlabel metal1 121394 8602 121394 8602 0 col\[3\].zbuf_top_iw_I\[17\].z
rlabel metal2 133446 9316 133446 9316 0 col\[3\].zbuf_top_iw_I\[1\].z
rlabel metal2 132894 8058 132894 8058 0 col\[3\].zbuf_top_iw_I\[2\].z
rlabel metal2 132158 8636 132158 8636 0 col\[3\].zbuf_top_iw_I\[3\].z
rlabel metal2 131422 9350 131422 9350 0 col\[3\].zbuf_top_iw_I\[4\].z
rlabel metal1 131192 8466 131192 8466 0 col\[3\].zbuf_top_iw_I\[5\].z
rlabel metal1 129398 9588 129398 9588 0 col\[3\].zbuf_top_iw_I\[6\].z
rlabel metal1 129076 8602 129076 8602 0 col\[3\].zbuf_top_iw_I\[7\].z
rlabel metal1 127650 8976 127650 8976 0 col\[3\].zbuf_top_iw_I\[8\].z
rlabel metal2 128018 9078 128018 9078 0 col\[3\].zbuf_top_iw_I\[9\].z
rlabel metal1 160632 3706 160632 3706 0 col\[4\].genblk1.mux4_I\[0\].x
rlabel metal1 150466 6290 150466 6290 0 col\[4\].genblk1.mux4_I\[10\].x
rlabel metal2 148258 6188 148258 6188 0 col\[4\].genblk1.mux4_I\[11\].x
rlabel metal1 146510 6324 146510 6324 0 col\[4\].genblk1.mux4_I\[12\].x
rlabel metal1 150328 2414 150328 2414 0 col\[4\].genblk1.mux4_I\[13\].x
rlabel metal1 150328 2958 150328 2958 0 col\[4\].genblk1.mux4_I\[14\].x
rlabel metal2 147522 3332 147522 3332 0 col\[4\].genblk1.mux4_I\[15\].x
rlabel metal2 147982 3842 147982 3842 0 col\[4\].genblk1.mux4_I\[16\].x
rlabel metal1 145314 2550 145314 2550 0 col\[4\].genblk1.mux4_I\[17\].x
rlabel metal1 144900 3638 144900 3638 0 col\[4\].genblk1.mux4_I\[18\].x
rlabel metal1 143244 3162 143244 3162 0 col\[4\].genblk1.mux4_I\[19\].x
rlabel metal1 160310 3094 160310 3094 0 col\[4\].genblk1.mux4_I\[1\].x
rlabel metal2 143106 6188 143106 6188 0 col\[4\].genblk1.mux4_I\[20\].x
rlabel metal1 141588 1734 141588 1734 0 col\[4\].genblk1.mux4_I\[21\].x
rlabel metal2 139978 2176 139978 2176 0 col\[4\].genblk1.mux4_I\[22\].x
rlabel metal1 139288 3162 139288 3162 0 col\[4\].genblk1.mux4_I\[23\].x
rlabel metal1 160632 4046 160632 4046 0 col\[4\].genblk1.mux4_I\[2\].x
rlabel metal1 157872 3094 157872 3094 0 col\[4\].genblk1.mux4_I\[3\].x
rlabel metal1 157918 3706 157918 3706 0 col\[4\].genblk1.mux4_I\[4\].x
rlabel metal1 155526 4590 155526 4590 0 col\[4\].genblk1.mux4_I\[5\].x
rlabel metal1 154146 4046 154146 4046 0 col\[4\].genblk1.mux4_I\[6\].x
rlabel metal1 152950 5338 152950 5338 0 col\[4\].genblk1.mux4_I\[7\].x
rlabel metal2 152398 4862 152398 4862 0 col\[4\].genblk1.mux4_I\[8\].x
rlabel metal2 152398 7140 152398 7140 0 col\[4\].genblk1.mux4_I\[9\].x
rlabel metal1 171120 5848 171120 5848 0 col\[4\].genblk1.tbuf_row_ena_I.t
rlabel metal1 161506 5678 161506 5678 0 col\[4\].genblk1.tbuf_row_ena_I.tx
rlabel metal1 157458 1292 157458 1292 0 col\[4\].zbuf_bot_ena_I.e
rlabel metal1 168452 1326 168452 1326 0 col\[4\].zbuf_bot_ena_I.z
rlabel metal1 168544 1938 168544 1938 0 col\[4\].zbuf_bot_iw_I\[0\].z
rlabel metal2 161506 1530 161506 1530 0 col\[4\].zbuf_bot_iw_I\[10\].z
rlabel metal1 160770 2380 160770 2380 0 col\[4\].zbuf_bot_iw_I\[11\].z
rlabel metal1 159942 1326 159942 1326 0 col\[4\].zbuf_bot_iw_I\[12\].z
rlabel metal2 160218 1530 160218 1530 0 col\[4\].zbuf_bot_iw_I\[13\].z
rlabel metal1 155158 1904 155158 1904 0 col\[4\].zbuf_bot_iw_I\[14\].z
rlabel metal1 158332 1190 158332 1190 0 col\[4\].zbuf_bot_iw_I\[15\].z
rlabel metal1 157504 1530 157504 1530 0 col\[4\].zbuf_bot_iw_I\[16\].z
rlabel metal1 156768 1530 156768 1530 0 col\[4\].zbuf_bot_iw_I\[17\].z
rlabel metal1 167624 1326 167624 1326 0 col\[4\].zbuf_bot_iw_I\[1\].z
rlabel metal2 167486 2244 167486 2244 0 col\[4\].zbuf_bot_iw_I\[2\].z
rlabel metal1 166290 2074 166290 2074 0 col\[4\].zbuf_bot_iw_I\[3\].z
rlabel metal2 165646 2244 165646 2244 0 col\[4\].zbuf_bot_iw_I\[4\].z
rlabel metal2 164542 1530 164542 1530 0 col\[4\].zbuf_bot_iw_I\[5\].z
rlabel metal1 164266 1326 164266 1326 0 col\[4\].zbuf_bot_iw_I\[6\].z
rlabel metal2 163990 2244 163990 2244 0 col\[4\].zbuf_bot_iw_I\[7\].z
rlabel metal1 162748 1326 162748 1326 0 col\[4\].zbuf_bot_iw_I\[8\].z
rlabel metal2 162334 2244 162334 2244 0 col\[4\].zbuf_bot_iw_I\[9\].z
rlabel metal1 163254 7344 163254 7344 0 col\[4\].zbuf_top_ena_I.e
rlabel metal2 169970 8772 169970 8772 0 col\[4\].zbuf_top_ena_I.z
rlabel metal2 168866 8602 168866 8602 0 col\[4\].zbuf_top_iw_I\[0\].z
rlabel metal2 161138 8364 161138 8364 0 col\[4\].zbuf_top_iw_I\[10\].z
rlabel metal2 160126 8058 160126 8058 0 col\[4\].zbuf_top_iw_I\[11\].z
rlabel metal2 159390 9078 159390 9078 0 col\[4\].zbuf_top_iw_I\[12\].z
rlabel metal1 158838 8602 158838 8602 0 col\[4\].zbuf_top_iw_I\[13\].z
rlabel metal2 157826 9350 157826 9350 0 col\[4\].zbuf_top_iw_I\[14\].z
rlabel metal2 157458 9078 157458 9078 0 col\[4\].zbuf_top_iw_I\[15\].z
rlabel metal2 156998 9350 156998 9350 0 col\[4\].zbuf_top_iw_I\[16\].z
rlabel metal2 156170 9350 156170 9350 0 col\[4\].zbuf_top_iw_I\[17\].z
rlabel metal2 167670 8330 167670 8330 0 col\[4\].zbuf_top_iw_I\[1\].z
rlabel metal2 167486 8602 167486 8602 0 col\[4\].zbuf_top_iw_I\[2\].z
rlabel metal2 166198 8602 166198 8602 0 col\[4\].zbuf_top_iw_I\[3\].z
rlabel metal2 165370 7548 165370 7548 0 col\[4\].zbuf_top_iw_I\[4\].z
rlabel metal2 164634 7548 164634 7548 0 col\[4\].zbuf_top_iw_I\[5\].z
rlabel metal2 165186 9078 165186 9078 0 col\[4\].zbuf_top_iw_I\[6\].z
rlabel metal2 163898 7548 163898 7548 0 col\[4\].zbuf_top_iw_I\[7\].z
rlabel metal2 162426 7820 162426 7820 0 col\[4\].zbuf_top_iw_I\[8\].z
rlabel metal1 162012 7854 162012 7854 0 col\[4\].zbuf_top_iw_I\[9\].z
rlabel metal2 190946 3026 190946 3026 0 col\[5\].zbuf_bot_ena_I.e
rlabel metal1 202952 1326 202952 1326 0 col\[5\].zbuf_bot_ena_I.z
rlabel metal1 202584 2414 202584 2414 0 col\[5\].zbuf_bot_iw_I\[0\].z
rlabel metal1 196098 1326 196098 1326 0 col\[5\].zbuf_bot_iw_I\[10\].z
rlabel metal2 195730 2244 195730 2244 0 col\[5\].zbuf_bot_iw_I\[11\].z
rlabel metal2 194626 1530 194626 1530 0 col\[5\].zbuf_bot_iw_I\[12\].z
rlabel metal2 193338 1530 193338 1530 0 col\[5\].zbuf_bot_iw_I\[13\].z
rlabel metal1 192878 1326 192878 1326 0 col\[5\].zbuf_bot_iw_I\[14\].z
rlabel metal2 192418 2244 192418 2244 0 col\[5\].zbuf_bot_iw_I\[15\].z
rlabel metal2 191406 1938 191406 1938 0 col\[5\].zbuf_bot_iw_I\[16\].z
rlabel metal2 190394 2244 190394 2244 0 col\[5\].zbuf_bot_iw_I\[17\].z
rlabel metal1 202952 1938 202952 1938 0 col\[5\].zbuf_bot_iw_I\[1\].z
rlabel metal1 201434 1190 201434 1190 0 col\[5\].zbuf_bot_iw_I\[2\].z
rlabel metal1 200514 1292 200514 1292 0 col\[5\].zbuf_bot_iw_I\[3\].z
rlabel metal2 200882 2244 200882 2244 0 col\[5\].zbuf_bot_iw_I\[4\].z
rlabel metal2 199778 1530 199778 1530 0 col\[5\].zbuf_bot_iw_I\[5\].z
rlabel metal2 199226 2244 199226 2244 0 col\[5\].zbuf_bot_iw_I\[6\].z
rlabel metal2 197938 1530 197938 1530 0 col\[5\].zbuf_bot_iw_I\[7\].z
rlabel metal1 197340 1326 197340 1326 0 col\[5\].zbuf_bot_iw_I\[8\].z
rlabel metal1 196926 2074 196926 2074 0 col\[5\].zbuf_bot_iw_I\[9\].z
rlabel metal2 190854 9282 190854 9282 0 col\[5\].zbuf_top_ena_I.e
rlabel metal2 203550 8772 203550 8772 0 col\[5\].zbuf_top_ena_I.z
rlabel metal2 203458 9248 203458 9248 0 col\[5\].zbuf_top_iw_I\[0\].z
rlabel metal2 196374 8636 196374 8636 0 col\[5\].zbuf_top_iw_I\[10\].z
rlabel metal2 195822 9350 195822 9350 0 col\[5\].zbuf_top_iw_I\[11\].z
rlabel metal2 194074 8636 194074 8636 0 col\[5\].zbuf_top_iw_I\[12\].z
rlabel metal2 193614 9078 193614 9078 0 col\[5\].zbuf_top_iw_I\[13\].z
rlabel metal1 193016 9146 193016 9146 0 col\[5\].zbuf_top_iw_I\[14\].z
rlabel metal2 192050 8636 192050 8636 0 col\[5\].zbuf_top_iw_I\[15\].z
rlabel metal1 191544 8466 191544 8466 0 col\[5\].zbuf_top_iw_I\[16\].z
rlabel metal2 190394 8636 190394 8636 0 col\[5\].zbuf_top_iw_I\[17\].z
rlabel metal2 202722 9078 202722 9078 0 col\[5\].zbuf_top_iw_I\[1\].z
rlabel metal1 201940 8466 201940 8466 0 col\[5\].zbuf_top_iw_I\[2\].z
rlabel metal1 200882 8466 200882 8466 0 col\[5\].zbuf_top_iw_I\[3\].z
rlabel metal1 200422 9146 200422 9146 0 col\[5\].zbuf_top_iw_I\[4\].z
rlabel metal2 199318 8636 199318 8636 0 col\[5\].zbuf_top_iw_I\[5\].z
rlabel metal2 198858 9078 198858 9078 0 col\[5\].zbuf_top_iw_I\[6\].z
rlabel metal1 198444 9146 198444 9146 0 col\[5\].zbuf_top_iw_I\[7\].z
rlabel metal2 197570 9078 197570 9078 0 col\[5\].zbuf_top_iw_I\[8\].z
rlabel metal2 196650 9078 196650 9078 0 col\[5\].zbuf_top_iw_I\[9\].z
rlabel metal2 227378 3876 227378 3876 0 col\[6\].genblk1.mux4_I\[0\].x
rlabel metal1 214222 6324 214222 6324 0 col\[6\].genblk1.mux4_I\[10\].x
rlabel viali 212842 5754 212842 5754 0 col\[6\].genblk1.mux4_I\[11\].x
rlabel metal1 213256 6834 213256 6834 0 col\[6\].genblk1.mux4_I\[12\].x
rlabel metal2 217258 3332 217258 3332 0 col\[6\].genblk1.mux4_I\[13\].x
rlabel metal2 214038 4964 214038 4964 0 col\[6\].genblk1.mux4_I\[14\].x
rlabel metal2 215142 4352 215142 4352 0 col\[6\].genblk1.mux4_I\[15\].x
rlabel metal1 210542 3638 210542 3638 0 col\[6\].genblk1.mux4_I\[16\].x
rlabel metal1 209806 4148 209806 4148 0 col\[6\].genblk1.mux4_I\[17\].x
rlabel metal1 212382 3366 212382 3366 0 col\[6\].genblk1.mux4_I\[18\].x
rlabel metal2 214498 3451 214498 3451 0 col\[6\].genblk1.mux4_I\[19\].x
rlabel metal2 226182 4352 226182 4352 0 col\[6\].genblk1.mux4_I\[1\].x
rlabel metal2 212106 6494 212106 6494 0 col\[6\].genblk1.mux4_I\[20\].x
rlabel metal1 204930 2550 204930 2550 0 col\[6\].genblk1.mux4_I\[21\].x
rlabel metal2 204930 3332 204930 3332 0 col\[6\].genblk1.mux4_I\[22\].x
rlabel metal1 204286 2890 204286 2890 0 col\[6\].genblk1.mux4_I\[23\].x
rlabel metal1 225722 5236 225722 5236 0 col\[6\].genblk1.mux4_I\[2\].x
rlabel metal2 225538 7038 225538 7038 0 col\[6\].genblk1.mux4_I\[3\].x
rlabel metal2 223698 6460 223698 6460 0 col\[6\].genblk1.mux4_I\[4\].x
rlabel metal1 222640 5202 222640 5202 0 col\[6\].genblk1.mux4_I\[5\].x
rlabel metal1 221950 5746 221950 5746 0 col\[6\].genblk1.mux4_I\[6\].x
rlabel metal2 220662 5372 220662 5372 0 col\[6\].genblk1.mux4_I\[7\].x
rlabel via1 219282 5219 219282 5219 0 col\[6\].genblk1.mux4_I\[8\].x
rlabel metal1 216890 6834 216890 6834 0 col\[6\].genblk1.mux4_I\[9\].x
rlabel metal2 230046 5440 230046 5440 0 col\[6\].genblk1.tbuf_row_ena_I.t
rlabel metal1 228482 5236 228482 5236 0 col\[6\].genblk1.tbuf_row_ena_I.tx
rlabel metal1 236348 1938 236348 1938 0 col\[6\].zbuf_bot_ena_I.e
rlabel metal1 237176 1938 237176 1938 0 col\[6\].zbuf_bot_ena_I.z
rlabel metal1 236394 1530 236394 1530 0 col\[6\].zbuf_bot_iw_I\[0\].z
rlabel metal1 229126 1326 229126 1326 0 col\[6\].zbuf_bot_iw_I\[10\].z
rlabel metal1 228666 1530 228666 1530 0 col\[6\].zbuf_bot_iw_I\[11\].z
rlabel metal1 228298 2074 228298 2074 0 col\[6\].zbuf_bot_iw_I\[12\].z
rlabel metal1 227010 3026 227010 3026 0 col\[6\].zbuf_bot_iw_I\[13\].z
rlabel metal2 227010 2244 227010 2244 0 col\[6\].zbuf_bot_iw_I\[14\].z
rlabel metal1 226090 1530 226090 1530 0 col\[6\].zbuf_bot_iw_I\[15\].z
rlabel metal2 226182 2244 226182 2244 0 col\[6\].zbuf_bot_iw_I\[16\].z
rlabel metal2 225354 2244 225354 2244 0 col\[6\].zbuf_bot_iw_I\[17\].z
rlabel metal2 236118 2244 236118 2244 0 col\[6\].zbuf_bot_iw_I\[1\].z
rlabel metal2 234738 1530 234738 1530 0 col\[6\].zbuf_bot_iw_I\[2\].z
rlabel metal2 234002 1530 234002 1530 0 col\[6\].zbuf_bot_iw_I\[3\].z
rlabel metal2 233266 1530 233266 1530 0 col\[6\].zbuf_bot_iw_I\[4\].z
rlabel metal1 232576 1530 232576 1530 0 col\[6\].zbuf_bot_iw_I\[5\].z
rlabel metal1 232254 2006 232254 2006 0 col\[6\].zbuf_bot_iw_I\[6\].z
rlabel metal2 231794 2210 231794 2210 0 col\[6\].zbuf_bot_iw_I\[7\].z
rlabel metal2 230690 1530 230690 1530 0 col\[6\].zbuf_bot_iw_I\[8\].z
rlabel metal2 229678 1530 229678 1530 0 col\[6\].zbuf_bot_iw_I\[9\].z
rlabel metal1 230506 8942 230506 8942 0 col\[6\].zbuf_top_ena_I.e
rlabel metal1 236072 8602 236072 8602 0 col\[6\].zbuf_top_ena_I.z
rlabel metal1 236348 8466 236348 8466 0 col\[6\].zbuf_top_iw_I\[0\].z
rlabel metal2 228942 8636 228942 8636 0 col\[6\].zbuf_top_iw_I\[10\].z
rlabel metal2 228390 9350 228390 9350 0 col\[6\].zbuf_top_iw_I\[11\].z
rlabel metal2 228114 8636 228114 8636 0 col\[6\].zbuf_top_iw_I\[12\].z
rlabel metal2 226550 8636 226550 8636 0 col\[6\].zbuf_top_iw_I\[13\].z
rlabel metal2 225814 8636 225814 8636 0 col\[6\].zbuf_top_iw_I\[14\].z
rlabel metal1 225262 9554 225262 9554 0 col\[6\].zbuf_top_iw_I\[15\].z
rlabel metal1 224848 8466 224848 8466 0 col\[6\].zbuf_top_iw_I\[16\].z
rlabel metal1 223238 8976 223238 8976 0 col\[6\].zbuf_top_iw_I\[17\].z
rlabel viali 236670 8939 236670 8939 0 col\[6\].zbuf_top_iw_I\[1\].z
rlabel metal2 234922 9078 234922 9078 0 col\[6\].zbuf_top_iw_I\[2\].z
rlabel metal2 234186 9350 234186 9350 0 col\[6\].zbuf_top_iw_I\[3\].z
rlabel metal2 234094 9350 234094 9350 0 col\[6\].zbuf_top_iw_I\[4\].z
rlabel metal2 233266 8636 233266 8636 0 col\[6\].zbuf_top_iw_I\[5\].z
rlabel metal2 231794 8636 231794 8636 0 col\[6\].zbuf_top_iw_I\[6\].z
rlabel metal2 231058 9078 231058 9078 0 col\[6\].zbuf_top_iw_I\[7\].z
rlabel metal1 230644 7854 230644 7854 0 col\[6\].zbuf_top_iw_I\[8\].z
rlabel metal2 230046 9282 230046 9282 0 col\[6\].zbuf_top_iw_I\[9\].z
rlabel metal1 264224 2414 264224 2414 0 col\[7\].zbuf_bot_ena_I.e
rlabel metal2 270526 2244 270526 2244 0 col\[7\].zbuf_bot_ena_I.z
rlabel metal1 269790 1326 269790 1326 0 col\[7\].zbuf_bot_iw_I\[0\].z
rlabel metal2 263074 1530 263074 1530 0 col\[7\].zbuf_bot_iw_I\[10\].z
rlabel metal2 262338 1530 262338 1530 0 col\[7\].zbuf_bot_iw_I\[11\].z
rlabel metal1 261740 2074 261740 2074 0 col\[7\].zbuf_bot_iw_I\[12\].z
rlabel metal2 261602 1530 261602 1530 0 col\[7\].zbuf_bot_iw_I\[13\].z
rlabel metal2 260314 1530 260314 1530 0 col\[7\].zbuf_bot_iw_I\[14\].z
rlabel metal1 259532 2414 259532 2414 0 col\[7\].zbuf_bot_iw_I\[15\].z
rlabel metal1 259210 2074 259210 2074 0 col\[7\].zbuf_bot_iw_I\[16\].z
rlabel metal1 258060 1326 258060 1326 0 col\[7\].zbuf_bot_iw_I\[17\].z
rlabel metal1 270066 1326 270066 1326 0 col\[7\].zbuf_bot_iw_I\[1\].z
rlabel metal2 269698 2244 269698 2244 0 col\[7\].zbuf_bot_iw_I\[2\].z
rlabel metal2 268226 1530 268226 1530 0 col\[7\].zbuf_bot_iw_I\[3\].z
rlabel metal2 267858 1530 267858 1530 0 col\[7\].zbuf_bot_iw_I\[4\].z
rlabel metal2 266754 1530 266754 1530 0 col\[7\].zbuf_bot_iw_I\[5\].z
rlabel metal2 265926 1530 265926 1530 0 col\[7\].zbuf_bot_iw_I\[6\].z
rlabel metal2 265190 1530 265190 1530 0 col\[7\].zbuf_bot_iw_I\[7\].z
rlabel metal1 264592 2414 264592 2414 0 col\[7\].zbuf_bot_iw_I\[8\].z
rlabel metal2 264178 1530 264178 1530 0 col\[7\].zbuf_bot_iw_I\[9\].z
rlabel metal2 235290 7871 235290 7871 0 col\[7\].zbuf_top_ena_I.e
rlabel viali 269885 3502 269885 3502 0 col\[7\].zbuf_top_ena_I.z
rlabel metal1 270388 4114 270388 4114 0 col\[7\].zbuf_top_iw_I\[0\].z
rlabel metal2 263074 7548 263074 7548 0 col\[7\].zbuf_top_iw_I\[10\].z
rlabel metal2 262338 7548 262338 7548 0 col\[7\].zbuf_top_iw_I\[11\].z
rlabel metal2 261602 8364 261602 8364 0 col\[7\].zbuf_top_iw_I\[12\].z
rlabel metal1 262246 9588 262246 9588 0 col\[7\].zbuf_top_iw_I\[13\].z
rlabel metal2 260314 8058 260314 8058 0 col\[7\].zbuf_top_iw_I\[14\].z
rlabel metal1 259624 9554 259624 9554 0 col\[7\].zbuf_top_iw_I\[15\].z
rlabel metal2 258842 8058 258842 8058 0 col\[7\].zbuf_top_iw_I\[16\].z
rlabel metal2 258106 8908 258106 8908 0 col\[7\].zbuf_top_iw_I\[17\].z
rlabel metal1 269008 3502 269008 3502 0 col\[7\].zbuf_top_iw_I\[1\].z
rlabel metal1 269514 4114 269514 4114 0 col\[7\].zbuf_top_iw_I\[2\].z
rlabel metal2 267674 5644 267674 5644 0 col\[7\].zbuf_top_iw_I\[3\].z
rlabel metal1 267536 5202 267536 5202 0 col\[7\].zbuf_top_iw_I\[4\].z
rlabel metal1 266432 4590 266432 4590 0 col\[7\].zbuf_top_iw_I\[5\].z
rlabel metal2 265650 7888 265650 7888 0 col\[7\].zbuf_top_iw_I\[6\].z
rlabel metal2 265558 8058 265558 8058 0 col\[7\].zbuf_top_iw_I\[7\].z
rlabel metal2 264086 8058 264086 8058 0 col\[7\].zbuf_top_iw_I\[8\].z
rlabel metal2 264178 7548 264178 7548 0 col\[7\].zbuf_top_iw_I\[9\].z
rlabel metal1 267260 8466 267260 8466 0 net1
rlabel metal1 268962 3162 268962 3162 0 net10
rlabel metal2 109894 1088 109894 1088 0 net100
rlabel metal2 37490 3145 37490 3145 0 net101
rlabel metal2 108882 1088 108882 1088 0 net102
rlabel metal1 107962 1190 107962 1190 0 net103
rlabel metal1 106950 1190 106950 1190 0 net104
rlabel metal1 105386 1802 105386 1802 0 net105
rlabel metal1 106214 1224 106214 1224 0 net106
rlabel metal2 105478 1513 105478 1513 0 net107
rlabel metal1 104696 1190 104696 1190 0 net108
rlabel metal1 103730 1224 103730 1224 0 net109
rlabel metal1 270802 2924 270802 2924 0 net11
rlabel metal2 121026 7276 121026 7276 0 net110
rlabel metal2 120106 4403 120106 4403 0 net111
rlabel metal1 36524 4658 36524 4658 0 net112
rlabel metal2 119186 6970 119186 6970 0 net113
rlabel via1 118367 5134 118367 5134 0 net114
rlabel metal1 115782 3570 115782 3570 0 net115
rlabel metal2 115598 6460 115598 6460 0 net116
rlabel metal1 113206 4046 113206 4046 0 net117
rlabel metal1 112654 5134 112654 5134 0 net118
rlabel metal2 110722 4998 110722 4998 0 net119
rlabel metal1 269008 3706 269008 3706 0 net12
rlabel metal2 110538 7548 110538 7548 0 net120
rlabel metal2 109066 6698 109066 6698 0 net121
rlabel metal2 112746 9248 112746 9248 0 net122
rlabel metal2 9430 816 9430 816 0 net123
rlabel metal1 105800 7922 105800 7922 0 net124
rlabel metal1 108054 4046 108054 4046 0 net125
rlabel metal2 110630 7242 110630 7242 0 net126
rlabel metal2 109894 9078 109894 9078 0 net127
rlabel metal2 105846 4267 105846 4267 0 net128
rlabel metal1 106306 9010 106306 9010 0 net129
rlabel metal1 268962 3366 268962 3366 0 net13
rlabel viali 102635 3026 102635 3026 0 net130
rlabel metal1 100510 2958 100510 2958 0 net131
rlabel metal2 100372 6834 100372 6834 0 net132
rlabel metal1 97520 2958 97520 2958 0 net133
rlabel metal2 5474 884 5474 884 0 net134
rlabel metal2 97658 2533 97658 2533 0 net135
rlabel metal2 97566 6868 97566 6868 0 net136
rlabel metal1 155112 2550 155112 2550 0 net137
rlabel metal1 155388 1190 155388 1190 0 net138
rlabel metal1 154054 1224 154054 1224 0 net139
rlabel metal2 267030 5372 267030 5372 0 net14
rlabel metal1 153686 1190 153686 1190 0 net140
rlabel metal2 152122 1054 152122 1054 0 net141
rlabel metal1 151478 1224 151478 1224 0 net142
rlabel metal1 150880 1190 150880 1190 0 net143
rlabel metal1 150374 2074 150374 2074 0 net144
rlabel metal2 4830 2244 4830 2244 0 net145
rlabel metal2 17986 850 17986 850 0 net146
rlabel metal1 150144 1190 150144 1190 0 net147
rlabel metal1 148902 1224 148902 1224 0 net148
rlabel metal2 148258 1975 148258 1975 0 net149
rlabel metal1 268548 2890 268548 2890 0 net15
rlabel metal1 146694 1190 146694 1190 0 net150
rlabel metal1 146234 1190 146234 1190 0 net151
rlabel metal2 147798 1666 147798 1666 0 net152
rlabel metal2 148166 2380 148166 2380 0 net153
rlabel metal1 144486 2958 144486 2958 0 net154
rlabel metal1 143796 1190 143796 1190 0 net155
rlabel metal2 142830 2108 142830 2108 0 net156
rlabel metal2 4186 986 4186 986 0 net157
rlabel metal2 143152 3094 143152 3094 0 net158
rlabel metal1 141864 1190 141864 1190 0 net159
rlabel metal2 239154 6902 239154 6902 0 net16
rlabel metal1 141036 1190 141036 1190 0 net160
rlabel metal1 140622 1462 140622 1462 0 net161
rlabel metal1 138782 1462 138782 1462 0 net162
rlabel metal2 137954 2074 137954 2074 0 net163
rlabel metal2 158378 6324 158378 6324 0 net164
rlabel metal1 155802 9520 155802 9520 0 net165
rlabel metal1 155710 9452 155710 9452 0 net166
rlabel metal2 155986 6307 155986 6307 0 net167
rlabel metal2 2898 850 2898 850 0 net168
rlabel metal1 155158 3570 155158 3570 0 net169
rlabel metal1 267812 3706 267812 3706 0 net17
rlabel metal1 152582 4658 152582 4658 0 net170
rlabel metal1 151524 4046 151524 4046 0 net171
rlabel metal1 150282 5202 150282 5202 0 net172
rlabel metal1 150512 4658 150512 4658 0 net173
rlabel metal2 150558 8126 150558 8126 0 net174
rlabel metal2 148258 8092 148258 8092 0 net175
rlabel metal2 145866 8126 145866 8126 0 net176
rlabel metal1 145682 7446 145682 7446 0 net177
rlabel metal1 147246 2482 147246 2482 0 net178
rlabel metal2 2622 2142 2622 2142 0 net179
rlabel metal2 266386 4726 266386 4726 0 net18
rlabel metal2 147798 5916 147798 5916 0 net180
rlabel metal1 145636 2958 145636 2958 0 net181
rlabel metal2 145406 6494 145406 6494 0 net182
rlabel metal1 143152 2482 143152 2482 0 net183
rlabel metal1 143060 3570 143060 3570 0 net184
rlabel metal1 142784 2958 142784 2958 0 net185
rlabel metal1 140622 6834 140622 6834 0 net186
rlabel metal1 140484 1938 140484 1938 0 net187
rlabel metal1 138690 9350 138690 9350 0 net188
rlabel metal2 137770 6188 137770 6188 0 net189
rlabel metal2 265190 4964 265190 4964 0 net19
rlabel metal2 36662 2244 36662 2244 0 net190
rlabel metal1 187082 2482 187082 2482 0 net191
rlabel metal2 189750 1088 189750 1088 0 net192
rlabel metal1 161046 2618 161046 2618 0 net193
rlabel metal1 187266 2550 187266 2550 0 net194
rlabel metal2 167578 2210 167578 2210 0 net195
rlabel metal1 161460 442 161460 442 0 net196
rlabel metal2 185058 2091 185058 2091 0 net197
rlabel metal3 182620 1088 182620 1088 0 net198
rlabel metal2 173834 3349 173834 3349 0 net199
rlabel metal1 264638 3910 264638 3910 0 net2
rlabel metal1 268318 2278 268318 2278 0 net20
rlabel metal2 182850 1122 182850 1122 0 net200
rlabel metal2 52854 6188 52854 6188 0 net201
rlabel metal3 166060 1904 166060 1904 0 net202
rlabel metal2 171442 1020 171442 1020 0 net203
rlabel metal2 146786 7446 146786 7446 0 net204
rlabel metal1 153318 2516 153318 2516 0 net205
rlabel metal1 179446 1972 179446 1972 0 net206
rlabel metal2 179446 1020 179446 1020 0 net207
rlabel metal1 178158 1836 178158 1836 0 net208
rlabel metal2 176962 1938 176962 1938 0 net209
rlabel metal1 267306 2924 267306 2924 0 net21
rlabel metal2 176870 2023 176870 2023 0 net210
rlabel metal2 176870 986 176870 986 0 net211
rlabel metal2 20378 8432 20378 8432 0 net212
rlabel metal2 174754 2142 174754 2142 0 net213
rlabel metal2 174294 1156 174294 1156 0 net214
rlabel metal2 173282 2159 173282 2159 0 net215
rlabel metal2 172546 952 172546 952 0 net216
rlabel metal1 168958 7888 168958 7888 0 net217
rlabel metal1 174662 9520 174662 9520 0 net218
rlabel metal2 170614 9384 170614 9384 0 net219
rlabel metal1 267766 2312 267766 2312 0 net22
rlabel metal2 187082 9180 187082 9180 0 net220
rlabel metal1 171120 6324 171120 6324 0 net221
rlabel metal1 187174 9418 187174 9418 0 net222
rlabel metal2 17342 9792 17342 9792 0 net223
rlabel metal2 170062 8466 170062 8466 0 net224
rlabel metal1 151478 5134 151478 5134 0 net225
rlabel metal2 173466 8211 173466 8211 0 net226
rlabel metal2 151478 7276 151478 7276 0 net227
rlabel metal2 149178 7344 149178 7344 0 net228
rlabel metal2 151754 9316 151754 9316 0 net229
rlabel metal2 266662 3944 266662 3944 0 net23
rlabel metal1 152582 7310 152582 7310 0 net230
rlabel via2 149178 2499 149178 2499 0 net231
rlabel metal2 148902 3230 148902 3230 0 net232
rlabel metal2 146602 5355 146602 5355 0 net233
rlabel metal2 51106 7684 51106 7684 0 net234
rlabel metal2 146326 4437 146326 4437 0 net235
rlabel metal1 144256 2482 144256 2482 0 net236
rlabel metal2 144026 5644 144026 5644 0 net237
rlabel metal2 175950 7344 175950 7344 0 net238
rlabel metal2 174754 8636 174754 8636 0 net239
rlabel metal2 266018 4454 266018 4454 0 net24
rlabel metal2 174202 6069 174202 6069 0 net240
rlabel metal2 173190 6528 173190 6528 0 net241
rlabel metal2 172546 9962 172546 9962 0 net242
rlabel metal2 225722 3332 225722 3332 0 net243
rlabel metal1 223560 3706 223560 3706 0 net244
rlabel metal2 15594 7922 15594 7922 0 net245
rlabel metal1 225400 5678 225400 5678 0 net246
rlabel metal1 223054 1190 223054 1190 0 net247
rlabel metal1 222870 6732 222870 6732 0 net248
rlabel metal1 221168 1530 221168 1530 0 net249
rlabel metal1 265466 4250 265466 4250 0 net25
rlabel metal1 220984 1190 220984 1190 0 net250
rlabel metal1 220432 6222 220432 6222 0 net251
rlabel metal2 219650 1088 219650 1088 0 net252
rlabel metal1 216568 2074 216568 2074 0 net253
rlabel metal1 216522 1224 216522 1224 0 net254
rlabel metal1 215740 1190 215740 1190 0 net255
rlabel metal1 18469 9486 18469 9486 0 net256
rlabel metal2 17250 1020 17250 1020 0 net257
rlabel metal2 215142 7412 215142 7412 0 net258
rlabel metal1 214176 1190 214176 1190 0 net259
rlabel metal1 267766 2618 267766 2618 0 net26
rlabel metal1 213302 1360 213302 1360 0 net260
rlabel metal1 214682 4046 214682 4046 0 net261
rlabel metal1 213486 2074 213486 2074 0 net262
rlabel metal1 212428 4046 212428 4046 0 net263
rlabel metal1 212612 3502 212612 3502 0 net264
rlabel metal1 210220 1190 210220 1190 0 net265
rlabel metal1 210174 6766 210174 6766 0 net266
rlabel metal1 208150 1224 208150 1224 0 net267
rlabel metal2 13754 7888 13754 7888 0 net268
rlabel metal2 207506 1088 207506 1088 0 net269
rlabel metal2 270434 9826 270434 9826 0 net27
rlabel metal1 207184 2958 207184 2958 0 net270
rlabel metal2 225170 6460 225170 6460 0 net271
rlabel metal1 223652 4046 223652 4046 0 net272
rlabel metal1 225239 5746 225239 5746 0 net273
rlabel metal1 222916 7378 222916 7378 0 net274
rlabel metal1 222410 6834 222410 6834 0 net275
rlabel metal1 220478 7378 220478 7378 0 net276
rlabel metal1 219788 6834 219788 6834 0 net277
rlabel metal1 219742 6222 219742 6222 0 net278
rlabel metal2 13570 8568 13570 8568 0 net279
rlabel via2 267766 7259 267766 7259 0 net28
rlabel metal2 217810 7820 217810 7820 0 net280
rlabel metal1 217258 7378 217258 7378 0 net281
rlabel metal1 217856 6766 217856 6766 0 net282
rlabel metal2 215418 7548 215418 7548 0 net283
rlabel metal2 214498 8364 214498 8364 0 net284
rlabel metal2 213946 9146 213946 9146 0 net285
rlabel metal1 214268 4658 214268 4658 0 net286
rlabel metal1 213808 9622 213808 9622 0 net287
rlabel metal1 214820 3570 214820 3570 0 net288
rlabel metal1 212750 4114 212750 4114 0 net289
rlabel metal2 263718 8160 263718 8160 0 net29
rlabel metal2 12834 9214 12834 9214 0 net290
rlabel metal1 211876 3570 211876 3570 0 net291
rlabel metal1 212428 3026 212428 3026 0 net292
rlabel metal1 209530 6834 209530 6834 0 net293
rlabel metal1 209116 2482 209116 2482 0 net294
rlabel metal1 209852 2958 209852 2958 0 net295
rlabel metal1 207598 3026 207598 3026 0 net296
rlabel metal1 248446 1292 248446 1292 0 net297
rlabel metal1 234002 1836 234002 1836 0 net298
rlabel metal2 252494 4896 252494 4896 0 net299
rlabel metal2 268226 6052 268226 6052 0 net3
rlabel via2 237038 7837 237038 7837 0 net30
rlabel metal1 234600 408 234600 408 0 net300
rlabel metal2 14766 8704 14766 8704 0 net301
rlabel metal2 244306 3485 244306 3485 0 net302
rlabel metal2 254058 1326 254058 1326 0 net303
rlabel metal2 229770 578 229770 578 0 net304
rlabel metal2 252586 4131 252586 4131 0 net305
rlabel metal2 251850 816 251850 816 0 net306
rlabel metal2 251482 2754 251482 2754 0 net307
rlabel metal2 250286 1020 250286 1020 0 net308
rlabel metal1 238096 1938 238096 1938 0 net309
rlabel metal2 259946 3145 259946 3145 0 net31
rlabel metal2 248078 1037 248078 1037 0 net310
rlabel metal2 248998 2686 248998 2686 0 net311
rlabel metal2 11362 7208 11362 7208 0 net312
rlabel metal2 248998 952 248998 952 0 net313
rlabel metal1 223790 2380 223790 2380 0 net314
rlabel metal1 246422 1836 246422 1836 0 net315
rlabel via1 213866 4046 213866 4046 0 net316
rlabel via1 213498 3502 213498 3502 0 net317
rlabel metal1 221766 2516 221766 2516 0 net318
rlabel via1 211347 6766 211347 6766 0 net319
rlabel metal2 268778 7871 268778 7871 0 net32
rlabel metal2 211094 1462 211094 1462 0 net320
rlabel via1 211106 3026 211106 3026 0 net321
rlabel via1 208863 2958 208863 2958 0 net322
rlabel metal2 17250 7514 17250 7514 0 net323
rlabel metal1 227424 1530 227424 1530 0 net324
rlabel metal2 225262 3876 225262 3876 0 net325
rlabel metal1 227562 5746 227562 5746 0 net326
rlabel metal1 248400 7276 248400 7276 0 net327
rlabel metal2 225630 6307 225630 6307 0 net328
rlabel metal2 221490 7446 221490 7446 0 net329
rlabel metal1 266570 9010 266570 9010 0 net33
rlabel metal1 226642 7956 226642 7956 0 net330
rlabel metal2 252862 7548 252862 7548 0 net331
rlabel metal2 251850 7089 251850 7089 0 net332
rlabel metal2 251390 8194 251390 8194 0 net333
rlabel metal2 9982 7888 9982 7888 0 net334
rlabel metal1 251528 9486 251528 9486 0 net335
rlabel metal2 249642 7293 249642 7293 0 net336
rlabel metal1 248998 8908 248998 8908 0 net337
rlabel metal2 248998 8381 248998 8381 0 net338
rlabel metal1 247112 8874 247112 8874 0 net339
rlabel metal1 266248 7922 266248 7922 0 net34
rlabel metal2 246698 8942 246698 8942 0 net340
rlabel metal1 246330 8942 246330 8942 0 net341
rlabel metal1 214590 3944 214590 3944 0 net342
rlabel metal2 213946 3043 213946 3043 0 net343
rlabel metal2 213578 3179 213578 3179 0 net344
rlabel metal2 8510 9792 8510 9792 0 net345
rlabel metal2 211186 6341 211186 6341 0 net346
rlabel metal1 211462 2482 211462 2482 0 net347
rlabel metal2 211002 3111 211002 3111 0 net348
rlabel metal2 208702 3315 208702 3315 0 net349
rlabel metal2 18722 1054 18722 1054 0 net35
rlabel metal2 8510 6664 8510 6664 0 net350
rlabel metal2 7682 9894 7682 9894 0 net351
rlabel metal2 17158 3502 17158 3502 0 net352
rlabel metal2 6946 8976 6946 8976 0 net353
rlabel metal2 5934 9860 5934 9860 0 net354
rlabel metal1 13662 9384 13662 9384 0 net355
rlabel metal1 5727 9554 5727 9554 0 net356
rlabel metal2 3450 8840 3450 8840 0 net357
rlabel metal1 36754 2346 36754 2346 0 net358
rlabel metal2 2530 9180 2530 9180 0 net359
rlabel metal2 82662 1360 82662 1360 0 net36
rlabel metal1 36340 2006 36340 2006 0 net360
rlabel metal1 52118 1190 52118 1190 0 net361
rlabel metal2 51566 2686 51566 2686 0 net362
rlabel via2 15870 1955 15870 1955 0 net363
rlabel metal1 50830 1190 50830 1190 0 net364
rlabel metal1 50508 1802 50508 1802 0 net365
rlabel metal2 49634 1975 49634 1975 0 net366
rlabel metal1 48944 1190 48944 1190 0 net367
rlabel metal1 48254 1224 48254 1224 0 net368
rlabel metal1 46966 1190 46966 1190 0 net369
rlabel metal2 82386 1666 82386 1666 0 net37
rlabel metal1 46138 1190 46138 1190 0 net370
rlabel metal1 45402 1190 45402 1190 0 net371
rlabel metal1 44942 1802 44942 1802 0 net372
rlabel metal1 43930 1462 43930 1462 0 net373
rlabel metal1 17250 3570 17250 3570 0 net374
rlabel metal1 43838 1224 43838 1224 0 net375
rlabel metal1 43056 4454 43056 4454 0 net376
rlabel metal1 41722 1190 41722 1190 0 net377
rlabel metal2 41262 2278 41262 2278 0 net378
rlabel metal2 40618 2686 40618 2686 0 net379
rlabel via2 82386 3043 82386 3043 0 net38
rlabel metal1 39606 1190 39606 1190 0 net380
rlabel metal2 38686 1734 38686 1734 0 net381
rlabel metal1 37950 3094 37950 3094 0 net382
rlabel metal1 37904 1802 37904 1802 0 net383
rlabel metal2 36754 1870 36754 1870 0 net384
rlabel metal2 14398 2992 14398 2992 0 net385
rlabel metal1 36294 3366 36294 3366 0 net386
rlabel metal1 35512 1530 35512 1530 0 net387
rlabel viali 52392 4590 52392 4590 0 net388
rlabel metal2 51290 6732 51290 6732 0 net389
rlabel metal2 81466 1326 81466 1326 0 net39
rlabel metal2 51198 7310 51198 7310 0 net390
rlabel metal1 50646 5678 50646 5678 0 net391
rlabel metal2 49266 6766 49266 6766 0 net392
rlabel metal2 47794 7004 47794 7004 0 net393
rlabel metal2 47058 3434 47058 3434 0 net394
rlabel metal2 46874 7514 46874 7514 0 net395
rlabel metal2 13570 1088 13570 1088 0 net396
rlabel metal2 46138 7310 46138 7310 0 net397
rlabel metal1 45448 6358 45448 6358 0 net398
rlabel metal1 43516 5678 43516 5678 0 net399
rlabel metal2 267766 9622 267766 9622 0 net4
rlabel metal1 80178 1258 80178 1258 0 net40
rlabel metal1 43608 5270 43608 5270 0 net400
rlabel metal1 43240 6358 43240 6358 0 net401
rlabel metal2 43286 6970 43286 6970 0 net402
rlabel metal2 41262 6834 41262 6834 0 net403
rlabel metal2 41538 3383 41538 3383 0 net404
rlabel metal2 40894 6732 40894 6732 0 net405
rlabel metal2 40158 5950 40158 5950 0 net406
rlabel metal2 12834 952 12834 952 0 net407
rlabel metal2 39330 5678 39330 5678 0 net408
rlabel metal2 38134 6222 38134 6222 0 net409
rlabel metal2 80178 4556 80178 4556 0 net41
rlabel metal2 37950 7310 37950 7310 0 net410
rlabel metal1 37168 2346 37168 2346 0 net411
rlabel metal1 36708 3502 36708 3502 0 net412
rlabel metal1 35650 9350 35650 9350 0 net413
rlabel metal2 87078 765 87078 765 0 net414
rlabel metal2 86434 2023 86434 2023 0 net415
rlabel metal3 87492 1088 87492 1088 0 net416
rlabel metal2 82754 969 82754 969 0 net417
rlabel metal2 12190 3060 12190 3060 0 net418
rlabel metal1 260406 8466 260406 8466 0 net419
rlabel metal2 80086 6069 80086 6069 0 net42
rlabel metal2 269514 9010 269514 9010 0 net420
rlabel metal2 229862 9146 229862 9146 0 net421
rlabel metal1 233910 8976 233910 8976 0 net422
rlabel metal1 195638 8908 195638 8908 0 net423
rlabel metal1 197478 8942 197478 8942 0 net424
rlabel metal1 162610 8466 162610 8466 0 net425
rlabel metal1 167716 9554 167716 9554 0 net426
rlabel metal1 128570 8908 128570 8908 0 net427
rlabel metal1 133262 8976 133262 8976 0 net428
rlabel metal2 89194 9248 89194 9248 0 net429
rlabel metal2 77602 1105 77602 1105 0 net43
rlabel metal1 98670 8908 98670 8908 0 net430
rlabel metal2 59846 8772 59846 8772 0 net431
rlabel metal2 60950 8704 60950 8704 0 net432
rlabel metal1 23460 8942 23460 8942 0 net433
rlabel metal2 32522 8636 32522 8636 0 net434
rlabel metal1 213348 6698 213348 6698 0 net435
rlabel metal1 211646 4658 211646 4658 0 net436
rlabel metal2 228298 4386 228298 4386 0 net437
rlabel metal2 148166 3604 148166 3604 0 net438
rlabel metal1 150880 2482 150880 2482 0 net439
rlabel metal2 78246 4998 78246 4998 0 net44
rlabel metal2 151846 4233 151846 4233 0 net440
rlabel metal1 99682 2482 99682 2482 0 net441
rlabel metal1 116702 2924 116702 2924 0 net442
rlabel metal2 112102 6732 112102 6732 0 net443
rlabel metal1 81788 4522 81788 4522 0 net444
rlabel metal1 89654 5100 89654 5100 0 net445
rlabel metal2 88090 5032 88090 5032 0 net446
rlabel metal1 39652 1938 39652 1938 0 net447
rlabel metal2 43654 5729 43654 5729 0 net448
rlabel metal2 47978 5287 47978 5287 0 net449
rlabel metal1 77510 1972 77510 1972 0 net45
rlabel metal2 109342 6596 109342 6596 0 net450
rlabel metal1 106536 2278 106536 2278 0 net451
rlabel metal2 110998 5950 110998 5950 0 net452
rlabel metal2 80914 4692 80914 4692 0 net453
rlabel metal2 149178 3196 149178 3196 0 net454
rlabel metal2 151846 4794 151846 4794 0 net455
rlabel metal1 156722 2958 156722 2958 0 net456
rlabel via1 211462 2958 211462 2958 0 net457
rlabel metal2 219006 7548 219006 7548 0 net458
rlabel metal2 221490 6239 221490 6239 0 net459
rlabel metal2 11178 2380 11178 2380 0 net46
rlabel metal1 189244 4998 189244 4998 0 net460
rlabel metal1 39974 1911 39974 1911 0 net461
rlabel metal2 48070 4420 48070 4420 0 net462
rlabel metal1 46690 4114 46690 4114 0 net463
rlabel metal2 108790 7276 108790 7276 0 net464
rlabel metal1 99038 3400 99038 3400 0 net465
rlabel metal1 110354 4726 110354 4726 0 net466
rlabel metal1 79994 5134 79994 5134 0 net467
rlabel metal2 148902 2655 148902 2655 0 net468
rlabel metal2 154514 3876 154514 3876 0 net469
rlabel metal2 76774 1564 76774 1564 0 net47
rlabel metal1 170016 6630 170016 6630 0 net470
rlabel metal1 213302 2856 213302 2856 0 net471
rlabel metal2 213486 4386 213486 4386 0 net472
rlabel metal1 230230 6630 230230 6630 0 net473
rlabel metal2 172546 7038 172546 7038 0 net474
rlabel metal1 58788 2618 58788 2618 0 net475
rlabel metal1 196834 1938 196834 1938 0 net476
rlabel metal1 59570 1326 59570 1326 0 net477
rlabel via1 212566 9707 212566 9707 0 net478
rlabel metal2 137310 9520 137310 9520 0 net479
rlabel metal1 76038 2006 76038 2006 0 net48
rlabel metal2 231518 2349 231518 2349 0 net480
rlabel metal1 129398 1972 129398 1972 0 net481
rlabel metal1 212014 6664 212014 6664 0 net482
rlabel metal2 61594 4419 61594 4419 0 net483
rlabel metal3 266593 2652 266593 2652 0 net484
rlabel metal2 62422 9656 62422 9656 0 net485
rlabel metal1 267122 1870 267122 1870 0 net486
rlabel metal2 63250 9792 63250 9792 0 net487
rlabel metal3 268157 2516 268157 2516 0 net488
rlabel metal1 132894 1326 132894 1326 0 net489
rlabel metal2 75026 952 75026 952 0 net49
rlabel metal1 270112 1870 270112 1870 0 net490
rlabel metal1 133170 1938 133170 1938 0 net491
rlabel metal1 202308 1938 202308 1938 0 net492
rlabel metal1 120934 1972 120934 1972 0 net493
rlabel metal2 190854 2159 190854 2159 0 net494
rlabel metal2 121670 1717 121670 1717 0 net495
rlabel metal2 191130 1445 191130 1445 0 net496
rlabel metal1 78154 2448 78154 2448 0 net497
rlabel metal1 192142 1972 192142 1972 0 net498
rlabel metal1 158838 2346 158838 2346 0 net499
rlabel metal1 269330 7922 269330 7922 0 net5
rlabel metal1 74566 1836 74566 1836 0 net50
rlabel metal1 192970 1972 192970 1972 0 net500
rlabel metal1 55476 1938 55476 1938 0 net501
rlabel metal1 193476 1938 193476 1938 0 net502
rlabel metal1 159252 1394 159252 1394 0 net503
rlabel metal1 227930 1938 227930 1938 0 net504
rlabel metal2 137310 8738 137310 8738 0 net505
rlabel metal2 195454 4419 195454 4419 0 net506
rlabel metal1 58236 1870 58236 1870 0 net507
rlabel metal1 209760 8500 209760 8500 0 net508
rlabel metal1 133952 1326 133952 1326 0 net509
rlabel metal2 73830 1530 73830 1530 0 net51
rlabel metal3 267559 1700 267559 1700 0 net510
rlabel metal1 226458 3094 226458 3094 0 net511
rlabel metal2 239246 4794 239246 4794 0 net512
rlabel metal2 251482 4896 251482 4896 0 net513
rlabel metal1 270710 6732 270710 6732 0 net514
rlabel metal1 265374 5644 265374 5644 0 net515
rlabel metal2 264730 5916 264730 5916 0 net516
rlabel metal3 272121 8772 272121 8772 0 net517
rlabel metal1 266248 3026 266248 3026 0 net518
rlabel metal3 272121 1020 272121 1020 0 net519
rlabel metal2 72450 884 72450 884 0 net52
rlabel metal4 828 779 828 779 0 net520
rlabel metal1 1610 9146 1610 9146 0 net521
rlabel metal4 34960 235 34960 235 0 net522
rlabel metal2 35190 9707 35190 9707 0 net523
rlabel metal4 69092 439 69092 439 0 net524
rlabel via2 69138 9571 69138 9571 0 net525
rlabel metal4 103224 303 103224 303 0 net526
rlabel metal2 103270 9911 103270 9911 0 net527
rlabel metal4 137356 779 137356 779 0 net528
rlabel via2 137402 9571 137402 9571 0 net529
rlabel metal1 79534 6392 79534 6392 0 net53
rlabel metal4 171488 235 171488 235 0 net530
rlabel metal2 171718 9911 171718 9911 0 net531
rlabel metal4 205620 235 205620 235 0 net532
rlabel via2 205850 9571 205850 9571 0 net533
rlabel metal4 239752 235 239752 235 0 net534
rlabel metal2 239706 9911 239706 9911 0 net535
rlabel metal1 32430 1972 32430 1972 0 net536
rlabel metal1 32752 8398 32752 8398 0 net537
rlabel metal2 66654 2108 66654 2108 0 net538
rlabel metal1 67068 8398 67068 8398 0 net539
rlabel metal2 73186 2652 73186 2652 0 net54
rlabel metal2 99866 1598 99866 1598 0 net540
rlabel metal1 100050 7922 100050 7922 0 net541
rlabel metal1 134182 1972 134182 1972 0 net542
rlabel metal2 134274 8636 134274 8636 0 net543
rlabel metal2 167762 2686 167762 2686 0 net544
rlabel metal2 169602 8160 169602 8160 0 net545
rlabel metal2 202354 2176 202354 2176 0 net546
rlabel metal1 202998 7922 202998 7922 0 net547
rlabel metal1 236210 1870 236210 1870 0 net548
rlabel metal1 235796 7854 235796 7854 0 net549
rlabel metal2 70886 2244 70886 2244 0 net55
rlabel metal2 267582 2142 267582 2142 0 net550
rlabel metal1 266386 5678 266386 5678 0 net551
rlabel metal3 272190 8908 272190 8908 0 net552
rlabel metal2 69874 1156 69874 1156 0 net56
rlabel metal3 16560 1088 16560 1088 0 net57
rlabel metal2 87078 8517 87078 8517 0 net58
rlabel metal2 86618 8245 86618 8245 0 net59
rlabel metal1 270802 4046 270802 4046 0 net6
rlabel metal2 85606 8432 85606 8432 0 net60
rlabel metal2 84870 8874 84870 8874 0 net61
rlabel metal2 84134 8449 84134 8449 0 net62
rlabel metal2 82754 8653 82754 8653 0 net63
rlabel metal2 82662 8177 82662 8177 0 net64
rlabel metal2 81926 8160 81926 8160 0 net65
rlabel metal1 80776 9486 80776 9486 0 net66
rlabel metal2 80178 8126 80178 8126 0 net67
rlabel metal2 9706 952 9706 952 0 net68
rlabel metal1 79718 8330 79718 8330 0 net69
rlabel metal1 269146 7922 269146 7922 0 net7
rlabel metal2 78890 8092 78890 8092 0 net70
rlabel metal2 77602 8466 77602 8466 0 net71
rlabel metal2 77510 9588 77510 9588 0 net72
rlabel metal2 76774 9214 76774 9214 0 net73
rlabel metal1 77786 6834 77786 6834 0 net74
rlabel metal2 75026 9826 75026 9826 0 net75
rlabel metal1 78752 4794 78752 4794 0 net76
rlabel metal2 82202 5593 82202 5593 0 net77
rlabel metal1 74520 9588 74520 9588 0 net78
rlabel metal2 9246 2992 9246 2992 0 net79
rlabel metal1 267030 5848 267030 5848 0 net8
rlabel metal1 72358 8874 72358 8874 0 net80
rlabel metal1 79534 6256 79534 6256 0 net81
rlabel metal1 96738 2516 96738 2516 0 net82
rlabel metal2 69874 8364 69874 8364 0 net83
rlabel metal1 120888 1190 120888 1190 0 net84
rlabel via1 120210 3502 120210 3502 0 net85
rlabel metal1 119232 1190 119232 1190 0 net86
rlabel via1 118519 5134 118519 5134 0 net87
rlabel metal1 117576 1190 117576 1190 0 net88
rlabel metal1 116840 2074 116840 2074 0 net89
rlabel metal2 268226 6885 268226 6885 0 net9
rlabel metal2 40296 2652 40296 2652 0 net90
rlabel metal1 116196 1190 116196 1190 0 net91
rlabel metal2 113390 1343 113390 1343 0 net92
rlabel metal1 113758 4522 113758 4522 0 net93
rlabel metal1 113482 1292 113482 1292 0 net94
rlabel metal2 113298 1360 113298 1360 0 net95
rlabel metal2 112746 952 112746 952 0 net96
rlabel metal1 109342 2074 109342 2074 0 net97
rlabel metal2 111366 2618 111366 2618 0 net98
rlabel metal1 110630 1224 110630 1224 0 net99
rlabel metal3 272190 7276 272190 7276 0 spine_iw[10]
rlabel metal2 262522 6953 262522 6953 0 spine_iw[11]
rlabel metal3 270212 7004 270212 7004 0 spine_iw[12]
rlabel metal3 270258 6868 270258 6868 0 spine_iw[13]
rlabel metal3 272236 6732 272236 6732 0 spine_iw[14]
rlabel metal3 272144 6596 272144 6596 0 spine_iw[15]
rlabel metal3 272121 6460 272121 6460 0 spine_iw[16]
rlabel metal3 272190 6324 272190 6324 0 spine_iw[17]
rlabel metal3 270672 6188 270672 6188 0 spine_iw[18]
rlabel metal3 272098 6052 272098 6052 0 spine_iw[19]
rlabel metal3 271500 8500 271500 8500 0 spine_iw[1]
rlabel metal3 272052 5916 272052 5916 0 spine_iw[20]
rlabel metal3 271937 5780 271937 5780 0 spine_iw[21]
rlabel metal3 271845 5644 271845 5644 0 spine_iw[22]
rlabel metal3 272098 5508 272098 5508 0 spine_iw[23]
rlabel metal3 272190 5372 272190 5372 0 spine_iw[24]
rlabel metal1 268410 2346 268410 2346 0 spine_iw[25]
rlabel metal3 272190 5100 272190 5100 0 spine_iw[26]
rlabel metal3 270258 4964 270258 4964 0 spine_iw[27]
rlabel metal3 270626 4828 270626 4828 0 spine_iw[28]
rlabel metal3 272282 4692 272282 4692 0 spine_iw[29]
rlabel metal3 271822 8364 271822 8364 0 spine_iw[2]
rlabel metal1 270342 7378 270342 7378 0 spine_iw[3]
rlabel metal3 271362 8092 271362 8092 0 spine_iw[4]
rlabel metal3 271270 7956 271270 7956 0 spine_iw[5]
rlabel metal3 270212 7820 270212 7820 0 spine_iw[6]
rlabel metal3 272098 7684 272098 7684 0 spine_iw[7]
rlabel metal3 272098 7548 272098 7548 0 spine_iw[8]
rlabel metal3 270212 7412 270212 7412 0 spine_iw[9]
rlabel metal2 252402 3264 252402 3264 0 spine_ow[10]
rlabel metal3 272190 2924 272190 2924 0 spine_ow[11]
rlabel metal3 271592 2788 271592 2788 0 spine_ow[12]
rlabel metal3 269798 2652 269798 2652 0 spine_ow[13]
rlabel via2 223238 3043 223238 3043 0 spine_ow[14]
rlabel metal3 272190 2380 272190 2380 0 spine_ow[15]
rlabel metal3 272121 2244 272121 2244 0 spine_ow[16]
rlabel metal3 272098 2108 272098 2108 0 spine_ow[17]
rlabel metal3 272282 1972 272282 1972 0 spine_ow[18]
rlabel metal3 271293 1836 271293 1836 0 spine_ow[19]
rlabel metal2 245410 4352 245410 4352 0 spine_ow[1]
rlabel metal3 271201 1700 271201 1700 0 spine_ow[20]
rlabel metal3 270718 1564 270718 1564 0 spine_ow[21]
rlabel metal3 270626 1428 270626 1428 0 spine_ow[22]
rlabel metal3 270649 1292 270649 1292 0 spine_ow[23]
rlabel metal3 272098 1156 272098 1156 0 spine_ow[24]
rlabel metal2 244214 4063 244214 4063 0 spine_ow[2]
rlabel metal3 271845 4012 271845 4012 0 spine_ow[3]
rlabel metal3 271937 3876 271937 3876 0 spine_ow[4]
rlabel metal3 272006 3740 272006 3740 0 spine_ow[5]
rlabel metal3 270166 3604 270166 3604 0 spine_ow[6]
rlabel metal3 272190 3468 272190 3468 0 spine_ow[7]
rlabel metal3 272121 3332 272121 3332 0 spine_ow[8]
rlabel metal3 272098 3196 272098 3196 0 spine_ow[9]
rlabel metal1 264684 7378 264684 7378 0 tbuf_row_ena_I.t
rlabel metal1 239108 5202 239108 5202 0 tbuf_row_ena_I.tx
rlabel metal1 244858 4522 244858 4522 0 tbuf_spine_ow_I\[0\].z
rlabel metal1 260636 4182 260636 4182 0 tbuf_spine_ow_I\[10\].z
rlabel metal1 258658 3502 258658 3502 0 tbuf_spine_ow_I\[11\].z
rlabel metal1 259808 3094 259808 3094 0 tbuf_spine_ow_I\[12\].z
rlabel metal1 222594 3026 222594 3026 0 tbuf_spine_ow_I\[13\].z
rlabel metal1 219190 1938 219190 1938 0 tbuf_spine_ow_I\[14\].z
rlabel metal2 216430 2108 216430 2108 0 tbuf_spine_ow_I\[15\].z
rlabel metal1 217994 2822 217994 2822 0 tbuf_spine_ow_I\[16\].z
rlabel metal1 218454 1326 218454 1326 0 tbuf_spine_ow_I\[17\].z
rlabel metal1 219834 1972 219834 1972 0 tbuf_spine_ow_I\[18\].z
rlabel metal2 220754 2142 220754 2142 0 tbuf_spine_ow_I\[19\].z
rlabel metal1 243616 4182 243616 4182 0 tbuf_spine_ow_I\[1\].z
rlabel metal1 227792 2414 227792 2414 0 tbuf_spine_ow_I\[20\].z
rlabel metal1 222732 1938 222732 1938 0 tbuf_spine_ow_I\[21\].z
rlabel metal1 223882 1972 223882 1972 0 tbuf_spine_ow_I\[22\].z
rlabel metal2 223790 1802 223790 1802 0 tbuf_spine_ow_I\[23\].z
rlabel metal1 241960 4182 241960 4182 0 tbuf_spine_ow_I\[2\].z
rlabel metal1 240074 4182 240074 4182 0 tbuf_spine_ow_I\[3\].z
rlabel metal1 253253 3978 253253 3978 0 tbuf_spine_ow_I\[4\].z
rlabel metal1 259992 3434 259992 3434 0 tbuf_spine_ow_I\[5\].z
rlabel metal2 260222 4233 260222 4233 0 tbuf_spine_ow_I\[6\].z
rlabel metal2 258106 3706 258106 3706 0 tbuf_spine_ow_I\[7\].z
rlabel metal1 258704 4182 258704 4182 0 tbuf_spine_ow_I\[8\].z
rlabel metal1 252034 3502 252034 3502 0 tbuf_spine_ow_I\[9\].z
rlabel metal4 32476 779 32476 779 0 um_ena[0]
rlabel metal4 203136 235 203136 235 0 um_ena[10]
rlabel metal2 204102 9707 204102 9707 0 um_ena[11]
rlabel metal4 237268 779 237268 779 0 um_ena[12]
rlabel metal1 237452 9146 237452 9146 0 um_ena[13]
rlabel metal4 271400 235 271400 235 0 um_ena[14]
rlabel metal1 270342 3706 270342 3706 0 um_ena[15]
rlabel metal2 32614 9503 32614 9503 0 um_ena[1]
rlabel metal4 66608 303 66608 303 0 um_ena[2]
rlabel metal2 66930 9979 66930 9979 0 um_ena[3]
rlabel metal4 100740 507 100740 507 0 um_ena[4]
rlabel via2 100694 9707 100694 9707 0 um_ena[5]
rlabel metal4 134872 235 134872 235 0 um_ena[6]
rlabel metal2 134918 9673 134918 9673 0 um_ena[7]
rlabel metal4 169004 371 169004 371 0 um_ena[8]
rlabel metal1 169786 9146 169786 9146 0 um_ena[9]
rlabel metal2 32522 833 32522 833 0 um_iw[0]
rlabel metal2 93334 8177 93334 8177 0 um_iw[100]
rlabel metal1 92276 8602 92276 8602 0 um_iw[101]
rlabel metal2 91862 8687 91862 8687 0 um_iw[102]
rlabel metal1 90804 8602 90804 8602 0 um_iw[103]
rlabel metal2 90390 9979 90390 9979 0 um_iw[104]
rlabel metal4 88964 9421 88964 9421 0 um_iw[105]
rlabel metal1 88412 9146 88412 9146 0 um_iw[106]
rlabel metal1 88688 8602 88688 8602 0 um_iw[107]
rlabel metal4 134136 371 134136 371 0 um_iw[108]
rlabel metal4 133400 371 133400 371 0 um_iw[109]
rlabel metal3 24449 3332 24449 3332 0 um_iw[10]
rlabel metal4 132664 371 132664 371 0 um_iw[110]
rlabel metal4 131928 371 131928 371 0 um_iw[111]
rlabel metal4 131192 371 131192 371 0 um_iw[112]
rlabel metal4 130456 235 130456 235 0 um_iw[113]
rlabel metal4 129720 371 129720 371 0 um_iw[114]
rlabel metal4 128984 371 128984 371 0 um_iw[115]
rlabel metal4 128248 235 128248 235 0 um_iw[116]
rlabel metal4 127512 371 127512 371 0 um_iw[117]
rlabel metal4 126776 371 126776 371 0 um_iw[118]
rlabel metal4 126040 371 126040 371 0 um_iw[119]
rlabel metal4 23644 371 23644 371 0 um_iw[11]
rlabel metal4 125304 371 125304 371 0 um_iw[120]
rlabel metal4 124568 371 124568 371 0 um_iw[121]
rlabel metal4 123832 371 123832 371 0 um_iw[122]
rlabel metal4 123096 371 123096 371 0 um_iw[123]
rlabel metal4 122360 371 122360 371 0 um_iw[124]
rlabel metal4 121624 371 121624 371 0 um_iw[125]
rlabel metal2 134274 9979 134274 9979 0 um_iw[126]
rlabel metal2 133538 9979 133538 9979 0 um_iw[127]
rlabel metal2 133078 9163 133078 9163 0 um_iw[128]
rlabel metal2 132342 9435 132342 9435 0 um_iw[129]
rlabel via3 22931 2924 22931 2924 0 um_iw[12]
rlabel metal2 131514 9979 131514 9979 0 um_iw[130]
rlabel metal1 131054 8602 131054 8602 0 um_iw[131]
rlabel metal1 129628 9690 129628 9690 0 um_iw[132]
rlabel metal2 128846 9979 128846 9979 0 um_iw[133]
rlabel metal2 127834 9775 127834 9775 0 um_iw[134]
rlabel metal2 127926 9979 127926 9979 0 um_iw[135]
rlabel metal1 126960 8602 126960 8602 0 um_iw[136]
rlabel metal2 126362 9435 126362 9435 0 um_iw[137]
rlabel metal1 125488 8602 125488 8602 0 um_iw[138]
rlabel metal2 125258 9979 125258 9979 0 um_iw[139]
rlabel metal1 23736 2618 23736 2618 0 um_iw[13]
rlabel metal2 123970 9435 123970 9435 0 um_iw[140]
rlabel metal2 123234 9435 123234 9435 0 um_iw[141]
rlabel metal2 122682 9979 122682 9979 0 um_iw[142]
rlabel metal1 121210 9146 121210 9146 0 um_iw[143]
rlabel metal4 168268 779 168268 779 0 um_iw[144]
rlabel metal4 167532 371 167532 371 0 um_iw[145]
rlabel metal4 166796 643 166796 643 0 um_iw[146]
rlabel metal4 166060 643 166060 643 0 um_iw[147]
rlabel metal4 165324 643 165324 643 0 um_iw[148]
rlabel metal4 164588 371 164588 371 0 um_iw[149]
rlabel metal4 21436 915 21436 915 0 um_iw[14]
rlabel metal4 163852 779 163852 779 0 um_iw[150]
rlabel metal4 163116 643 163116 643 0 um_iw[151]
rlabel metal4 162380 371 162380 371 0 um_iw[152]
rlabel metal4 161644 643 161644 643 0 um_iw[153]
rlabel metal4 160908 371 160908 371 0 um_iw[154]
rlabel metal4 160172 643 160172 643 0 um_iw[155]
rlabel metal1 160356 2618 160356 2618 0 um_iw[156]
rlabel metal4 158700 371 158700 371 0 um_iw[157]
rlabel metal4 157964 779 157964 779 0 um_iw[158]
rlabel metal1 157642 2618 157642 2618 0 um_iw[159]
rlabel metal4 20700 779 20700 779 0 um_iw[15]
rlabel metal2 157458 1853 157458 1853 0 um_iw[160]
rlabel metal4 155756 779 155756 779 0 um_iw[161]
rlabel metal1 168728 8058 168728 8058 0 um_iw[162]
rlabel metal2 167854 8211 167854 8211 0 um_iw[163]
rlabel metal4 166796 9489 166796 9489 0 um_iw[164]
rlabel metal2 166382 8211 166382 8211 0 um_iw[165]
rlabel metal2 165554 7939 165554 7939 0 um_iw[166]
rlabel metal2 164818 7939 164818 7939 0 um_iw[167]
rlabel metal1 164772 9690 164772 9690 0 um_iw[168]
rlabel metal2 164082 7939 164082 7939 0 um_iw[169]
rlabel via3 19987 2788 19987 2788 0 um_iw[16]
rlabel metal2 162610 7939 162610 7939 0 um_iw[170]
rlabel metal1 162380 8058 162380 8058 0 um_iw[171]
rlabel metal2 161322 7939 161322 7939 0 um_iw[172]
rlabel metal2 160310 8211 160310 8211 0 um_iw[173]
rlabel metal1 159850 9690 159850 9690 0 um_iw[174]
rlabel via2 159482 9435 159482 9435 0 um_iw[175]
rlabel metal1 158378 9690 158378 9690 0 um_iw[176]
rlabel metal4 157228 10509 157228 10509 0 um_iw[177]
rlabel via2 156906 9707 156906 9707 0 um_iw[178]
rlabel metal1 156078 9690 156078 9690 0 um_iw[179]
rlabel via3 19251 2924 19251 2924 0 um_iw[17]
rlabel metal4 202400 235 202400 235 0 um_iw[180]
rlabel metal4 201664 235 201664 235 0 um_iw[181]
rlabel metal4 200928 235 200928 235 0 um_iw[182]
rlabel metal4 200192 235 200192 235 0 um_iw[183]
rlabel metal4 199456 235 199456 235 0 um_iw[184]
rlabel metal4 198720 235 198720 235 0 um_iw[185]
rlabel metal4 197984 235 197984 235 0 um_iw[186]
rlabel metal4 197248 235 197248 235 0 um_iw[187]
rlabel metal4 196512 235 196512 235 0 um_iw[188]
rlabel metal4 195776 235 195776 235 0 um_iw[189]
rlabel metal1 32706 9146 32706 9146 0 um_iw[18]
rlabel metal4 195040 235 195040 235 0 um_iw[190]
rlabel metal4 194304 235 194304 235 0 um_iw[191]
rlabel metal4 193568 235 193568 235 0 um_iw[192]
rlabel metal4 192832 235 192832 235 0 um_iw[193]
rlabel metal4 192096 235 192096 235 0 um_iw[194]
rlabel metal4 191360 235 191360 235 0 um_iw[195]
rlabel metal4 190624 235 190624 235 0 um_iw[196]
rlabel metal1 190532 2618 190532 2618 0 um_iw[197]
rlabel metal1 202952 9690 202952 9690 0 um_iw[198]
rlabel metal2 202538 9979 202538 9979 0 um_iw[199]
rlabel via2 31326 8619 31326 8619 0 um_iw[19]
rlabel metal4 31004 235 31004 235 0 um_iw[1]
rlabel metal1 201296 8602 201296 8602 0 um_iw[200]
rlabel metal2 200882 9435 200882 9435 0 um_iw[201]
rlabel metal2 200054 9979 200054 9979 0 um_iw[202]
rlabel metal2 199502 9503 199502 9503 0 um_iw[203]
rlabel metal1 198444 9690 198444 9690 0 um_iw[204]
rlabel metal1 197708 9418 197708 9418 0 um_iw[205]
rlabel metal1 196972 9690 196972 9690 0 um_iw[206]
rlabel metal2 195822 9979 195822 9979 0 um_iw[207]
rlabel metal2 195638 9435 195638 9435 0 um_iw[208]
rlabel metal1 194626 9690 194626 9690 0 um_iw[209]
rlabel metal1 30360 8602 30360 8602 0 um_iw[20]
rlabel metal2 194258 9503 194258 9503 0 um_iw[210]
rlabel metal1 193154 9690 193154 9690 0 um_iw[211]
rlabel metal2 192602 9979 192602 9979 0 um_iw[212]
rlabel metal1 191820 8602 191820 8602 0 um_iw[213]
rlabel metal2 191314 9503 191314 9503 0 um_iw[214]
rlabel metal4 189888 10509 189888 10509 0 um_iw[215]
rlabel metal4 236532 643 236532 643 0 um_iw[216]
rlabel metal3 235865 2788 235865 2788 0 um_iw[217]
rlabel metal4 235060 303 235060 303 0 um_iw[218]
rlabel metal4 234324 235 234324 235 0 um_iw[219]
rlabel via2 29670 8619 29670 8619 0 um_iw[21]
rlabel metal4 233588 235 233588 235 0 um_iw[220]
rlabel metal4 232852 643 232852 643 0 um_iw[221]
rlabel metal4 232116 643 232116 643 0 um_iw[222]
rlabel metal4 231380 643 231380 643 0 um_iw[223]
rlabel metal4 230644 235 230644 235 0 um_iw[224]
rlabel metal4 229908 235 229908 235 0 um_iw[225]
rlabel metal4 229172 235 229172 235 0 um_iw[226]
rlabel metal4 228436 643 228436 643 0 um_iw[227]
rlabel metal4 227700 711 227700 711 0 um_iw[228]
rlabel metal4 226964 711 226964 711 0 um_iw[229]
rlabel via2 28842 9435 28842 9435 0 um_iw[22]
rlabel metal1 226734 2618 226734 2618 0 um_iw[230]
rlabel metal4 225492 779 225492 779 0 um_iw[231]
rlabel metal1 225446 2618 225446 2618 0 um_iw[232]
rlabel metal1 225538 2312 225538 2312 0 um_iw[233]
rlabel via2 236670 8619 236670 8619 0 um_iw[234]
rlabel metal1 236440 9146 236440 9146 0 um_iw[235]
rlabel via2 235106 9707 235106 9707 0 um_iw[236]
rlabel via2 234370 9707 234370 9707 0 um_iw[237]
rlabel via2 233542 9707 233542 9707 0 um_iw[238]
rlabel metal1 233174 8602 233174 8602 0 um_iw[239]
rlabel metal2 28382 8211 28382 8211 0 um_iw[23]
rlabel via2 231978 8619 231978 8619 0 um_iw[240]
rlabel metal2 231610 9537 231610 9537 0 um_iw[241]
rlabel metal2 230874 8211 230874 8211 0 um_iw[242]
rlabel via2 229862 9707 229862 9707 0 um_iw[243]
rlabel via2 229126 8619 229126 8619 0 um_iw[244]
rlabel metal1 228344 9350 228344 9350 0 um_iw[245]
rlabel via2 228298 8619 228298 8619 0 um_iw[246]
rlabel via2 226734 8619 226734 8619 0 um_iw[247]
rlabel via2 225998 8619 225998 8619 0 um_iw[248]
rlabel via2 225722 9707 225722 9707 0 um_iw[249]
rlabel metal1 28520 7718 28520 7718 0 um_iw[24]
rlabel metal4 224756 9557 224756 9557 0 um_iw[250]
rlabel metal1 223468 9078 223468 9078 0 um_iw[251]
rlabel metal4 270664 235 270664 235 0 um_iw[252]
rlabel metal4 269928 371 269928 371 0 um_iw[253]
rlabel metal4 269192 303 269192 303 0 um_iw[254]
rlabel metal4 268456 371 268456 371 0 um_iw[255]
rlabel metal2 267674 901 267674 901 0 um_iw[256]
rlabel metal4 266984 371 266984 371 0 um_iw[257]
rlabel metal4 266248 371 266248 371 0 um_iw[258]
rlabel metal4 265512 371 265512 371 0 um_iw[259]
rlabel metal2 26726 7497 26726 7497 0 um_iw[25]
rlabel metal4 264776 235 264776 235 0 um_iw[260]
rlabel metal4 264040 371 264040 371 0 um_iw[261]
rlabel metal4 263304 371 263304 371 0 um_iw[262]
rlabel metal4 262568 371 262568 371 0 um_iw[263]
rlabel metal4 261832 303 261832 303 0 um_iw[264]
rlabel metal4 261096 371 261096 371 0 um_iw[265]
rlabel metal4 260360 371 260360 371 0 um_iw[266]
rlabel metal4 259624 371 259624 371 0 um_iw[267]
rlabel metal4 258888 371 258888 371 0 um_iw[268]
rlabel metal4 258152 371 258152 371 0 um_iw[269]
rlabel metal1 29118 9350 29118 9350 0 um_iw[26]
rlabel metal1 270388 3910 270388 3910 0 um_iw[270]
rlabel metal1 269468 3638 269468 3638 0 um_iw[271]
rlabel metal1 269468 3910 269468 3910 0 um_iw[272]
rlabel metal1 267904 3978 267904 3978 0 um_iw[273]
rlabel metal2 267766 5491 267766 5491 0 um_iw[274]
rlabel metal2 266938 5219 266938 5219 0 um_iw[275]
rlabel metal4 266248 10645 266248 10645 0 um_iw[276]
rlabel metal2 265742 8449 265742 8449 0 um_iw[277]
rlabel metal1 264362 6630 264362 6630 0 um_iw[278]
rlabel metal2 264362 8891 264362 8891 0 um_iw[279]
rlabel metal1 27140 7174 27140 7174 0 um_iw[27]
rlabel metal2 263258 8891 263258 8891 0 um_iw[280]
rlabel metal2 262522 8891 262522 8891 0 um_iw[281]
rlabel metal2 261786 8891 261786 8891 0 um_iw[282]
rlabel metal1 262338 9690 262338 9690 0 um_iw[283]
rlabel metal2 260498 9163 260498 9163 0 um_iw[284]
rlabel metal2 260038 9979 260038 9979 0 um_iw[285]
rlabel metal2 259026 9163 259026 9163 0 um_iw[286]
rlabel metal2 258290 9435 258290 9435 0 um_iw[287]
rlabel via2 23506 8619 23506 8619 0 um_iw[28]
rlabel metal1 25300 6630 25300 6630 0 um_iw[29]
rlabel metal4 30268 371 30268 371 0 um_iw[2]
rlabel metal1 24104 7174 24104 7174 0 um_iw[30]
rlabel metal4 22172 10441 22172 10441 0 um_iw[31]
rlabel metal4 21436 10305 21436 10305 0 um_iw[32]
rlabel metal4 20700 10645 20700 10645 0 um_iw[33]
rlabel metal4 19964 8809 19964 8809 0 um_iw[34]
rlabel metal4 19228 8809 19228 8809 0 um_iw[35]
rlabel metal4 65872 303 65872 303 0 um_iw[36]
rlabel metal4 65136 371 65136 371 0 um_iw[37]
rlabel metal4 64400 371 64400 371 0 um_iw[38]
rlabel metal4 63664 371 63664 371 0 um_iw[39]
rlabel metal4 29532 303 29532 303 0 um_iw[3]
rlabel metal4 62928 371 62928 371 0 um_iw[40]
rlabel metal4 62192 371 62192 371 0 um_iw[41]
rlabel metal4 61456 371 61456 371 0 um_iw[42]
rlabel metal4 60720 371 60720 371 0 um_iw[43]
rlabel metal4 59984 235 59984 235 0 um_iw[44]
rlabel metal4 59248 235 59248 235 0 um_iw[45]
rlabel metal4 58512 371 58512 371 0 um_iw[46]
rlabel metal4 57776 371 57776 371 0 um_iw[47]
rlabel metal4 57040 371 57040 371 0 um_iw[48]
rlabel metal4 56304 371 56304 371 0 um_iw[49]
rlabel metal4 28796 371 28796 371 0 um_iw[4]
rlabel metal4 55568 371 55568 371 0 um_iw[50]
rlabel metal4 54832 371 54832 371 0 um_iw[51]
rlabel metal4 54096 235 54096 235 0 um_iw[52]
rlabel metal4 53360 371 53360 371 0 um_iw[53]
rlabel metal2 66194 9979 66194 9979 0 um_iw[54]
rlabel metal2 65458 9299 65458 9299 0 um_iw[55]
rlabel metal2 64630 9435 64630 9435 0 um_iw[56]
rlabel metal2 63802 9435 63802 9435 0 um_iw[57]
rlabel metal2 63434 9979 63434 9979 0 um_iw[58]
rlabel metal2 62330 9435 62330 9435 0 um_iw[59]
rlabel metal4 28060 303 28060 303 0 um_iw[5]
rlabel metal2 61594 9435 61594 9435 0 um_iw[60]
rlabel metal2 60858 9979 60858 9979 0 um_iw[61]
rlabel metal2 60030 9979 60030 9979 0 um_iw[62]
rlabel metal2 59294 9979 59294 9979 0 um_iw[63]
rlabel metal2 58650 9435 58650 9435 0 um_iw[64]
rlabel metal1 58052 9690 58052 9690 0 um_iw[65]
rlabel metal2 57086 9435 57086 9435 0 um_iw[66]
rlabel metal2 56258 9435 56258 9435 0 um_iw[67]
rlabel metal2 55522 9435 55522 9435 0 um_iw[68]
rlabel metal2 54786 9435 54786 9435 0 um_iw[69]
rlabel metal4 27324 711 27324 711 0 um_iw[6]
rlabel metal2 54694 10047 54694 10047 0 um_iw[70]
rlabel metal2 53222 9707 53222 9707 0 um_iw[71]
rlabel metal4 100004 303 100004 303 0 um_iw[72]
rlabel metal4 99268 847 99268 847 0 um_iw[73]
rlabel metal4 98532 439 98532 439 0 um_iw[74]
rlabel metal4 97796 439 97796 439 0 um_iw[75]
rlabel metal4 97060 303 97060 303 0 um_iw[76]
rlabel metal4 96324 643 96324 643 0 um_iw[77]
rlabel metal4 95588 643 95588 643 0 um_iw[78]
rlabel metal4 94852 643 94852 643 0 um_iw[79]
rlabel metal4 26588 711 26588 711 0 um_iw[7]
rlabel metal4 94116 643 94116 643 0 um_iw[80]
rlabel metal4 93380 439 93380 439 0 um_iw[81]
rlabel metal4 92644 235 92644 235 0 um_iw[82]
rlabel metal4 91908 439 91908 439 0 um_iw[83]
rlabel metal4 91172 235 91172 235 0 um_iw[84]
rlabel metal4 90436 439 90436 439 0 um_iw[85]
rlabel metal4 89700 235 89700 235 0 um_iw[86]
rlabel metal4 88964 711 88964 711 0 um_iw[87]
rlabel metal4 88228 643 88228 643 0 um_iw[88]
rlabel metal4 87492 711 87492 711 0 um_iw[89]
rlabel metal4 25852 711 25852 711 0 um_iw[8]
rlabel metal1 100602 8602 100602 8602 0 um_iw[90]
rlabel metal4 99268 9489 99268 9489 0 um_iw[91]
rlabel via2 98670 8619 98670 8619 0 um_iw[92]
rlabel metal1 98118 9690 98118 9690 0 um_iw[93]
rlabel via2 97474 8619 97474 8619 0 um_iw[94]
rlabel metal1 96646 9690 96646 9690 0 um_iw[95]
rlabel via2 96002 9707 96002 9707 0 um_iw[96]
rlabel metal1 95128 8602 95128 8602 0 um_iw[97]
rlabel via2 94622 8619 94622 8619 0 um_iw[98]
rlabel via2 93518 9707 93518 9707 0 um_iw[99]
rlabel metal3 26611 2788 26611 2788 0 um_iw[9]
rlabel metal4 18492 371 18492 371 0 um_ow[0]
rlabel metal4 83812 847 83812 847 0 um_ow[100]
rlabel metal4 83076 847 83076 847 0 um_ow[101]
rlabel metal4 82340 711 82340 711 0 um_ow[102]
rlabel metal4 81604 847 81604 847 0 um_ow[103]
rlabel metal4 80868 439 80868 439 0 um_ow[104]
rlabel metal4 80132 847 80132 847 0 um_ow[105]
rlabel metal4 79396 711 79396 711 0 um_ow[106]
rlabel metal4 78660 439 78660 439 0 um_ow[107]
rlabel metal4 77924 711 77924 711 0 um_ow[108]
rlabel metal4 77188 575 77188 575 0 um_ow[109]
rlabel metal4 11132 371 11132 371 0 um_ow[10]
rlabel metal4 76452 711 76452 711 0 um_ow[110]
rlabel metal4 75716 575 75716 575 0 um_ow[111]
rlabel metal4 74980 371 74980 371 0 um_ow[112]
rlabel metal4 74244 575 74244 575 0 um_ow[113]
rlabel metal4 73508 711 73508 711 0 um_ow[114]
rlabel metal4 72772 371 72772 371 0 um_ow[115]
rlabel metal4 72036 575 72036 575 0 um_ow[116]
rlabel metal4 71300 711 71300 711 0 um_ow[117]
rlabel metal4 70564 575 70564 575 0 um_ow[118]
rlabel metal4 69828 439 69828 439 0 um_ow[119]
rlabel metal4 10396 371 10396 371 0 um_ow[11]
rlabel metal4 86756 10645 86756 10645 0 um_ow[120]
rlabel metal4 86020 10305 86020 10305 0 um_ow[121]
rlabel metal4 85284 10305 85284 10305 0 um_ow[122]
rlabel metal4 84548 10645 84548 10645 0 um_ow[123]
rlabel metal4 83812 10577 83812 10577 0 um_ow[124]
rlabel metal1 82570 9554 82570 9554 0 um_ow[125]
rlabel metal4 82340 10577 82340 10577 0 um_ow[126]
rlabel metal4 81604 10237 81604 10237 0 um_ow[127]
rlabel metal1 79948 9554 79948 9554 0 um_ow[128]
rlabel metal1 79948 9010 79948 9010 0 um_ow[129]
rlabel metal4 9660 371 9660 371 0 um_ow[12]
rlabel metal4 79396 10237 79396 10237 0 um_ow[130]
rlabel via2 78614 9027 78614 9027 0 um_ow[131]
rlabel via2 77326 9571 77326 9571 0 um_ow[132]
rlabel metal4 77188 10577 77188 10577 0 um_ow[133]
rlabel metal4 76452 10237 76452 10237 0 um_ow[134]
rlabel via2 74750 9571 74750 9571 0 um_ow[135]
rlabel via2 74750 9027 74750 9027 0 um_ow[136]
rlabel metal4 74244 10645 74244 10645 0 um_ow[137]
rlabel via2 73462 9027 73462 9027 0 um_ow[138]
rlabel via2 72174 9571 72174 9571 0 um_ow[139]
rlabel metal4 8924 439 8924 439 0 um_ow[13]
rlabel metal4 72036 10577 72036 10577 0 um_ow[140]
rlabel metal4 71300 10645 71300 10645 0 um_ow[141]
rlabel metal1 69966 9554 69966 9554 0 um_ow[142]
rlabel via2 69598 9027 69598 9027 0 um_ow[143]
rlabel metal4 120888 371 120888 371 0 um_ow[144]
rlabel metal4 120152 371 120152 371 0 um_ow[145]
rlabel metal4 119416 371 119416 371 0 um_ow[146]
rlabel metal4 118680 371 118680 371 0 um_ow[147]
rlabel metal4 117944 371 117944 371 0 um_ow[148]
rlabel metal4 117208 235 117208 235 0 um_ow[149]
rlabel metal4 8188 371 8188 371 0 um_ow[14]
rlabel metal4 116472 371 116472 371 0 um_ow[150]
rlabel metal4 115736 371 115736 371 0 um_ow[151]
rlabel metal4 115000 371 115000 371 0 um_ow[152]
rlabel metal4 114264 371 114264 371 0 um_ow[153]
rlabel metal4 113528 235 113528 235 0 um_ow[154]
rlabel metal4 112792 303 112792 303 0 um_ow[155]
rlabel metal4 112056 303 112056 303 0 um_ow[156]
rlabel metal4 111320 303 111320 303 0 um_ow[157]
rlabel metal4 110584 303 110584 303 0 um_ow[158]
rlabel metal4 109848 303 109848 303 0 um_ow[159]
rlabel metal4 7452 439 7452 439 0 um_ow[15]
rlabel metal4 109112 303 109112 303 0 um_ow[160]
rlabel metal4 108376 303 108376 303 0 um_ow[161]
rlabel metal4 107640 303 107640 303 0 um_ow[162]
rlabel metal4 106904 303 106904 303 0 um_ow[163]
rlabel metal4 106168 303 106168 303 0 um_ow[164]
rlabel metal4 105432 303 105432 303 0 um_ow[165]
rlabel metal4 104696 303 104696 303 0 um_ow[166]
rlabel metal4 103960 303 103960 303 0 um_ow[167]
rlabel metal4 120888 10509 120888 10509 0 um_ow[168]
rlabel metal4 120152 10509 120152 10509 0 um_ow[169]
rlabel metal4 6716 575 6716 575 0 um_ow[16]
rlabel metal4 119416 10509 119416 10509 0 um_ow[170]
rlabel metal4 118680 10509 118680 10509 0 um_ow[171]
rlabel metal4 117944 10509 117944 10509 0 um_ow[172]
rlabel metal4 117208 10509 117208 10509 0 um_ow[173]
rlabel metal4 116472 10509 116472 10509 0 um_ow[174]
rlabel metal4 115736 10509 115736 10509 0 um_ow[175]
rlabel metal4 115000 10509 115000 10509 0 um_ow[176]
rlabel metal4 114264 10509 114264 10509 0 um_ow[177]
rlabel metal4 113528 10509 113528 10509 0 um_ow[178]
rlabel metal4 112792 10509 112792 10509 0 um_ow[179]
rlabel metal4 5980 439 5980 439 0 um_ow[17]
rlabel metal4 112056 10509 112056 10509 0 um_ow[180]
rlabel metal4 111320 10509 111320 10509 0 um_ow[181]
rlabel metal4 110584 10509 110584 10509 0 um_ow[182]
rlabel metal4 109848 10509 109848 10509 0 um_ow[183]
rlabel metal4 109112 10509 109112 10509 0 um_ow[184]
rlabel metal4 108376 10509 108376 10509 0 um_ow[185]
rlabel metal4 107640 10509 107640 10509 0 um_ow[186]
rlabel metal4 106904 10509 106904 10509 0 um_ow[187]
rlabel metal4 106168 10509 106168 10509 0 um_ow[188]
rlabel metal4 105432 10509 105432 10509 0 um_ow[189]
rlabel metal4 5244 439 5244 439 0 um_ow[18]
rlabel metal4 104696 10509 104696 10509 0 um_ow[190]
rlabel metal4 103960 10509 103960 10509 0 um_ow[191]
rlabel metal4 155020 711 155020 711 0 um_ow[192]
rlabel metal4 154284 439 154284 439 0 um_ow[193]
rlabel metal4 153548 371 153548 371 0 um_ow[194]
rlabel metal4 152812 439 152812 439 0 um_ow[195]
rlabel metal4 152076 439 152076 439 0 um_ow[196]
rlabel metal4 151340 439 151340 439 0 um_ow[197]
rlabel metal4 150604 439 150604 439 0 um_ow[198]
rlabel metal4 149868 575 149868 575 0 um_ow[199]
rlabel metal4 4508 575 4508 575 0 um_ow[19]
rlabel metal4 17756 371 17756 371 0 um_ow[1]
rlabel metal4 149132 439 149132 439 0 um_ow[200]
rlabel metal4 148396 439 148396 439 0 um_ow[201]
rlabel metal2 148442 969 148442 969 0 um_ow[202]
rlabel metal4 146924 439 146924 439 0 um_ow[203]
rlabel metal4 146188 439 146188 439 0 um_ow[204]
rlabel metal4 145452 439 145452 439 0 um_ow[205]
rlabel metal4 144716 779 144716 779 0 um_ow[206]
rlabel metal4 143980 439 143980 439 0 um_ow[207]
rlabel metal4 143244 439 143244 439 0 um_ow[208]
rlabel metal4 142508 575 142508 575 0 um_ow[209]
rlabel metal4 3772 371 3772 371 0 um_ow[20]
rlabel metal4 141772 371 141772 371 0 um_ow[210]
rlabel metal4 141036 439 141036 439 0 um_ow[211]
rlabel metal4 140300 711 140300 711 0 um_ow[212]
rlabel metal4 139564 303 139564 303 0 um_ow[213]
rlabel metal4 138828 439 138828 439 0 um_ow[214]
rlabel metal4 138092 371 138092 371 0 um_ow[215]
rlabel metal4 155020 10305 155020 10305 0 um_ow[216]
rlabel metal4 154284 10441 154284 10441 0 um_ow[217]
rlabel metal4 153548 10509 153548 10509 0 um_ow[218]
rlabel metal4 152812 10441 152812 10441 0 um_ow[219]
rlabel metal4 3036 439 3036 439 0 um_ow[21]
rlabel metal4 152076 10441 152076 10441 0 um_ow[220]
rlabel metal4 151340 10441 151340 10441 0 um_ow[221]
rlabel metal4 150604 10441 150604 10441 0 um_ow[222]
rlabel metal4 149868 10305 149868 10305 0 um_ow[223]
rlabel metal4 149132 10441 149132 10441 0 um_ow[224]
rlabel metal4 148396 10441 148396 10441 0 um_ow[225]
rlabel metal2 148442 9979 148442 9979 0 um_ow[226]
rlabel metal4 146924 10441 146924 10441 0 um_ow[227]
rlabel metal4 146188 10441 146188 10441 0 um_ow[228]
rlabel metal4 145452 10441 145452 10441 0 um_ow[229]
rlabel metal4 2300 575 2300 575 0 um_ow[22]
rlabel metal4 144716 10305 144716 10305 0 um_ow[230]
rlabel metal4 143980 10441 143980 10441 0 um_ow[231]
rlabel metal4 143244 10441 143244 10441 0 um_ow[232]
rlabel metal4 142508 10509 142508 10509 0 um_ow[233]
rlabel metal4 141772 10441 141772 10441 0 um_ow[234]
rlabel metal4 141036 10441 141036 10441 0 um_ow[235]
rlabel metal4 140300 10441 140300 10441 0 um_ow[236]
rlabel metal4 139564 10305 139564 10305 0 um_ow[237]
rlabel metal4 138828 10441 138828 10441 0 um_ow[238]
rlabel metal4 138092 10509 138092 10509 0 um_ow[239]
rlabel metal4 1564 711 1564 711 0 um_ow[23]
rlabel metal4 189152 235 189152 235 0 um_ow[240]
rlabel metal4 188416 235 188416 235 0 um_ow[241]
rlabel metal4 187680 235 187680 235 0 um_ow[242]
rlabel metal4 186944 235 186944 235 0 um_ow[243]
rlabel metal4 186208 235 186208 235 0 um_ow[244]
rlabel metal4 185472 235 185472 235 0 um_ow[245]
rlabel metal4 184736 235 184736 235 0 um_ow[246]
rlabel metal4 184000 235 184000 235 0 um_ow[247]
rlabel metal4 183264 235 183264 235 0 um_ow[248]
rlabel metal4 182528 235 182528 235 0 um_ow[249]
rlabel metal4 18492 10441 18492 10441 0 um_ow[24]
rlabel metal4 181792 235 181792 235 0 um_ow[250]
rlabel metal4 181056 235 181056 235 0 um_ow[251]
rlabel metal4 180320 235 180320 235 0 um_ow[252]
rlabel metal4 179584 235 179584 235 0 um_ow[253]
rlabel metal4 178848 235 178848 235 0 um_ow[254]
rlabel metal4 178112 235 178112 235 0 um_ow[255]
rlabel metal4 177376 235 177376 235 0 um_ow[256]
rlabel metal4 176640 235 176640 235 0 um_ow[257]
rlabel metal4 175904 235 175904 235 0 um_ow[258]
rlabel metal4 175168 235 175168 235 0 um_ow[259]
rlabel metal4 17756 10441 17756 10441 0 um_ow[25]
rlabel metal4 174432 235 174432 235 0 um_ow[260]
rlabel metal4 173696 235 173696 235 0 um_ow[261]
rlabel metal4 172960 235 172960 235 0 um_ow[262]
rlabel metal4 172224 235 172224 235 0 um_ow[263]
rlabel metal4 189152 10509 189152 10509 0 um_ow[264]
rlabel metal4 188416 10509 188416 10509 0 um_ow[265]
rlabel metal4 187680 10509 187680 10509 0 um_ow[266]
rlabel metal4 186944 10509 186944 10509 0 um_ow[267]
rlabel metal4 186208 10509 186208 10509 0 um_ow[268]
rlabel metal4 185472 10509 185472 10509 0 um_ow[269]
rlabel metal4 17020 10441 17020 10441 0 um_ow[26]
rlabel metal4 184736 10509 184736 10509 0 um_ow[270]
rlabel metal4 184000 10509 184000 10509 0 um_ow[271]
rlabel metal4 183264 10509 183264 10509 0 um_ow[272]
rlabel metal4 182528 10509 182528 10509 0 um_ow[273]
rlabel metal4 181792 10577 181792 10577 0 um_ow[274]
rlabel metal4 181056 10509 181056 10509 0 um_ow[275]
rlabel metal4 180320 10509 180320 10509 0 um_ow[276]
rlabel metal4 179584 10509 179584 10509 0 um_ow[277]
rlabel metal4 178848 10509 178848 10509 0 um_ow[278]
rlabel metal1 177882 9554 177882 9554 0 um_ow[279]
rlabel metal4 16284 10441 16284 10441 0 um_ow[27]
rlabel metal4 177376 10509 177376 10509 0 um_ow[280]
rlabel metal4 176640 10509 176640 10509 0 um_ow[281]
rlabel metal4 175904 10509 175904 10509 0 um_ow[282]
rlabel metal4 175168 10509 175168 10509 0 um_ow[283]
rlabel metal4 174432 10509 174432 10509 0 um_ow[284]
rlabel metal4 173696 10509 173696 10509 0 um_ow[285]
rlabel metal4 172960 10509 172960 10509 0 um_ow[286]
rlabel metal4 172224 10509 172224 10509 0 um_ow[287]
rlabel via3 223307 2788 223307 2788 0 um_ow[288]
rlabel metal4 222548 711 222548 711 0 um_ow[289]
rlabel metal4 15548 10441 15548 10441 0 um_ow[28]
rlabel metal4 221812 235 221812 235 0 um_ow[290]
rlabel metal4 221076 507 221076 507 0 um_ow[291]
rlabel metal4 220340 779 220340 779 0 um_ow[292]
rlabel metal4 219604 235 219604 235 0 um_ow[293]
rlabel metal4 218868 235 218868 235 0 um_ow[294]
rlabel metal4 218132 507 218132 507 0 um_ow[295]
rlabel metal4 217396 507 217396 507 0 um_ow[296]
rlabel metal4 216660 779 216660 779 0 um_ow[297]
rlabel metal4 215924 507 215924 507 0 um_ow[298]
rlabel metal4 215188 507 215188 507 0 um_ow[299]
rlabel metal4 14812 10441 14812 10441 0 um_ow[29]
rlabel metal4 17020 371 17020 371 0 um_ow[2]
rlabel metal4 214452 507 214452 507 0 um_ow[300]
rlabel metal4 213716 507 213716 507 0 um_ow[301]
rlabel metal4 212980 507 212980 507 0 um_ow[302]
rlabel metal4 212244 507 212244 507 0 um_ow[303]
rlabel metal4 211508 575 211508 575 0 um_ow[304]
rlabel metal4 210772 711 210772 711 0 um_ow[305]
rlabel metal4 210036 575 210036 575 0 um_ow[306]
rlabel metal4 209300 507 209300 507 0 um_ow[307]
rlabel metal4 208564 507 208564 507 0 um_ow[308]
rlabel metal4 207828 507 207828 507 0 um_ow[309]
rlabel metal4 14076 10441 14076 10441 0 um_ow[30]
rlabel metal4 207092 507 207092 507 0 um_ow[310]
rlabel metal4 206356 507 206356 507 0 um_ow[311]
rlabel metal4 223284 10441 223284 10441 0 um_ow[312]
rlabel metal4 222548 10509 222548 10509 0 um_ow[313]
rlabel metal4 221812 10509 221812 10509 0 um_ow[314]
rlabel metal4 221076 10577 221076 10577 0 um_ow[315]
rlabel metal4 220340 10509 220340 10509 0 um_ow[316]
rlabel metal4 219604 10441 219604 10441 0 um_ow[317]
rlabel metal4 218868 10441 218868 10441 0 um_ow[318]
rlabel metal4 218132 10645 218132 10645 0 um_ow[319]
rlabel metal4 13340 10305 13340 10305 0 um_ow[31]
rlabel metal4 217396 10441 217396 10441 0 um_ow[320]
rlabel metal4 216660 10305 216660 10305 0 um_ow[321]
rlabel metal4 215924 10441 215924 10441 0 um_ow[322]
rlabel metal4 215188 10509 215188 10509 0 um_ow[323]
rlabel metal4 214452 10441 214452 10441 0 um_ow[324]
rlabel metal4 213716 10441 213716 10441 0 um_ow[325]
rlabel metal4 212980 10441 212980 10441 0 um_ow[326]
rlabel metal3 212359 6868 212359 6868 0 um_ow[327]
rlabel metal4 211508 10577 211508 10577 0 um_ow[328]
rlabel metal4 210772 10441 210772 10441 0 um_ow[329]
rlabel metal4 12604 10441 12604 10441 0 um_ow[32]
rlabel metal4 210036 10577 210036 10577 0 um_ow[330]
rlabel metal4 209300 10441 209300 10441 0 um_ow[331]
rlabel metal4 208564 10441 208564 10441 0 um_ow[332]
rlabel metal4 207828 10645 207828 10645 0 um_ow[333]
rlabel metal4 207092 10441 207092 10441 0 um_ow[334]
rlabel metal4 206356 10441 206356 10441 0 um_ow[335]
rlabel metal4 257416 371 257416 371 0 um_ow[336]
rlabel metal4 256680 371 256680 371 0 um_ow[337]
rlabel metal4 255944 371 255944 371 0 um_ow[338]
rlabel metal4 255208 371 255208 371 0 um_ow[339]
rlabel metal4 11868 10441 11868 10441 0 um_ow[33]
rlabel metal4 254472 235 254472 235 0 um_ow[340]
rlabel metal4 253736 371 253736 371 0 um_ow[341]
rlabel metal4 253000 371 253000 371 0 um_ow[342]
rlabel metal4 252264 371 252264 371 0 um_ow[343]
rlabel metal4 251528 371 251528 371 0 um_ow[344]
rlabel metal4 250792 235 250792 235 0 um_ow[345]
rlabel metal4 250056 371 250056 371 0 um_ow[346]
rlabel metal4 249320 235 249320 235 0 um_ow[347]
rlabel metal4 248584 303 248584 303 0 um_ow[348]
rlabel metal2 248446 1649 248446 1649 0 um_ow[349]
rlabel metal4 11132 10305 11132 10305 0 um_ow[34]
rlabel metal2 248538 1241 248538 1241 0 um_ow[350]
rlabel metal4 246376 303 246376 303 0 um_ow[351]
rlabel metal4 245640 303 245640 303 0 um_ow[352]
rlabel metal4 244904 303 244904 303 0 um_ow[353]
rlabel metal2 244306 1649 244306 1649 0 um_ow[354]
rlabel metal4 243432 303 243432 303 0 um_ow[355]
rlabel metal4 242696 235 242696 235 0 um_ow[356]
rlabel metal4 241960 303 241960 303 0 um_ow[357]
rlabel metal4 241224 303 241224 303 0 um_ow[358]
rlabel metal4 240488 235 240488 235 0 um_ow[359]
rlabel metal4 10396 10305 10396 10305 0 um_ow[35]
rlabel metal4 257416 10509 257416 10509 0 um_ow[360]
rlabel metal4 256680 10509 256680 10509 0 um_ow[361]
rlabel metal4 255944 10509 255944 10509 0 um_ow[362]
rlabel metal4 255208 10509 255208 10509 0 um_ow[363]
rlabel metal4 254472 10509 254472 10509 0 um_ow[364]
rlabel metal4 253736 10509 253736 10509 0 um_ow[365]
rlabel metal4 253000 10509 253000 10509 0 um_ow[366]
rlabel metal4 252264 10509 252264 10509 0 um_ow[367]
rlabel metal4 251528 10509 251528 10509 0 um_ow[368]
rlabel metal4 250792 10509 250792 10509 0 um_ow[369]
rlabel metal4 9660 10645 9660 10645 0 um_ow[36]
rlabel metal4 250056 10509 250056 10509 0 um_ow[370]
rlabel metal4 249320 10509 249320 10509 0 um_ow[371]
rlabel metal4 248584 10509 248584 10509 0 um_ow[372]
rlabel metal4 247848 10509 247848 10509 0 um_ow[373]
rlabel metal4 247112 10509 247112 10509 0 um_ow[374]
rlabel metal4 246376 10509 246376 10509 0 um_ow[375]
rlabel metal4 245640 10509 245640 10509 0 um_ow[376]
rlabel metal4 244904 10509 244904 10509 0 um_ow[377]
rlabel metal4 244168 10509 244168 10509 0 um_ow[378]
rlabel metal4 243432 10509 243432 10509 0 um_ow[379]
rlabel metal4 8924 10441 8924 10441 0 um_ow[37]
rlabel metal4 242696 10509 242696 10509 0 um_ow[380]
rlabel metal4 241960 10509 241960 10509 0 um_ow[381]
rlabel metal4 241224 10509 241224 10509 0 um_ow[382]
rlabel metal4 240488 10509 240488 10509 0 um_ow[383]
rlabel metal4 8188 10305 8188 10305 0 um_ow[38]
rlabel metal4 7452 10441 7452 10441 0 um_ow[39]
rlabel metal2 16606 1683 16606 1683 0 um_ow[3]
rlabel metal4 6716 10441 6716 10441 0 um_ow[40]
rlabel metal4 5980 10441 5980 10441 0 um_ow[41]
rlabel metal4 5244 10441 5244 10441 0 um_ow[42]
rlabel metal4 4508 10441 4508 10441 0 um_ow[43]
rlabel metal4 3772 10441 3772 10441 0 um_ow[44]
rlabel metal4 3036 10305 3036 10305 0 um_ow[45]
rlabel metal4 2300 10441 2300 10441 0 um_ow[46]
rlabel metal4 1564 10441 1564 10441 0 um_ow[47]
rlabel metal4 52624 371 52624 371 0 um_ow[48]
rlabel metal4 51888 371 51888 371 0 um_ow[49]
rlabel metal4 15548 439 15548 439 0 um_ow[4]
rlabel metal4 51152 371 51152 371 0 um_ow[50]
rlabel metal4 50416 371 50416 371 0 um_ow[51]
rlabel metal4 49680 371 49680 371 0 um_ow[52]
rlabel metal4 48944 371 48944 371 0 um_ow[53]
rlabel metal4 48208 371 48208 371 0 um_ow[54]
rlabel metal4 47472 371 47472 371 0 um_ow[55]
rlabel metal4 46736 371 46736 371 0 um_ow[56]
rlabel metal4 46000 371 46000 371 0 um_ow[57]
rlabel metal4 45264 371 45264 371 0 um_ow[58]
rlabel metal4 44528 371 44528 371 0 um_ow[59]
rlabel metal4 14812 439 14812 439 0 um_ow[5]
rlabel metal4 43792 371 43792 371 0 um_ow[60]
rlabel metal4 43056 371 43056 371 0 um_ow[61]
rlabel metal4 42320 371 42320 371 0 um_ow[62]
rlabel metal4 41584 371 41584 371 0 um_ow[63]
rlabel metal4 40848 371 40848 371 0 um_ow[64]
rlabel metal4 40112 371 40112 371 0 um_ow[65]
rlabel metal4 39376 235 39376 235 0 um_ow[66]
rlabel metal4 38640 371 38640 371 0 um_ow[67]
rlabel metal4 37904 371 37904 371 0 um_ow[68]
rlabel metal4 37168 371 37168 371 0 um_ow[69]
rlabel metal4 14076 575 14076 575 0 um_ow[6]
rlabel metal4 36432 371 36432 371 0 um_ow[70]
rlabel metal4 35696 371 35696 371 0 um_ow[71]
rlabel metal4 52624 10509 52624 10509 0 um_ow[72]
rlabel metal4 51888 10509 51888 10509 0 um_ow[73]
rlabel metal4 51152 10509 51152 10509 0 um_ow[74]
rlabel metal4 50416 10509 50416 10509 0 um_ow[75]
rlabel metal4 49680 10509 49680 10509 0 um_ow[76]
rlabel metal4 48944 10509 48944 10509 0 um_ow[77]
rlabel metal4 48208 10509 48208 10509 0 um_ow[78]
rlabel metal4 47472 10509 47472 10509 0 um_ow[79]
rlabel metal4 13340 371 13340 371 0 um_ow[7]
rlabel metal4 46736 10509 46736 10509 0 um_ow[80]
rlabel metal4 46000 10509 46000 10509 0 um_ow[81]
rlabel metal4 45264 10509 45264 10509 0 um_ow[82]
rlabel metal4 44528 10509 44528 10509 0 um_ow[83]
rlabel metal4 43792 10509 43792 10509 0 um_ow[84]
rlabel metal4 43056 10509 43056 10509 0 um_ow[85]
rlabel metal4 42320 10509 42320 10509 0 um_ow[86]
rlabel metal4 41584 10509 41584 10509 0 um_ow[87]
rlabel metal4 40848 10509 40848 10509 0 um_ow[88]
rlabel metal4 40112 10509 40112 10509 0 um_ow[89]
rlabel metal4 12604 371 12604 371 0 um_ow[8]
rlabel metal4 39376 10509 39376 10509 0 um_ow[90]
rlabel metal4 38640 10509 38640 10509 0 um_ow[91]
rlabel metal4 37904 10509 37904 10509 0 um_ow[92]
rlabel metal4 37168 10509 37168 10509 0 um_ow[93]
rlabel metal4 36432 10509 36432 10509 0 um_ow[94]
rlabel metal4 35696 10509 35696 10509 0 um_ow[95]
rlabel metal4 86756 439 86756 439 0 um_ow[96]
rlabel metal4 86020 575 86020 575 0 um_ow[97]
rlabel metal4 85284 439 85284 439 0 um_ow[98]
rlabel metal1 82478 1292 82478 1292 0 um_ow[99]
rlabel metal4 11868 371 11868 371 0 um_ow[9]
rlabel metal2 231150 6426 231150 6426 0 zbuf_bus_ena_I.genblk1.l
rlabel via2 82018 5763 82018 5763 0 zbuf_bus_ena_I.z
rlabel metal1 268134 6800 268134 6800 0 zbuf_bus_iw_I\[0\].genblk1.l
rlabel metal1 266938 5338 266938 5338 0 zbuf_bus_iw_I\[10\].genblk1.l
rlabel metal2 261234 6086 261234 6086 0 zbuf_bus_iw_I\[11\].genblk1.l
rlabel metal2 261694 5882 261694 5882 0 zbuf_bus_iw_I\[12\].genblk1.l
rlabel metal1 260406 5236 260406 5236 0 zbuf_bus_iw_I\[13\].genblk1.l
rlabel metal2 262246 5542 262246 5542 0 zbuf_bus_iw_I\[14\].genblk1.l
rlabel metal2 261970 5406 261970 5406 0 zbuf_bus_iw_I\[15\].genblk1.l
rlabel metal1 263810 4624 263810 4624 0 zbuf_bus_iw_I\[16\].genblk1.l
rlabel metal1 268502 4250 268502 4250 0 zbuf_bus_iw_I\[17\].genblk1.l
rlabel metal2 269422 6732 269422 6732 0 zbuf_bus_iw_I\[1\].genblk1.l
rlabel metal1 269376 5338 269376 5338 0 zbuf_bus_iw_I\[2\].genblk1.l
rlabel metal1 268272 5338 268272 5338 0 zbuf_bus_iw_I\[3\].genblk1.l
rlabel metal1 266984 5678 266984 5678 0 zbuf_bus_iw_I\[4\].genblk1.l
rlabel metal1 266662 6324 266662 6324 0 zbuf_bus_iw_I\[5\].genblk1.l
rlabel metal1 265650 6290 265650 6290 0 zbuf_bus_iw_I\[6\].genblk1.l
rlabel metal1 266984 4726 266984 4726 0 zbuf_bus_iw_I\[7\].genblk1.l
rlabel metal1 268916 5270 268916 5270 0 zbuf_bus_iw_I\[8\].genblk1.l
rlabel via2 267766 5797 267766 5797 0 zbuf_bus_iw_I\[9\].genblk1.l
rlabel metal2 231242 7582 231242 7582 0 zbuf_bus_sel_I\[0\].genblk1.l
rlabel metal2 130318 6885 130318 6885 0 zbuf_bus_sel_I\[0\].z
rlabel metal2 235658 6732 235658 6732 0 zbuf_bus_sel_I\[1\].genblk1.l
rlabel metal1 128662 5814 128662 5814 0 zbuf_bus_sel_I\[1\].z
rlabel metal1 236118 6766 236118 6766 0 zbuf_bus_sel_I\[2\].genblk1.l
rlabel metal1 189106 6324 189106 6324 0 zbuf_bus_sel_I\[2\].z
rlabel metal1 236808 6290 236808 6290 0 zbuf_bus_sel_I\[3\].genblk1.l
rlabel metal1 190440 5848 190440 5848 0 zbuf_bus_sel_I\[3\].z
rlabel metal2 236210 7548 236210 7548 0 zbuf_bus_sel_I\[4\].genblk1.l
rlabel metal2 228114 6698 228114 6698 0 zbuf_bus_sel_I\[4\].z
<< properties >>
string FIXED_BBOX 0 0 272600 11000
<< end >>
