magic
tech sky130A
magscale 1 2
timestamp 1684775848
<< obsli1 >>
rect 1104 1071 271492 9809
<< obsm1 >>
rect 842 212 272214 10872
<< obsm2 >>
rect 846 31 272210 10878
<< metal3 >>
rect 272198 9558 272504 9618
rect 272014 9422 272504 9482
rect 268990 9286 272504 9346
rect 268070 9150 272504 9210
rect 268162 9014 272504 9074
rect 272026 8878 272504 8938
rect 271830 8742 272504 8802
rect 272304 8606 272504 8666
rect 270646 8470 272504 8530
rect 271290 8334 272504 8394
rect 270554 8198 272504 8258
rect 270370 8062 272504 8122
rect 270186 7926 272504 7986
rect 268070 7790 272504 7850
rect 271842 7654 272504 7714
rect 271842 7518 272504 7578
rect 268070 7382 272504 7442
rect 272026 7246 272504 7306
rect 262550 7110 272504 7170
rect 268070 6974 272504 7034
rect 268162 6838 272504 6898
rect 272118 6702 272504 6762
rect 271934 6566 272504 6626
rect 271830 6430 272504 6490
rect 272026 6294 272504 6354
rect 268990 6158 272504 6218
rect 271842 6022 272504 6082
rect 271750 5886 272504 5946
rect 271462 5750 272504 5810
rect 271278 5614 272504 5674
rect 271842 5478 272504 5538
rect 272026 5342 272504 5402
rect 268990 5206 272504 5266
rect 272026 5070 272504 5130
rect 268162 4934 272504 4994
rect 268898 4798 272504 4858
rect 272210 4662 272504 4722
rect 272304 4526 272504 4586
rect 271968 4390 272504 4450
rect 271830 4254 272504 4314
rect 244242 4118 272504 4178
rect 271278 3982 272504 4042
rect 271462 3846 272504 3906
rect 271658 3710 272504 3770
rect 267978 3574 272504 3634
rect 272026 3438 272504 3498
rect 271830 3302 272504 3362
rect 271842 3166 272504 3226
rect 262274 3030 272504 3090
rect 272026 2894 272504 2954
rect 270830 2758 272504 2818
rect 267242 2622 272504 2682
rect 268530 2486 272504 2546
rect 272026 2350 272504 2410
rect 271830 2214 272504 2274
rect 271842 2078 272504 2138
rect 272210 1942 272504 2002
rect 270174 1806 272504 1866
rect 269990 1670 272504 1730
rect 269082 1534 272504 1594
rect 268898 1398 272504 1458
rect 268886 1262 272504 1322
rect 271842 1126 272504 1186
rect 271830 990 272504 1050
<< obsm3 >>
rect 750 9698 272442 10845
rect 750 9562 272118 9698
rect 750 9426 271934 9562
rect 750 9290 268910 9426
rect 750 9070 267990 9290
rect 750 8934 268082 9070
rect 750 8882 271946 8934
rect 750 8662 271750 8882
rect 750 8610 272224 8662
rect 750 8390 270566 8610
rect 750 8338 271210 8390
rect 750 8202 270474 8338
rect 750 8066 270290 8202
rect 750 7930 270106 8066
rect 750 7710 267990 7930
rect 750 7522 271762 7710
rect 750 7302 267990 7522
rect 750 7250 271946 7302
rect 750 7030 262470 7250
rect 750 6894 267990 7030
rect 750 6758 268082 6894
rect 750 6706 272038 6758
rect 750 6570 271854 6706
rect 750 6350 271750 6570
rect 750 6298 271946 6350
rect 750 6078 268910 6298
rect 750 6026 271762 6078
rect 750 5890 271670 6026
rect 750 5754 271382 5890
rect 750 5534 271198 5754
rect 750 5398 271762 5534
rect 750 5346 271946 5398
rect 750 5126 268910 5346
rect 750 5074 271946 5126
rect 750 4854 268082 5074
rect 750 4718 268818 4854
rect 750 4582 272130 4718
rect 750 4530 272224 4582
rect 750 4394 271888 4530
rect 750 4258 271750 4394
rect 750 4038 244162 4258
rect 750 3902 271198 4038
rect 750 3766 271382 3902
rect 750 3714 271578 3766
rect 750 3494 267898 3714
rect 750 3442 271946 3494
rect 750 3222 271750 3442
rect 750 3170 271762 3222
rect 750 2950 262194 3170
rect 750 2898 271946 2950
rect 750 2762 270750 2898
rect 750 2542 267162 2762
rect 750 2406 268450 2542
rect 750 2354 271946 2406
rect 750 2134 271750 2354
rect 750 1998 271762 2134
rect 750 1946 272130 1998
rect 750 1810 270094 1946
rect 750 1674 269910 1810
rect 750 1538 269002 1674
rect 750 1402 268818 1538
rect 750 1182 268806 1402
rect 750 1130 271762 1182
rect 750 910 271750 1130
rect 750 35 272442 910
<< metal4 >>
rect 798 9212 858 10880
rect 1534 10164 1594 10880
rect 2270 10164 2330 10880
rect 3006 9892 3066 10880
rect 3742 10164 3802 10880
rect 4478 10164 4538 10880
rect 5214 10164 5274 10880
rect 5950 10164 6010 10880
rect 6686 10164 6746 10880
rect 7422 10164 7482 10880
rect 8158 9892 8218 10880
rect 8894 10164 8954 10880
rect 9630 10572 9690 10880
rect 10366 9892 10426 10880
rect 11102 9892 11162 10880
rect 11838 10164 11898 10880
rect 12574 10164 12634 10880
rect 13310 9892 13370 10880
rect 14046 10164 14106 10880
rect 14782 10164 14842 10880
rect 15518 10164 15578 10880
rect 16254 10164 16314 10880
rect 16990 10164 17050 10880
rect 17726 10164 17786 10880
rect 18462 10164 18522 10880
rect 19198 6900 19258 10880
rect 19934 6900 19994 10880
rect 20670 10572 20730 10880
rect 21406 9892 21466 10880
rect 22142 10164 22202 10880
rect 22878 6900 22938 10880
rect 23614 6900 23674 10880
rect 24350 8668 24410 10880
rect 25086 6900 25146 10880
rect 25822 9620 25882 10880
rect 26558 8396 26618 10880
rect 27294 7852 27354 10880
rect 28030 8396 28090 10880
rect 28766 9484 28826 10880
rect 29502 8668 29562 10880
rect 30238 8668 30298 10880
rect 30974 8668 31034 10880
rect 31710 10300 31770 10880
rect 32446 9620 32506 10880
rect 34930 10300 34990 10880
rect 35666 10300 35726 10880
rect 36402 10300 36462 10880
rect 37138 10300 37198 10880
rect 37874 10300 37934 10880
rect 38610 10300 38670 10880
rect 39346 10300 39406 10880
rect 40082 10300 40142 10880
rect 40818 10300 40878 10880
rect 41554 10300 41614 10880
rect 42290 10300 42350 10880
rect 43026 10300 43086 10880
rect 43762 10300 43822 10880
rect 44498 10300 44558 10880
rect 45234 10300 45294 10880
rect 45970 10300 46030 10880
rect 46706 10300 46766 10880
rect 47442 10300 47502 10880
rect 48178 10300 48238 10880
rect 48914 10300 48974 10880
rect 49650 10300 49710 10880
rect 50386 10300 50446 10880
rect 51122 10300 51182 10880
rect 51858 10300 51918 10880
rect 52594 10300 52654 10880
rect 53330 10300 53390 10880
rect 54066 10436 54126 10880
rect 54802 10300 54862 10880
rect 55538 10300 55598 10880
rect 56274 10300 56334 10880
rect 57010 10300 57070 10880
rect 57746 10300 57806 10880
rect 58482 10300 58542 10880
rect 59218 10300 59278 10880
rect 59954 10300 60014 10880
rect 60690 10300 60750 10880
rect 61426 10300 61486 10880
rect 62162 10300 62222 10880
rect 62898 10300 62958 10880
rect 63634 10300 63694 10880
rect 64370 10300 64430 10880
rect 65106 10300 65166 10880
rect 65842 10300 65902 10880
rect 66578 10300 66638 10880
rect 798 0 858 1396
rect 1534 0 1594 1260
rect 2270 0 2330 988
rect 3006 0 3066 716
rect 3742 0 3802 580
rect 4478 0 4538 988
rect 5214 0 5274 716
rect 5950 0 6010 716
rect 6686 0 6746 988
rect 7422 0 7482 716
rect 8158 0 8218 580
rect 8894 0 8954 716
rect 9630 0 9690 580
rect 10366 0 10426 580
rect 11102 0 11162 580
rect 11838 0 11898 580
rect 12574 0 12634 580
rect 13310 0 13370 580
rect 14046 0 14106 988
rect 14782 0 14842 716
rect 15518 0 15578 716
rect 16254 0 16314 1396
rect 16990 0 17050 580
rect 17726 0 17786 580
rect 18462 0 18522 580
rect 19198 0 19258 2892
rect 19934 0 19994 2756
rect 20670 0 20730 1396
rect 21406 0 21466 1668
rect 22142 0 22202 2756
rect 22878 0 22938 2892
rect 23614 0 23674 580
rect 24350 0 24410 3300
rect 25086 0 25146 2756
rect 25822 0 25882 1260
rect 26558 0 26618 1260
rect 27294 0 27354 1260
rect 28030 0 28090 444
rect 28766 0 28826 580
rect 29502 0 29562 444
rect 30238 0 30298 580
rect 30974 0 31034 308
rect 31710 0 31770 444
rect 32446 0 32506 1396
rect 34742 1040 35062 9840
rect 68540 1040 68860 9840
rect 69062 9620 69122 10880
rect 69798 9076 69858 10880
rect 70534 9620 70594 10880
rect 71270 10572 71330 10880
rect 72006 10436 72066 10880
rect 72742 9620 72802 10880
rect 73478 9076 73538 10880
rect 74214 10572 74274 10880
rect 74950 9076 75010 10880
rect 75686 9620 75746 10880
rect 76422 9756 76482 10880
rect 77158 10436 77218 10880
rect 77894 9620 77954 10880
rect 78630 9076 78690 10880
rect 79366 9756 79426 10880
rect 80102 9076 80162 10880
rect 80838 9620 80898 10880
rect 81574 9756 81634 10880
rect 82310 10436 82370 10880
rect 83046 9620 83106 10880
rect 83782 10436 83842 10880
rect 84518 10572 84578 10880
rect 85254 9892 85314 10880
rect 85990 9892 86050 10880
rect 86726 10572 86786 10880
rect 87462 8668 87522 10880
rect 88198 9212 88258 10880
rect 88934 8124 88994 10880
rect 89670 10300 89730 10880
rect 90406 8668 90466 10880
rect 91142 8804 91202 10880
rect 91878 8668 91938 10880
rect 92614 8396 92674 10880
rect 93350 9756 93410 10880
rect 94086 8668 94146 10880
rect 94822 8668 94882 10880
rect 95558 9756 95618 10880
rect 96294 9756 96354 10880
rect 97030 8668 97090 10880
rect 97766 9756 97826 10880
rect 98502 8668 98562 10880
rect 99238 8260 99298 10880
rect 99974 8668 100034 10880
rect 100710 9756 100770 10880
rect 103194 10300 103254 10880
rect 103930 10300 103990 10880
rect 104666 10300 104726 10880
rect 105402 10300 105462 10880
rect 106138 10300 106198 10880
rect 106874 10300 106934 10880
rect 107610 10300 107670 10880
rect 108346 10300 108406 10880
rect 109082 10300 109142 10880
rect 109818 10300 109878 10880
rect 110554 10300 110614 10880
rect 111290 10300 111350 10880
rect 112026 10300 112086 10880
rect 112762 10300 112822 10880
rect 113498 10300 113558 10880
rect 114234 10300 114294 10880
rect 114970 10300 115030 10880
rect 115706 10300 115766 10880
rect 116442 10300 116502 10880
rect 117178 10300 117238 10880
rect 117914 10300 117974 10880
rect 118650 10300 118710 10880
rect 119386 10300 119446 10880
rect 120122 10300 120182 10880
rect 120858 10300 120918 10880
rect 121594 10300 121654 10880
rect 122330 10300 122390 10880
rect 123066 10300 123126 10880
rect 123802 10300 123862 10880
rect 124538 10300 124598 10880
rect 125274 10436 125334 10880
rect 126010 10300 126070 10880
rect 126746 10300 126806 10880
rect 127482 10300 127542 10880
rect 128218 10436 128278 10880
rect 128954 10300 129014 10880
rect 129690 10300 129750 10880
rect 130426 10300 130486 10880
rect 131162 10300 131222 10880
rect 131898 10300 131958 10880
rect 132634 10300 132694 10880
rect 133370 10300 133430 10880
rect 134106 10300 134166 10880
rect 134842 10300 134902 10880
rect 34930 0 34990 308
rect 35666 0 35726 580
rect 36402 0 36462 580
rect 37138 0 37198 580
rect 37874 0 37934 580
rect 38610 0 38670 580
rect 39346 0 39406 308
rect 40082 0 40142 580
rect 40818 0 40878 580
rect 41554 0 41614 580
rect 42290 0 42350 580
rect 43026 0 43086 580
rect 43762 0 43822 580
rect 44498 0 44558 580
rect 45234 0 45294 580
rect 45970 0 46030 580
rect 46706 0 46766 580
rect 47442 0 47502 580
rect 48178 0 48238 580
rect 48914 0 48974 580
rect 49650 0 49710 580
rect 50386 0 50446 580
rect 51122 0 51182 580
rect 51858 0 51918 580
rect 52594 0 52654 580
rect 53330 0 53390 580
rect 54066 0 54126 370
rect 54802 0 54862 580
rect 55538 0 55598 580
rect 56274 0 56334 580
rect 57010 0 57070 580
rect 57746 0 57806 580
rect 58482 0 58542 580
rect 59218 0 59278 370
rect 59954 0 60014 370
rect 60690 0 60750 580
rect 61426 0 61486 580
rect 62162 0 62222 580
rect 62898 0 62958 580
rect 63634 0 63694 580
rect 64370 0 64430 580
rect 65106 0 65166 580
rect 65842 0 65902 444
rect 66578 0 66638 444
rect 69062 0 69122 716
rect 69798 0 69858 716
rect 70534 0 70594 988
rect 71270 0 71330 1260
rect 72006 0 72066 988
rect 72742 0 72802 580
rect 73478 0 73538 1260
rect 74214 0 74274 988
rect 74950 0 75010 580
rect 75686 0 75746 988
rect 76422 0 76482 1260
rect 77158 0 77218 988
rect 77894 0 77954 1260
rect 78630 0 78690 716
rect 79366 0 79426 1260
rect 80102 0 80162 1532
rect 80838 0 80898 716
rect 81574 0 81634 1532
rect 82310 0 82370 1260
rect 83046 0 83106 1532
rect 83782 0 83842 1532
rect 84518 0 84578 716
rect 85254 0 85314 716
rect 85990 0 86050 988
rect 86726 0 86786 716
rect 87462 0 87522 1260
rect 88198 0 88258 1124
rect 88934 0 88994 1260
rect 89670 0 89730 308
rect 90406 0 90466 716
rect 91142 0 91202 308
rect 91878 0 91938 716
rect 92614 0 92674 308
rect 93350 0 93410 716
rect 94086 0 94146 1124
rect 94822 0 94882 1124
rect 95558 0 95618 1124
rect 96294 0 96354 1124
rect 97030 0 97090 444
rect 97766 0 97826 716
rect 98502 0 98562 716
rect 99238 0 99298 1532
rect 102339 1040 102659 9840
rect 136137 1040 136457 9840
rect 137326 9620 137386 10880
rect 138062 10300 138122 10880
rect 138798 10164 138858 10880
rect 139534 9892 139594 10880
rect 140270 10164 140330 10880
rect 141006 10164 141066 10880
rect 141742 10164 141802 10880
rect 142478 10300 142538 10880
rect 143214 10164 143274 10880
rect 143950 10164 144010 10880
rect 144686 9892 144746 10880
rect 145422 10164 145482 10880
rect 146158 10164 146218 10880
rect 146894 10164 146954 10880
rect 147630 10436 147690 10880
rect 148366 10164 148426 10880
rect 149102 10164 149162 10880
rect 149838 9892 149898 10880
rect 150574 10164 150634 10880
rect 151310 10164 151370 10880
rect 152046 10164 152106 10880
rect 152782 10164 152842 10880
rect 153518 10300 153578 10880
rect 154254 10164 154314 10880
rect 154990 9892 155050 10880
rect 155726 9756 155786 10880
rect 156462 9756 156522 10880
rect 157198 10300 157258 10880
rect 157934 9756 157994 10880
rect 158670 9484 158730 10880
rect 159406 9756 159466 10880
rect 160142 8396 160202 10880
rect 160878 8396 160938 10880
rect 161614 8532 161674 10880
rect 162350 8396 162410 10880
rect 163086 8396 163146 10880
rect 163822 9756 163882 10880
rect 164558 8396 164618 10880
rect 165294 8396 165354 10880
rect 166030 8396 166090 10880
rect 166766 8260 166826 10880
rect 167502 8396 167562 10880
rect 168238 8124 168298 10880
rect 168974 9212 169034 10880
rect 171458 10300 171518 10880
rect 172194 10300 172254 10880
rect 172930 10300 172990 10880
rect 173666 10300 173726 10880
rect 174402 10300 174462 10880
rect 175138 10300 175198 10880
rect 175874 10300 175934 10880
rect 176610 10300 176670 10880
rect 177346 10300 177406 10880
rect 178082 10300 178142 10880
rect 178818 10300 178878 10880
rect 179554 10300 179614 10880
rect 180290 10300 180350 10880
rect 181026 10300 181086 10880
rect 181762 10436 181822 10880
rect 182498 10300 182558 10880
rect 183234 10300 183294 10880
rect 183970 10300 184030 10880
rect 184706 10300 184766 10880
rect 185442 10300 185502 10880
rect 186178 10300 186238 10880
rect 186914 10300 186974 10880
rect 187650 10300 187710 10880
rect 188386 10300 188446 10880
rect 189122 10300 189182 10880
rect 189858 10300 189918 10880
rect 190594 10436 190654 10880
rect 191330 10300 191390 10880
rect 192066 10300 192126 10880
rect 192802 10300 192862 10880
rect 193538 10436 193598 10880
rect 194274 10300 194334 10880
rect 195010 10300 195070 10880
rect 195746 10300 195806 10880
rect 196482 10300 196542 10880
rect 197218 10300 197278 10880
rect 197954 10300 198014 10880
rect 198690 10436 198750 10880
rect 199426 10300 199486 10880
rect 200162 10300 200222 10880
rect 200898 10436 200958 10880
rect 201634 10300 201694 10880
rect 202370 10436 202430 10880
rect 203106 10300 203166 10880
rect 99974 0 100034 444
rect 100710 0 100770 852
rect 103194 0 103254 444
rect 103930 0 103990 444
rect 104666 0 104726 444
rect 105402 0 105462 444
rect 106138 0 106198 444
rect 106874 0 106934 444
rect 107610 0 107670 444
rect 108346 0 108406 444
rect 109082 0 109142 444
rect 109818 0 109878 444
rect 110554 0 110614 444
rect 111290 0 111350 444
rect 112026 0 112086 444
rect 112762 0 112822 444
rect 113498 0 113558 308
rect 114234 0 114294 580
rect 114970 0 115030 580
rect 115706 0 115766 580
rect 116442 0 116502 580
rect 117178 0 117238 370
rect 117914 0 117974 580
rect 118650 0 118710 580
rect 119386 0 119446 580
rect 120122 0 120182 580
rect 120858 0 120918 580
rect 121594 0 121654 580
rect 122330 0 122390 580
rect 123066 0 123126 580
rect 123802 0 123862 580
rect 124538 0 124598 580
rect 125274 0 125334 580
rect 126010 0 126070 580
rect 126746 0 126806 580
rect 127482 0 127542 580
rect 128218 0 128278 370
rect 128954 0 129014 580
rect 129690 0 129750 580
rect 130426 0 130486 308
rect 131162 0 131222 580
rect 131898 0 131958 580
rect 132634 0 132694 580
rect 133370 0 133430 580
rect 134106 0 134166 580
rect 134842 0 134902 370
rect 137326 0 137386 1396
rect 138062 0 138122 580
rect 138798 0 138858 716
rect 139534 0 139594 444
rect 140270 0 140330 1260
rect 141006 0 141066 716
rect 141742 0 141802 580
rect 142478 0 142538 988
rect 143214 0 143274 716
rect 143950 0 144010 716
rect 144686 0 144746 1396
rect 145422 0 145482 716
rect 146158 0 146218 716
rect 146894 0 146954 716
rect 147630 0 147690 580
rect 148366 0 148426 716
rect 149102 0 149162 716
rect 149838 0 149898 988
rect 150574 0 150634 716
rect 151310 0 151370 716
rect 152046 0 152106 716
rect 152782 0 152842 716
rect 153518 0 153578 580
rect 154254 0 154314 716
rect 154990 0 155050 1260
rect 155726 0 155786 1396
rect 156462 0 156522 1396
rect 157198 0 157258 2756
rect 157934 0 157994 1396
rect 158670 0 158730 580
rect 159406 0 159466 2756
rect 160142 0 160202 1124
rect 160878 0 160938 580
rect 161614 0 161674 1124
rect 162350 0 162410 580
rect 163086 0 163146 1124
rect 163822 0 163882 1396
rect 164558 0 164618 580
rect 165294 0 165354 1124
rect 166030 0 166090 1124
rect 166766 0 166826 1124
rect 167502 0 167562 580
rect 168238 0 168298 1396
rect 169936 1040 170256 9840
rect 203734 1040 204054 9840
rect 205590 9620 205650 10880
rect 206326 10164 206386 10880
rect 207062 10164 207122 10880
rect 207798 10572 207858 10880
rect 208534 10164 208594 10880
rect 209270 10164 209330 10880
rect 210006 10436 210066 10880
rect 210742 10164 210802 10880
rect 211478 10436 211538 10880
rect 212214 6900 212274 10880
rect 212950 10164 213010 10880
rect 213686 10164 213746 10880
rect 214422 10164 214482 10880
rect 215158 10300 215218 10880
rect 215894 10164 215954 10880
rect 216630 9892 216690 10880
rect 217366 10164 217426 10880
rect 218102 10572 218162 10880
rect 218838 10164 218898 10880
rect 219574 10164 219634 10880
rect 220310 10300 220370 10880
rect 221046 10436 221106 10880
rect 221782 10300 221842 10880
rect 222518 10300 222578 10880
rect 223254 10164 223314 10880
rect 223990 9212 224050 10880
rect 224726 8396 224786 10880
rect 225462 9756 225522 10880
rect 226198 8668 226258 10880
rect 226934 8668 226994 10880
rect 227670 8668 227730 10880
rect 228406 9484 228466 10880
rect 229142 8668 229202 10880
rect 229878 9756 229938 10880
rect 230614 8396 230674 10880
rect 231350 9756 231410 10880
rect 232086 8668 232146 10880
rect 232822 8668 232882 10880
rect 233558 9756 233618 10880
rect 234294 9756 234354 10880
rect 235030 9756 235090 10880
rect 235766 9212 235826 10880
rect 236502 8668 236562 10880
rect 237238 9212 237298 10880
rect 239722 10300 239782 10880
rect 240458 10300 240518 10880
rect 241194 10300 241254 10880
rect 241930 10300 241990 10880
rect 242666 10300 242726 10880
rect 243402 10300 243462 10880
rect 244138 10300 244198 10880
rect 244874 10300 244934 10880
rect 245610 10300 245670 10880
rect 246346 10300 246406 10880
rect 247082 10300 247142 10880
rect 247818 10300 247878 10880
rect 248554 10300 248614 10880
rect 249290 10300 249350 10880
rect 250026 10300 250086 10880
rect 250762 10300 250822 10880
rect 251498 10300 251558 10880
rect 252234 10300 252294 10880
rect 252970 10300 253030 10880
rect 253706 10300 253766 10880
rect 254442 10300 254502 10880
rect 255178 10300 255238 10880
rect 255914 10300 255974 10880
rect 256650 10300 256710 10880
rect 257386 10300 257446 10880
rect 258122 10300 258182 10880
rect 258858 10300 258918 10880
rect 259594 10300 259654 10880
rect 260330 10300 260390 10880
rect 261066 10436 261126 10880
rect 261802 10300 261862 10880
rect 262538 10300 262598 10880
rect 263274 10300 263334 10880
rect 264010 10300 264070 10880
rect 264746 10436 264806 10880
rect 265482 10300 265542 10880
rect 266218 10510 266278 10880
rect 266954 10238 267014 10880
rect 267690 10238 267750 10880
rect 268426 10238 268486 10880
rect 269162 10238 269222 10880
rect 269898 10238 269958 10880
rect 270634 10238 270694 10880
rect 271370 10238 271430 10880
rect 168974 0 169034 580
rect 171458 0 171518 370
rect 172194 0 172254 370
rect 172930 0 172990 370
rect 173666 0 173726 370
rect 174402 0 174462 370
rect 175138 0 175198 370
rect 175874 0 175934 370
rect 176610 0 176670 370
rect 177346 0 177406 370
rect 178082 0 178142 370
rect 178818 0 178878 370
rect 179554 0 179614 370
rect 180290 0 180350 370
rect 181026 0 181086 370
rect 181762 0 181822 370
rect 182498 0 182558 370
rect 183234 0 183294 370
rect 183970 0 184030 370
rect 184706 0 184766 370
rect 185442 0 185502 370
rect 186178 0 186238 370
rect 186914 0 186974 370
rect 187650 0 187710 370
rect 188386 0 188446 370
rect 189122 0 189182 370
rect 189858 0 189918 370
rect 190594 0 190654 370
rect 191330 0 191390 370
rect 192066 0 192126 370
rect 192802 0 192862 370
rect 193538 0 193598 370
rect 194274 0 194334 370
rect 195010 0 195070 370
rect 195746 0 195806 370
rect 196482 0 196542 370
rect 197218 0 197278 370
rect 197954 0 198014 370
rect 198690 0 198750 370
rect 199426 0 199486 370
rect 200162 0 200222 370
rect 200898 0 200958 370
rect 201634 0 201694 370
rect 202370 0 202430 370
rect 203106 0 203166 370
rect 205590 0 205650 370
rect 206326 0 206386 852
rect 207062 0 207122 852
rect 207798 0 207858 852
rect 208534 0 208594 852
rect 209270 0 209330 852
rect 210006 0 210066 988
rect 210742 0 210802 1260
rect 211478 0 211538 988
rect 212214 0 212274 852
rect 212950 0 213010 852
rect 213686 0 213746 852
rect 214422 0 214482 852
rect 215158 0 215218 852
rect 215894 0 215954 852
rect 216630 0 216690 1396
rect 217366 0 217426 852
rect 218102 0 218162 852
rect 218838 0 218898 308
rect 219574 0 219634 308
rect 220310 0 220370 1396
rect 221046 0 221106 852
rect 221782 0 221842 308
rect 222518 0 222578 1260
rect 223254 0 223314 2756
rect 223990 0 224050 1396
rect 224726 0 224786 2756
rect 225462 0 225522 1396
rect 226198 0 226258 2756
rect 226934 0 226994 1260
rect 227670 0 227730 1260
rect 228406 0 228466 1124
rect 229142 0 229202 308
rect 229878 0 229938 308
rect 230614 0 230674 308
rect 231350 0 231410 1124
rect 232086 0 232146 1124
rect 232822 0 232882 1124
rect 233558 0 233618 308
rect 234294 0 234354 308
rect 235030 0 235090 444
rect 235766 0 235826 2756
rect 236502 0 236562 1124
rect 237238 0 237298 1396
rect 237533 1040 237853 9840
rect 271331 1040 271651 9840
rect 239722 0 239782 308
rect 240458 0 240518 308
rect 241194 0 241254 444
rect 241930 0 241990 444
rect 242666 0 242726 370
rect 243402 0 243462 444
rect 244138 0 244198 370
rect 244874 0 244934 444
rect 245610 0 245670 444
rect 246346 0 246406 444
rect 247082 0 247142 370
rect 247818 0 247878 370
rect 248554 0 248614 444
rect 249290 0 249350 370
rect 250026 0 250086 580
rect 250762 0 250822 370
rect 251498 0 251558 580
rect 252234 0 252294 580
rect 252970 0 253030 580
rect 253706 0 253766 580
rect 254442 0 254502 308
rect 255178 0 255238 580
rect 255914 0 255974 580
rect 256650 0 256710 580
rect 257386 0 257446 580
rect 258122 0 258182 642
rect 258858 0 258918 580
rect 259594 0 259654 580
rect 260330 0 260390 580
rect 261066 0 261126 580
rect 261802 0 261862 444
rect 262538 0 262598 580
rect 263274 0 263334 580
rect 264010 0 264070 580
rect 264746 0 264806 370
rect 265482 0 265542 580
rect 266218 0 266278 580
rect 266954 0 267014 580
rect 267690 0 267750 580
rect 268426 0 268486 580
rect 269162 0 269222 444
rect 269898 0 269958 580
rect 270634 0 270694 370
rect 271370 0 271430 308
<< obsm4 >>
rect 938 10084 1454 10573
rect 1674 10084 2190 10573
rect 2410 10084 2926 10573
rect 938 9812 2926 10084
rect 3146 10084 3662 10573
rect 3882 10084 4398 10573
rect 4618 10084 5134 10573
rect 5354 10084 5870 10573
rect 6090 10084 6606 10573
rect 6826 10084 7342 10573
rect 7562 10084 8078 10573
rect 3146 9812 8078 10084
rect 8298 10084 8814 10573
rect 9034 10492 9550 10573
rect 9770 10492 10286 10573
rect 9034 10084 10286 10492
rect 8298 9812 10286 10084
rect 10506 9812 11022 10573
rect 11242 10084 11758 10573
rect 11978 10084 12494 10573
rect 12714 10084 13230 10573
rect 11242 9812 13230 10084
rect 13450 10084 13966 10573
rect 14186 10084 14702 10573
rect 14922 10084 15438 10573
rect 15658 10084 16174 10573
rect 16394 10084 16910 10573
rect 17130 10084 17646 10573
rect 17866 10084 18382 10573
rect 18602 10084 19118 10573
rect 13450 9812 19118 10084
rect 938 9132 19118 9812
rect 795 6820 19118 9132
rect 19338 6820 19854 10573
rect 20074 10492 20590 10573
rect 20810 10492 21326 10573
rect 20074 9812 21326 10492
rect 21546 10084 22062 10573
rect 22282 10084 22798 10573
rect 21546 9812 22798 10084
rect 20074 6820 22798 9812
rect 23018 6820 23534 10573
rect 23754 8588 24270 10573
rect 24490 8588 25006 10573
rect 23754 6820 25006 8588
rect 25226 9540 25742 10573
rect 25962 9540 26478 10573
rect 25226 8316 26478 9540
rect 26698 8316 27214 10573
rect 25226 7772 27214 8316
rect 27434 8316 27950 10573
rect 28170 9404 28686 10573
rect 28906 9404 29422 10573
rect 28170 8588 29422 9404
rect 29642 8588 30158 10573
rect 30378 8588 30894 10573
rect 31114 10220 31630 10573
rect 31850 10220 32366 10573
rect 31114 9540 32366 10220
rect 32586 10220 34850 10573
rect 35070 10220 35586 10573
rect 35806 10220 36322 10573
rect 36542 10220 37058 10573
rect 37278 10220 37794 10573
rect 38014 10220 38530 10573
rect 38750 10220 39266 10573
rect 39486 10220 40002 10573
rect 40222 10220 40738 10573
rect 40958 10220 41474 10573
rect 41694 10220 42210 10573
rect 42430 10220 42946 10573
rect 43166 10220 43682 10573
rect 43902 10220 44418 10573
rect 44638 10220 45154 10573
rect 45374 10220 45890 10573
rect 46110 10220 46626 10573
rect 46846 10220 47362 10573
rect 47582 10220 48098 10573
rect 48318 10220 48834 10573
rect 49054 10220 49570 10573
rect 49790 10220 50306 10573
rect 50526 10220 51042 10573
rect 51262 10220 51778 10573
rect 51998 10220 52514 10573
rect 52734 10220 53250 10573
rect 53470 10356 53986 10573
rect 54206 10356 54722 10573
rect 53470 10220 54722 10356
rect 54942 10220 55458 10573
rect 55678 10220 56194 10573
rect 56414 10220 56930 10573
rect 57150 10220 57666 10573
rect 57886 10220 58402 10573
rect 58622 10220 59138 10573
rect 59358 10220 59874 10573
rect 60094 10220 60610 10573
rect 60830 10220 61346 10573
rect 61566 10220 62082 10573
rect 62302 10220 62818 10573
rect 63038 10220 63554 10573
rect 63774 10220 64290 10573
rect 64510 10220 65026 10573
rect 65246 10220 65762 10573
rect 65982 10220 66498 10573
rect 66718 10220 68982 10573
rect 32586 9920 68982 10220
rect 32586 9540 34662 9920
rect 31114 8588 34662 9540
rect 28170 8316 34662 8588
rect 27434 7772 34662 8316
rect 25226 6820 34662 7772
rect 795 3380 34662 6820
rect 795 2972 24270 3380
rect 795 1476 19118 2972
rect 938 1340 16174 1476
rect 938 307 1454 1340
rect 1674 1068 16174 1340
rect 1674 307 2190 1068
rect 2410 796 4398 1068
rect 2410 307 2926 796
rect 3146 660 4398 796
rect 3146 307 3662 660
rect 3882 307 4398 660
rect 4618 796 6606 1068
rect 4618 307 5134 796
rect 5354 307 5870 796
rect 6090 307 6606 796
rect 6826 796 13966 1068
rect 6826 307 7342 796
rect 7562 660 8814 796
rect 7562 307 8078 660
rect 8298 307 8814 660
rect 9034 660 13966 796
rect 9034 307 9550 660
rect 9770 307 10286 660
rect 10506 307 11022 660
rect 11242 307 11758 660
rect 11978 307 12494 660
rect 12714 307 13230 660
rect 13450 307 13966 660
rect 14186 796 16174 1068
rect 14186 307 14702 796
rect 14922 307 15438 796
rect 15658 307 16174 796
rect 16394 660 19118 1476
rect 16394 307 16910 660
rect 17130 307 17646 660
rect 17866 307 18382 660
rect 18602 307 19118 660
rect 19338 2836 22798 2972
rect 19338 307 19854 2836
rect 20074 1748 22062 2836
rect 20074 1476 21326 1748
rect 20074 307 20590 1476
rect 20810 307 21326 1476
rect 21546 307 22062 1748
rect 22282 307 22798 2836
rect 23018 660 24270 2972
rect 23018 307 23534 660
rect 23754 307 24270 660
rect 24490 2836 34662 3380
rect 24490 307 25006 2836
rect 25226 1476 34662 2836
rect 25226 1340 32366 1476
rect 25226 307 25742 1340
rect 25962 307 26478 1340
rect 26698 307 27214 1340
rect 27434 660 32366 1340
rect 27434 524 28686 660
rect 27434 307 27950 524
rect 28170 307 28686 524
rect 28906 524 30158 660
rect 28906 307 29422 524
rect 29642 307 30158 524
rect 30378 524 32366 660
rect 30378 388 31630 524
rect 30378 307 30894 388
rect 31114 307 31630 388
rect 31850 307 32366 524
rect 32586 960 34662 1476
rect 35142 960 68460 9920
rect 68940 9540 68982 9920
rect 69202 9540 69718 10573
rect 68940 8996 69718 9540
rect 69938 9540 70454 10573
rect 70674 10492 71190 10573
rect 71410 10492 71926 10573
rect 70674 10356 71926 10492
rect 72146 10356 72662 10573
rect 70674 9540 72662 10356
rect 72882 9540 73398 10573
rect 69938 8996 73398 9540
rect 73618 10492 74134 10573
rect 74354 10492 74870 10573
rect 73618 8996 74870 10492
rect 75090 9540 75606 10573
rect 75826 9676 76342 10573
rect 76562 10356 77078 10573
rect 77298 10356 77814 10573
rect 76562 9676 77814 10356
rect 75826 9540 77814 9676
rect 78034 9540 78550 10573
rect 75090 8996 78550 9540
rect 78770 9676 79286 10573
rect 79506 9676 80022 10573
rect 78770 8996 80022 9676
rect 80242 9540 80758 10573
rect 80978 9676 81494 10573
rect 81714 10356 82230 10573
rect 82450 10356 82966 10573
rect 81714 9676 82966 10356
rect 80978 9540 82966 9676
rect 83186 10356 83702 10573
rect 83922 10492 84438 10573
rect 84658 10492 85174 10573
rect 83922 10356 85174 10492
rect 83186 9812 85174 10356
rect 85394 9812 85910 10573
rect 86130 10492 86646 10573
rect 86866 10492 87382 10573
rect 86130 9812 87382 10492
rect 83186 9540 87382 9812
rect 80242 8996 87382 9540
rect 68940 8588 87382 8996
rect 87602 9132 88118 10573
rect 88338 9132 88854 10573
rect 87602 8588 88854 9132
rect 68940 8044 88854 8588
rect 89074 10220 89590 10573
rect 89810 10220 90326 10573
rect 89074 8588 90326 10220
rect 90546 8724 91062 10573
rect 91282 8724 91798 10573
rect 90546 8588 91798 8724
rect 92018 8588 92534 10573
rect 89074 8316 92534 8588
rect 92754 9676 93270 10573
rect 93490 9676 94006 10573
rect 92754 8588 94006 9676
rect 94226 8588 94742 10573
rect 94962 9676 95478 10573
rect 95698 9676 96214 10573
rect 96434 9676 96950 10573
rect 94962 8588 96950 9676
rect 97170 9676 97686 10573
rect 97906 9676 98422 10573
rect 97170 8588 98422 9676
rect 98642 8588 99158 10573
rect 92754 8316 99158 8588
rect 89074 8180 99158 8316
rect 99378 8588 99894 10573
rect 100114 9676 100630 10573
rect 100850 10220 103114 10573
rect 103334 10220 103850 10573
rect 104070 10220 104586 10573
rect 104806 10220 105322 10573
rect 105542 10220 106058 10573
rect 106278 10220 106794 10573
rect 107014 10220 107530 10573
rect 107750 10220 108266 10573
rect 108486 10220 109002 10573
rect 109222 10220 109738 10573
rect 109958 10220 110474 10573
rect 110694 10220 111210 10573
rect 111430 10220 111946 10573
rect 112166 10220 112682 10573
rect 112902 10220 113418 10573
rect 113638 10220 114154 10573
rect 114374 10220 114890 10573
rect 115110 10220 115626 10573
rect 115846 10220 116362 10573
rect 116582 10220 117098 10573
rect 117318 10220 117834 10573
rect 118054 10220 118570 10573
rect 118790 10220 119306 10573
rect 119526 10220 120042 10573
rect 120262 10220 120778 10573
rect 120998 10220 121514 10573
rect 121734 10220 122250 10573
rect 122470 10220 122986 10573
rect 123206 10220 123722 10573
rect 123942 10220 124458 10573
rect 124678 10356 125194 10573
rect 125414 10356 125930 10573
rect 124678 10220 125930 10356
rect 126150 10220 126666 10573
rect 126886 10220 127402 10573
rect 127622 10356 128138 10573
rect 128358 10356 128874 10573
rect 127622 10220 128874 10356
rect 129094 10220 129610 10573
rect 129830 10220 130346 10573
rect 130566 10220 131082 10573
rect 131302 10220 131818 10573
rect 132038 10220 132554 10573
rect 132774 10220 133290 10573
rect 133510 10220 134026 10573
rect 134246 10220 134762 10573
rect 134982 10220 137246 10573
rect 100850 9920 137246 10220
rect 100850 9676 102259 9920
rect 100114 8588 102259 9676
rect 99378 8180 102259 8588
rect 89074 8044 102259 8180
rect 68940 1612 102259 8044
rect 68940 1340 80022 1612
rect 68940 1068 71190 1340
rect 68940 960 70454 1068
rect 32586 796 70454 960
rect 32586 660 68982 796
rect 32586 388 35586 660
rect 32586 307 34850 388
rect 35070 307 35586 388
rect 35806 307 36322 660
rect 36542 307 37058 660
rect 37278 307 37794 660
rect 38014 307 38530 660
rect 38750 388 40002 660
rect 38750 307 39266 388
rect 39486 307 40002 388
rect 40222 307 40738 660
rect 40958 307 41474 660
rect 41694 307 42210 660
rect 42430 307 42946 660
rect 43166 307 43682 660
rect 43902 307 44418 660
rect 44638 307 45154 660
rect 45374 307 45890 660
rect 46110 307 46626 660
rect 46846 307 47362 660
rect 47582 307 48098 660
rect 48318 307 48834 660
rect 49054 307 49570 660
rect 49790 307 50306 660
rect 50526 307 51042 660
rect 51262 307 51778 660
rect 51998 307 52514 660
rect 52734 307 53250 660
rect 53470 450 54722 660
rect 53470 307 53986 450
rect 54206 307 54722 450
rect 54942 307 55458 660
rect 55678 307 56194 660
rect 56414 307 56930 660
rect 57150 307 57666 660
rect 57886 307 58402 660
rect 58622 450 60610 660
rect 58622 307 59138 450
rect 59358 307 59874 450
rect 60094 307 60610 450
rect 60830 307 61346 660
rect 61566 307 62082 660
rect 62302 307 62818 660
rect 63038 307 63554 660
rect 63774 307 64290 660
rect 64510 307 65026 660
rect 65246 524 68982 660
rect 65246 307 65762 524
rect 65982 307 66498 524
rect 66718 307 68982 524
rect 69202 307 69718 796
rect 69938 307 70454 796
rect 70674 307 71190 1068
rect 71410 1068 73398 1340
rect 71410 307 71926 1068
rect 72146 660 73398 1068
rect 72146 307 72662 660
rect 72882 307 73398 660
rect 73618 1068 76342 1340
rect 73618 307 74134 1068
rect 74354 660 75606 1068
rect 74354 307 74870 660
rect 75090 307 75606 660
rect 75826 307 76342 1068
rect 76562 1068 77814 1340
rect 76562 307 77078 1068
rect 77298 307 77814 1068
rect 78034 796 79286 1340
rect 78034 307 78550 796
rect 78770 307 79286 796
rect 79506 307 80022 1340
rect 80242 796 81494 1612
rect 80242 307 80758 796
rect 80978 307 81494 796
rect 81714 1340 82966 1612
rect 81714 307 82230 1340
rect 82450 307 82966 1340
rect 83186 307 83702 1612
rect 83922 1340 99158 1612
rect 83922 1068 87382 1340
rect 83922 796 85910 1068
rect 83922 307 84438 796
rect 84658 307 85174 796
rect 85394 307 85910 796
rect 86130 796 87382 1068
rect 86130 307 86646 796
rect 86866 307 87382 796
rect 87602 1204 88854 1340
rect 87602 307 88118 1204
rect 88338 307 88854 1204
rect 89074 1204 99158 1340
rect 89074 796 94006 1204
rect 89074 388 90326 796
rect 89074 307 89590 388
rect 89810 307 90326 388
rect 90546 388 91798 796
rect 90546 307 91062 388
rect 91282 307 91798 388
rect 92018 388 93270 796
rect 92018 307 92534 388
rect 92754 307 93270 388
rect 93490 307 94006 796
rect 94226 307 94742 1204
rect 94962 307 95478 1204
rect 95698 307 96214 1204
rect 96434 796 99158 1204
rect 96434 524 97686 796
rect 96434 307 96950 524
rect 97170 307 97686 524
rect 97906 307 98422 796
rect 98642 307 99158 796
rect 99378 960 102259 1612
rect 102739 960 136057 9920
rect 136537 9540 137246 9920
rect 137466 10220 137982 10573
rect 138202 10220 138718 10573
rect 137466 10084 138718 10220
rect 138938 10084 139454 10573
rect 137466 9812 139454 10084
rect 139674 10084 140190 10573
rect 140410 10084 140926 10573
rect 141146 10084 141662 10573
rect 141882 10220 142398 10573
rect 142618 10220 143134 10573
rect 141882 10084 143134 10220
rect 143354 10084 143870 10573
rect 144090 10084 144606 10573
rect 139674 9812 144606 10084
rect 144826 10084 145342 10573
rect 145562 10084 146078 10573
rect 146298 10084 146814 10573
rect 147034 10356 147550 10573
rect 147770 10356 148286 10573
rect 147034 10084 148286 10356
rect 148506 10084 149022 10573
rect 149242 10084 149758 10573
rect 144826 9812 149758 10084
rect 149978 10084 150494 10573
rect 150714 10084 151230 10573
rect 151450 10084 151966 10573
rect 152186 10084 152702 10573
rect 152922 10220 153438 10573
rect 153658 10220 154174 10573
rect 152922 10084 154174 10220
rect 154394 10084 154910 10573
rect 149978 9812 154910 10084
rect 155130 9812 155646 10573
rect 137466 9676 155646 9812
rect 155866 9676 156382 10573
rect 156602 10220 157118 10573
rect 157338 10220 157854 10573
rect 156602 9676 157854 10220
rect 158074 9676 158590 10573
rect 137466 9540 158590 9676
rect 136537 9404 158590 9540
rect 158810 9676 159326 10573
rect 159546 9676 160062 10573
rect 158810 9404 160062 9676
rect 136537 8316 160062 9404
rect 160282 8316 160798 10573
rect 161018 8452 161534 10573
rect 161754 8452 162270 10573
rect 161018 8316 162270 8452
rect 162490 8316 163006 10573
rect 163226 9676 163742 10573
rect 163962 9676 164478 10573
rect 163226 8316 164478 9676
rect 164698 8316 165214 10573
rect 165434 8316 165950 10573
rect 166170 8316 166686 10573
rect 136537 8180 166686 8316
rect 166906 8316 167422 10573
rect 167642 8316 168158 10573
rect 166906 8180 168158 8316
rect 136537 8044 168158 8180
rect 168378 9132 168894 10573
rect 169114 10220 171378 10573
rect 171598 10220 172114 10573
rect 172334 10220 172850 10573
rect 173070 10220 173586 10573
rect 173806 10220 174322 10573
rect 174542 10220 175058 10573
rect 175278 10220 175794 10573
rect 176014 10220 176530 10573
rect 176750 10220 177266 10573
rect 177486 10220 178002 10573
rect 178222 10220 178738 10573
rect 178958 10220 179474 10573
rect 179694 10220 180210 10573
rect 180430 10220 180946 10573
rect 181166 10356 181682 10573
rect 181902 10356 182418 10573
rect 181166 10220 182418 10356
rect 182638 10220 183154 10573
rect 183374 10220 183890 10573
rect 184110 10220 184626 10573
rect 184846 10220 185362 10573
rect 185582 10220 186098 10573
rect 186318 10220 186834 10573
rect 187054 10220 187570 10573
rect 187790 10220 188306 10573
rect 188526 10220 189042 10573
rect 189262 10220 189778 10573
rect 189998 10356 190514 10573
rect 190734 10356 191250 10573
rect 189998 10220 191250 10356
rect 191470 10220 191986 10573
rect 192206 10220 192722 10573
rect 192942 10356 193458 10573
rect 193678 10356 194194 10573
rect 192942 10220 194194 10356
rect 194414 10220 194930 10573
rect 195150 10220 195666 10573
rect 195886 10220 196402 10573
rect 196622 10220 197138 10573
rect 197358 10220 197874 10573
rect 198094 10356 198610 10573
rect 198830 10356 199346 10573
rect 198094 10220 199346 10356
rect 199566 10220 200082 10573
rect 200302 10356 200818 10573
rect 201038 10356 201554 10573
rect 200302 10220 201554 10356
rect 201774 10356 202290 10573
rect 202510 10356 203026 10573
rect 201774 10220 203026 10356
rect 203246 10220 205510 10573
rect 169114 9920 205510 10220
rect 169114 9132 169856 9920
rect 168378 8044 169856 9132
rect 136537 2836 169856 8044
rect 136537 1476 157118 2836
rect 136537 960 137246 1476
rect 99378 932 137246 960
rect 99378 524 100630 932
rect 99378 307 99894 524
rect 100114 307 100630 524
rect 100850 660 137246 932
rect 100850 524 114154 660
rect 100850 307 103114 524
rect 103334 307 103850 524
rect 104070 307 104586 524
rect 104806 307 105322 524
rect 105542 307 106058 524
rect 106278 307 106794 524
rect 107014 307 107530 524
rect 107750 307 108266 524
rect 108486 307 109002 524
rect 109222 307 109738 524
rect 109958 307 110474 524
rect 110694 307 111210 524
rect 111430 307 111946 524
rect 112166 307 112682 524
rect 112902 388 114154 524
rect 112902 307 113418 388
rect 113638 307 114154 388
rect 114374 307 114890 660
rect 115110 307 115626 660
rect 115846 307 116362 660
rect 116582 450 117834 660
rect 116582 307 117098 450
rect 117318 307 117834 450
rect 118054 307 118570 660
rect 118790 307 119306 660
rect 119526 307 120042 660
rect 120262 307 120778 660
rect 120998 307 121514 660
rect 121734 307 122250 660
rect 122470 307 122986 660
rect 123206 307 123722 660
rect 123942 307 124458 660
rect 124678 307 125194 660
rect 125414 307 125930 660
rect 126150 307 126666 660
rect 126886 307 127402 660
rect 127622 450 128874 660
rect 127622 307 128138 450
rect 128358 307 128874 450
rect 129094 307 129610 660
rect 129830 388 131082 660
rect 129830 307 130346 388
rect 130566 307 131082 388
rect 131302 307 131818 660
rect 132038 307 132554 660
rect 132774 307 133290 660
rect 133510 307 134026 660
rect 134246 450 137246 660
rect 134246 307 134762 450
rect 134982 307 137246 450
rect 137466 1340 144606 1476
rect 137466 796 140190 1340
rect 137466 660 138718 796
rect 137466 307 137982 660
rect 138202 307 138718 660
rect 138938 524 140190 796
rect 138938 307 139454 524
rect 139674 307 140190 524
rect 140410 1068 144606 1340
rect 140410 796 142398 1068
rect 140410 307 140926 796
rect 141146 660 142398 796
rect 141146 307 141662 660
rect 141882 307 142398 660
rect 142618 796 144606 1068
rect 142618 307 143134 796
rect 143354 307 143870 796
rect 144090 307 144606 796
rect 144826 1340 155646 1476
rect 144826 1068 154910 1340
rect 144826 796 149758 1068
rect 144826 307 145342 796
rect 145562 307 146078 796
rect 146298 307 146814 796
rect 147034 660 148286 796
rect 147034 307 147550 660
rect 147770 307 148286 660
rect 148506 307 149022 796
rect 149242 307 149758 796
rect 149978 796 154910 1068
rect 149978 307 150494 796
rect 150714 307 151230 796
rect 151450 307 151966 796
rect 152186 307 152702 796
rect 152922 660 154174 796
rect 152922 307 153438 660
rect 153658 307 154174 660
rect 154394 307 154910 796
rect 155130 307 155646 1340
rect 155866 307 156382 1476
rect 156602 307 157118 1476
rect 157338 1476 159326 2836
rect 157338 307 157854 1476
rect 158074 660 159326 1476
rect 158074 307 158590 660
rect 158810 307 159326 660
rect 159546 1476 169856 2836
rect 159546 1204 163742 1476
rect 159546 307 160062 1204
rect 160282 660 161534 1204
rect 160282 307 160798 660
rect 161018 307 161534 660
rect 161754 660 163006 1204
rect 161754 307 162270 660
rect 162490 307 163006 660
rect 163226 307 163742 1204
rect 163962 1204 168158 1476
rect 163962 660 165214 1204
rect 163962 307 164478 660
rect 164698 307 165214 660
rect 165434 307 165950 1204
rect 166170 307 166686 1204
rect 166906 660 168158 1204
rect 166906 307 167422 660
rect 167642 307 168158 660
rect 168378 960 169856 1476
rect 170336 960 203654 9920
rect 204134 9540 205510 9920
rect 205730 10084 206246 10573
rect 206466 10084 206982 10573
rect 207202 10492 207718 10573
rect 207938 10492 208454 10573
rect 207202 10084 208454 10492
rect 208674 10084 209190 10573
rect 209410 10356 209926 10573
rect 210146 10356 210662 10573
rect 209410 10084 210662 10356
rect 210882 10356 211398 10573
rect 211618 10356 212134 10573
rect 210882 10084 212134 10356
rect 205730 9540 212134 10084
rect 204134 6820 212134 9540
rect 212354 10084 212870 10573
rect 213090 10084 213606 10573
rect 213826 10084 214342 10573
rect 214562 10220 215078 10573
rect 215298 10220 215814 10573
rect 214562 10084 215814 10220
rect 216034 10084 216550 10573
rect 212354 9812 216550 10084
rect 216770 10084 217286 10573
rect 217506 10492 218022 10573
rect 218242 10492 218758 10573
rect 217506 10084 218758 10492
rect 218978 10084 219494 10573
rect 219714 10220 220230 10573
rect 220450 10356 220966 10573
rect 221186 10356 221702 10573
rect 220450 10220 221702 10356
rect 221922 10220 222438 10573
rect 222658 10220 223174 10573
rect 219714 10084 223174 10220
rect 223394 10084 223910 10573
rect 216770 9812 223910 10084
rect 212354 9132 223910 9812
rect 224130 9132 224646 10573
rect 212354 8316 224646 9132
rect 224866 9676 225382 10573
rect 225602 9676 226118 10573
rect 224866 8588 226118 9676
rect 226338 8588 226854 10573
rect 227074 8588 227590 10573
rect 227810 9404 228326 10573
rect 228546 9404 229062 10573
rect 227810 8588 229062 9404
rect 229282 9676 229798 10573
rect 230018 9676 230534 10573
rect 229282 8588 230534 9676
rect 224866 8316 230534 8588
rect 230754 9676 231270 10573
rect 231490 9676 232006 10573
rect 230754 8588 232006 9676
rect 232226 8588 232742 10573
rect 232962 9676 233478 10573
rect 233698 9676 234214 10573
rect 234434 9676 234950 10573
rect 235170 9676 235686 10573
rect 232962 9132 235686 9676
rect 235906 9132 236422 10573
rect 232962 8588 236422 9132
rect 236642 9132 237158 10573
rect 237378 10220 239642 10573
rect 239862 10220 240378 10573
rect 240598 10220 241114 10573
rect 241334 10220 241850 10573
rect 242070 10220 242586 10573
rect 242806 10220 243322 10573
rect 243542 10220 244058 10573
rect 244278 10220 244794 10573
rect 245014 10220 245530 10573
rect 245750 10220 246266 10573
rect 246486 10220 247002 10573
rect 247222 10220 247738 10573
rect 247958 10220 248474 10573
rect 248694 10220 249210 10573
rect 249430 10220 249946 10573
rect 250166 10220 250682 10573
rect 250902 10220 251418 10573
rect 251638 10220 252154 10573
rect 252374 10220 252890 10573
rect 253110 10220 253626 10573
rect 253846 10220 254362 10573
rect 254582 10220 255098 10573
rect 255318 10220 255834 10573
rect 256054 10220 256570 10573
rect 256790 10220 257306 10573
rect 257526 10220 258042 10573
rect 258262 10220 258778 10573
rect 258998 10220 259514 10573
rect 259734 10220 260250 10573
rect 260470 10356 260986 10573
rect 261206 10356 261722 10573
rect 260470 10220 261722 10356
rect 261942 10220 262458 10573
rect 262678 10220 263194 10573
rect 263414 10220 263930 10573
rect 264150 10356 264666 10573
rect 264886 10356 265402 10573
rect 264150 10220 265402 10356
rect 265622 10430 266138 10573
rect 266358 10430 266874 10573
rect 265622 10220 266874 10430
rect 237378 10158 266874 10220
rect 267094 10158 267610 10573
rect 267830 10158 268346 10573
rect 268566 10158 269082 10573
rect 269302 10158 269818 10573
rect 270038 10158 270554 10573
rect 270774 10158 271290 10573
rect 237378 9920 271433 10158
rect 237378 9132 237453 9920
rect 236642 8588 237453 9132
rect 230754 8316 237453 8588
rect 212354 6820 237453 8316
rect 204134 2836 237453 6820
rect 204134 1476 223174 2836
rect 204134 1340 216550 1476
rect 204134 1068 210662 1340
rect 204134 960 209926 1068
rect 168378 932 209926 960
rect 168378 660 206246 932
rect 168378 307 168894 660
rect 169114 450 206246 660
rect 169114 307 171378 450
rect 171598 307 172114 450
rect 172334 307 172850 450
rect 173070 307 173586 450
rect 173806 307 174322 450
rect 174542 307 175058 450
rect 175278 307 175794 450
rect 176014 307 176530 450
rect 176750 307 177266 450
rect 177486 307 178002 450
rect 178222 307 178738 450
rect 178958 307 179474 450
rect 179694 307 180210 450
rect 180430 307 180946 450
rect 181166 307 181682 450
rect 181902 307 182418 450
rect 182638 307 183154 450
rect 183374 307 183890 450
rect 184110 307 184626 450
rect 184846 307 185362 450
rect 185582 307 186098 450
rect 186318 307 186834 450
rect 187054 307 187570 450
rect 187790 307 188306 450
rect 188526 307 189042 450
rect 189262 307 189778 450
rect 189998 307 190514 450
rect 190734 307 191250 450
rect 191470 307 191986 450
rect 192206 307 192722 450
rect 192942 307 193458 450
rect 193678 307 194194 450
rect 194414 307 194930 450
rect 195150 307 195666 450
rect 195886 307 196402 450
rect 196622 307 197138 450
rect 197358 307 197874 450
rect 198094 307 198610 450
rect 198830 307 199346 450
rect 199566 307 200082 450
rect 200302 307 200818 450
rect 201038 307 201554 450
rect 201774 307 202290 450
rect 202510 307 203026 450
rect 203246 307 205510 450
rect 205730 307 206246 450
rect 206466 307 206982 932
rect 207202 307 207718 932
rect 207938 307 208454 932
rect 208674 307 209190 932
rect 209410 307 209926 932
rect 210146 307 210662 1068
rect 210882 1068 216550 1340
rect 210882 307 211398 1068
rect 211618 932 216550 1068
rect 211618 307 212134 932
rect 212354 307 212870 932
rect 213090 307 213606 932
rect 213826 307 214342 932
rect 214562 307 215078 932
rect 215298 307 215814 932
rect 216034 307 216550 932
rect 216770 932 220230 1476
rect 216770 307 217286 932
rect 217506 307 218022 932
rect 218242 388 220230 932
rect 218242 307 218758 388
rect 218978 307 219494 388
rect 219714 307 220230 388
rect 220450 1340 223174 1476
rect 220450 932 222438 1340
rect 220450 307 220966 932
rect 221186 388 222438 932
rect 221186 307 221702 388
rect 221922 307 222438 388
rect 222658 307 223174 1340
rect 223394 1476 224646 2836
rect 223394 307 223910 1476
rect 224130 307 224646 1476
rect 224866 1476 226118 2836
rect 224866 307 225382 1476
rect 225602 307 226118 1476
rect 226338 1340 235686 2836
rect 226338 307 226854 1340
rect 227074 307 227590 1340
rect 227810 1204 235686 1340
rect 227810 307 228326 1204
rect 228546 388 231270 1204
rect 228546 307 229062 388
rect 229282 307 229798 388
rect 230018 307 230534 388
rect 230754 307 231270 388
rect 231490 307 232006 1204
rect 232226 307 232742 1204
rect 232962 524 235686 1204
rect 232962 388 234950 524
rect 232962 307 233478 388
rect 233698 307 234214 388
rect 234434 307 234950 388
rect 235170 307 235686 524
rect 235906 1476 237453 2836
rect 235906 1204 237158 1476
rect 235906 307 236422 1204
rect 236642 307 237158 1204
rect 237378 960 237453 1476
rect 237933 960 271251 9920
rect 237378 722 271433 960
rect 237378 660 258042 722
rect 237378 524 249946 660
rect 237378 388 241114 524
rect 237378 307 239642 388
rect 239862 307 240378 388
rect 240598 307 241114 388
rect 241334 307 241850 524
rect 242070 450 243322 524
rect 242070 307 242586 450
rect 242806 307 243322 450
rect 243542 450 244794 524
rect 243542 307 244058 450
rect 244278 307 244794 450
rect 245014 307 245530 524
rect 245750 307 246266 524
rect 246486 450 248474 524
rect 246486 307 247002 450
rect 247222 307 247738 450
rect 247958 307 248474 450
rect 248694 450 249946 524
rect 248694 307 249210 450
rect 249430 307 249946 450
rect 250166 450 251418 660
rect 250166 307 250682 450
rect 250902 307 251418 450
rect 251638 307 252154 660
rect 252374 307 252890 660
rect 253110 307 253626 660
rect 253846 388 255098 660
rect 253846 307 254362 388
rect 254582 307 255098 388
rect 255318 307 255834 660
rect 256054 307 256570 660
rect 256790 307 257306 660
rect 257526 307 258042 660
rect 258262 660 271433 722
rect 258262 307 258778 660
rect 258998 307 259514 660
rect 259734 307 260250 660
rect 260470 307 260986 660
rect 261206 524 262458 660
rect 261206 307 261722 524
rect 261942 307 262458 524
rect 262678 307 263194 660
rect 263414 307 263930 660
rect 264150 450 265402 660
rect 264150 307 264666 450
rect 264886 307 265402 450
rect 265622 307 266138 660
rect 266358 307 266874 660
rect 267094 307 267610 660
rect 267830 307 268346 660
rect 268566 524 269818 660
rect 268566 307 269082 524
rect 269302 307 269818 524
rect 270038 450 271433 660
rect 270038 307 270554 450
rect 270774 388 271433 450
rect 270774 307 271290 388
<< labels >>
rlabel metal3 s 272198 9558 272504 9618 6 addr[0]
port 1 nsew signal input
rlabel metal3 s 272014 9422 272504 9482 6 addr[1]
port 2 nsew signal input
rlabel metal3 s 268990 9286 272504 9346 6 addr[2]
port 3 nsew signal input
rlabel metal3 s 268070 9150 272504 9210 6 addr[3]
port 4 nsew signal input
rlabel metal3 s 268162 9014 272504 9074 6 addr[4]
port 5 nsew signal input
rlabel metal3 s 272026 8878 272504 8938 6 k_one
port 6 nsew signal output
rlabel metal3 s 271830 8742 272504 8802 6 k_zero
port 7 nsew signal output
rlabel metal3 s 272304 8606 272504 8666 6 spine_iw[0]
port 8 nsew signal input
rlabel metal3 s 272026 7246 272504 7306 6 spine_iw[10]
port 9 nsew signal input
rlabel metal3 s 262550 7110 272504 7170 6 spine_iw[11]
port 10 nsew signal input
rlabel metal3 s 268070 6974 272504 7034 6 spine_iw[12]
port 11 nsew signal input
rlabel metal3 s 268162 6838 272504 6898 6 spine_iw[13]
port 12 nsew signal input
rlabel metal3 s 272118 6702 272504 6762 6 spine_iw[14]
port 13 nsew signal input
rlabel metal3 s 271934 6566 272504 6626 6 spine_iw[15]
port 14 nsew signal input
rlabel metal3 s 271830 6430 272504 6490 6 spine_iw[16]
port 15 nsew signal input
rlabel metal3 s 272026 6294 272504 6354 6 spine_iw[17]
port 16 nsew signal input
rlabel metal3 s 268990 6158 272504 6218 6 spine_iw[18]
port 17 nsew signal input
rlabel metal3 s 271842 6022 272504 6082 6 spine_iw[19]
port 18 nsew signal input
rlabel metal3 s 270646 8470 272504 8530 6 spine_iw[1]
port 19 nsew signal input
rlabel metal3 s 271750 5886 272504 5946 6 spine_iw[20]
port 20 nsew signal input
rlabel metal3 s 271462 5750 272504 5810 6 spine_iw[21]
port 21 nsew signal input
rlabel metal3 s 271278 5614 272504 5674 6 spine_iw[22]
port 22 nsew signal input
rlabel metal3 s 271842 5478 272504 5538 6 spine_iw[23]
port 23 nsew signal input
rlabel metal3 s 272026 5342 272504 5402 6 spine_iw[24]
port 24 nsew signal input
rlabel metal3 s 268990 5206 272504 5266 6 spine_iw[25]
port 25 nsew signal input
rlabel metal3 s 272026 5070 272504 5130 6 spine_iw[26]
port 26 nsew signal input
rlabel metal3 s 268162 4934 272504 4994 6 spine_iw[27]
port 27 nsew signal input
rlabel metal3 s 268898 4798 272504 4858 6 spine_iw[28]
port 28 nsew signal input
rlabel metal3 s 272210 4662 272504 4722 6 spine_iw[29]
port 29 nsew signal input
rlabel metal3 s 271290 8334 272504 8394 6 spine_iw[2]
port 30 nsew signal input
rlabel metal3 s 272304 4526 272504 4586 6 spine_iw[30]
port 31 nsew signal input
rlabel metal3 s 270554 8198 272504 8258 6 spine_iw[3]
port 32 nsew signal input
rlabel metal3 s 270370 8062 272504 8122 6 spine_iw[4]
port 33 nsew signal input
rlabel metal3 s 270186 7926 272504 7986 6 spine_iw[5]
port 34 nsew signal input
rlabel metal3 s 268070 7790 272504 7850 6 spine_iw[6]
port 35 nsew signal input
rlabel metal3 s 271842 7654 272504 7714 6 spine_iw[7]
port 36 nsew signal input
rlabel metal3 s 271842 7518 272504 7578 6 spine_iw[8]
port 37 nsew signal input
rlabel metal3 s 268070 7382 272504 7442 6 spine_iw[9]
port 38 nsew signal input
rlabel metal3 s 271968 4390 272504 4450 6 spine_ow[0]
port 39 nsew signal output
rlabel metal3 s 262274 3030 272504 3090 6 spine_ow[10]
port 40 nsew signal output
rlabel metal3 s 272026 2894 272504 2954 6 spine_ow[11]
port 41 nsew signal output
rlabel metal3 s 270830 2758 272504 2818 6 spine_ow[12]
port 42 nsew signal output
rlabel metal3 s 267242 2622 272504 2682 6 spine_ow[13]
port 43 nsew signal output
rlabel metal3 s 268530 2486 272504 2546 6 spine_ow[14]
port 44 nsew signal output
rlabel metal3 s 272026 2350 272504 2410 6 spine_ow[15]
port 45 nsew signal output
rlabel metal3 s 271830 2214 272504 2274 6 spine_ow[16]
port 46 nsew signal output
rlabel metal3 s 271842 2078 272504 2138 6 spine_ow[17]
port 47 nsew signal output
rlabel metal3 s 272210 1942 272504 2002 6 spine_ow[18]
port 48 nsew signal output
rlabel metal3 s 270174 1806 272504 1866 6 spine_ow[19]
port 49 nsew signal output
rlabel metal3 s 271830 4254 272504 4314 6 spine_ow[1]
port 50 nsew signal output
rlabel metal3 s 269990 1670 272504 1730 6 spine_ow[20]
port 51 nsew signal output
rlabel metal3 s 269082 1534 272504 1594 6 spine_ow[21]
port 52 nsew signal output
rlabel metal3 s 268898 1398 272504 1458 6 spine_ow[22]
port 53 nsew signal output
rlabel metal3 s 268886 1262 272504 1322 6 spine_ow[23]
port 54 nsew signal output
rlabel metal3 s 271842 1126 272504 1186 6 spine_ow[24]
port 55 nsew signal output
rlabel metal3 s 271830 990 272504 1050 6 spine_ow[25]
port 56 nsew signal output
rlabel metal3 s 244242 4118 272504 4178 6 spine_ow[2]
port 57 nsew signal output
rlabel metal3 s 271278 3982 272504 4042 6 spine_ow[3]
port 58 nsew signal output
rlabel metal3 s 271462 3846 272504 3906 6 spine_ow[4]
port 59 nsew signal output
rlabel metal3 s 271658 3710 272504 3770 6 spine_ow[5]
port 60 nsew signal output
rlabel metal3 s 267978 3574 272504 3634 6 spine_ow[6]
port 61 nsew signal output
rlabel metal3 s 272026 3438 272504 3498 6 spine_ow[7]
port 62 nsew signal output
rlabel metal3 s 271830 3302 272504 3362 6 spine_ow[8]
port 63 nsew signal output
rlabel metal3 s 271842 3166 272504 3226 6 spine_ow[9]
port 64 nsew signal output
rlabel metal4 s 32446 0 32506 1396 6 um_ena[0]
port 65 nsew signal output
rlabel metal4 s 203106 0 203166 370 6 um_ena[10]
port 66 nsew signal output
rlabel metal4 s 203106 10300 203166 10880 6 um_ena[11]
port 67 nsew signal output
rlabel metal4 s 237238 0 237298 1396 6 um_ena[12]
port 68 nsew signal output
rlabel metal4 s 237238 9212 237298 10880 6 um_ena[13]
port 69 nsew signal output
rlabel metal4 s 271370 0 271430 308 6 um_ena[14]
port 70 nsew signal output
rlabel metal4 s 271370 10238 271430 10880 6 um_ena[15]
port 71 nsew signal output
rlabel metal4 s 32446 9620 32506 10880 6 um_ena[1]
port 72 nsew signal output
rlabel metal4 s 66578 0 66638 444 6 um_ena[2]
port 73 nsew signal output
rlabel metal4 s 66578 10300 66638 10880 6 um_ena[3]
port 74 nsew signal output
rlabel metal4 s 100710 0 100770 852 6 um_ena[4]
port 75 nsew signal output
rlabel metal4 s 100710 9756 100770 10880 6 um_ena[5]
port 76 nsew signal output
rlabel metal4 s 134842 0 134902 370 6 um_ena[6]
port 77 nsew signal output
rlabel metal4 s 134842 10300 134902 10880 6 um_ena[7]
port 78 nsew signal output
rlabel metal4 s 168974 0 169034 580 6 um_ena[8]
port 79 nsew signal output
rlabel metal4 s 168974 9212 169034 10880 6 um_ena[9]
port 80 nsew signal output
rlabel metal4 s 31710 0 31770 444 6 um_iw[0]
port 81 nsew signal output
rlabel metal4 s 92614 8396 92674 10880 6 um_iw[100]
port 82 nsew signal output
rlabel metal4 s 91878 8668 91938 10880 6 um_iw[101]
port 83 nsew signal output
rlabel metal4 s 91142 8804 91202 10880 6 um_iw[102]
port 84 nsew signal output
rlabel metal4 s 90406 8668 90466 10880 6 um_iw[103]
port 85 nsew signal output
rlabel metal4 s 89670 10300 89730 10880 6 um_iw[104]
port 86 nsew signal output
rlabel metal4 s 88934 8124 88994 10880 6 um_iw[105]
port 87 nsew signal output
rlabel metal4 s 88198 9212 88258 10880 6 um_iw[106]
port 88 nsew signal output
rlabel metal4 s 87462 8668 87522 10880 6 um_iw[107]
port 89 nsew signal output
rlabel metal4 s 134106 0 134166 580 6 um_iw[108]
port 90 nsew signal output
rlabel metal4 s 133370 0 133430 580 6 um_iw[109]
port 91 nsew signal output
rlabel metal4 s 24350 0 24410 3300 6 um_iw[10]
port 92 nsew signal output
rlabel metal4 s 132634 0 132694 580 6 um_iw[110]
port 93 nsew signal output
rlabel metal4 s 131898 0 131958 580 6 um_iw[111]
port 94 nsew signal output
rlabel metal4 s 131162 0 131222 580 6 um_iw[112]
port 95 nsew signal output
rlabel metal4 s 130426 0 130486 308 6 um_iw[113]
port 96 nsew signal output
rlabel metal4 s 129690 0 129750 580 6 um_iw[114]
port 97 nsew signal output
rlabel metal4 s 128954 0 129014 580 6 um_iw[115]
port 98 nsew signal output
rlabel metal4 s 128218 0 128278 370 6 um_iw[116]
port 99 nsew signal output
rlabel metal4 s 127482 0 127542 580 6 um_iw[117]
port 100 nsew signal output
rlabel metal4 s 126746 0 126806 580 6 um_iw[118]
port 101 nsew signal output
rlabel metal4 s 126010 0 126070 580 6 um_iw[119]
port 102 nsew signal output
rlabel metal4 s 23614 0 23674 580 6 um_iw[11]
port 103 nsew signal output
rlabel metal4 s 125274 0 125334 580 6 um_iw[120]
port 104 nsew signal output
rlabel metal4 s 124538 0 124598 580 6 um_iw[121]
port 105 nsew signal output
rlabel metal4 s 123802 0 123862 580 6 um_iw[122]
port 106 nsew signal output
rlabel metal4 s 123066 0 123126 580 6 um_iw[123]
port 107 nsew signal output
rlabel metal4 s 122330 0 122390 580 6 um_iw[124]
port 108 nsew signal output
rlabel metal4 s 121594 0 121654 580 6 um_iw[125]
port 109 nsew signal output
rlabel metal4 s 134106 10300 134166 10880 6 um_iw[126]
port 110 nsew signal output
rlabel metal4 s 133370 10300 133430 10880 6 um_iw[127]
port 111 nsew signal output
rlabel metal4 s 132634 10300 132694 10880 6 um_iw[128]
port 112 nsew signal output
rlabel metal4 s 131898 10300 131958 10880 6 um_iw[129]
port 113 nsew signal output
rlabel metal4 s 22878 0 22938 2892 6 um_iw[12]
port 114 nsew signal output
rlabel metal4 s 131162 10300 131222 10880 6 um_iw[130]
port 115 nsew signal output
rlabel metal4 s 130426 10300 130486 10880 6 um_iw[131]
port 116 nsew signal output
rlabel metal4 s 129690 10300 129750 10880 6 um_iw[132]
port 117 nsew signal output
rlabel metal4 s 128954 10300 129014 10880 6 um_iw[133]
port 118 nsew signal output
rlabel metal4 s 128218 10436 128278 10880 6 um_iw[134]
port 119 nsew signal output
rlabel metal4 s 127482 10300 127542 10880 6 um_iw[135]
port 120 nsew signal output
rlabel metal4 s 126746 10300 126806 10880 6 um_iw[136]
port 121 nsew signal output
rlabel metal4 s 126010 10300 126070 10880 6 um_iw[137]
port 122 nsew signal output
rlabel metal4 s 125274 10436 125334 10880 6 um_iw[138]
port 123 nsew signal output
rlabel metal4 s 124538 10300 124598 10880 6 um_iw[139]
port 124 nsew signal output
rlabel metal4 s 22142 0 22202 2756 6 um_iw[13]
port 125 nsew signal output
rlabel metal4 s 123802 10300 123862 10880 6 um_iw[140]
port 126 nsew signal output
rlabel metal4 s 123066 10300 123126 10880 6 um_iw[141]
port 127 nsew signal output
rlabel metal4 s 122330 10300 122390 10880 6 um_iw[142]
port 128 nsew signal output
rlabel metal4 s 121594 10300 121654 10880 6 um_iw[143]
port 129 nsew signal output
rlabel metal4 s 168238 0 168298 1396 6 um_iw[144]
port 130 nsew signal output
rlabel metal4 s 167502 0 167562 580 6 um_iw[145]
port 131 nsew signal output
rlabel metal4 s 166766 0 166826 1124 6 um_iw[146]
port 132 nsew signal output
rlabel metal4 s 166030 0 166090 1124 6 um_iw[147]
port 133 nsew signal output
rlabel metal4 s 165294 0 165354 1124 6 um_iw[148]
port 134 nsew signal output
rlabel metal4 s 164558 0 164618 580 6 um_iw[149]
port 135 nsew signal output
rlabel metal4 s 21406 0 21466 1668 6 um_iw[14]
port 136 nsew signal output
rlabel metal4 s 163822 0 163882 1396 6 um_iw[150]
port 137 nsew signal output
rlabel metal4 s 163086 0 163146 1124 6 um_iw[151]
port 138 nsew signal output
rlabel metal4 s 162350 0 162410 580 6 um_iw[152]
port 139 nsew signal output
rlabel metal4 s 161614 0 161674 1124 6 um_iw[153]
port 140 nsew signal output
rlabel metal4 s 160878 0 160938 580 6 um_iw[154]
port 141 nsew signal output
rlabel metal4 s 160142 0 160202 1124 6 um_iw[155]
port 142 nsew signal output
rlabel metal4 s 159406 0 159466 2756 6 um_iw[156]
port 143 nsew signal output
rlabel metal4 s 158670 0 158730 580 6 um_iw[157]
port 144 nsew signal output
rlabel metal4 s 157934 0 157994 1396 6 um_iw[158]
port 145 nsew signal output
rlabel metal4 s 157198 0 157258 2756 6 um_iw[159]
port 146 nsew signal output
rlabel metal4 s 20670 0 20730 1396 6 um_iw[15]
port 147 nsew signal output
rlabel metal4 s 156462 0 156522 1396 6 um_iw[160]
port 148 nsew signal output
rlabel metal4 s 155726 0 155786 1396 6 um_iw[161]
port 149 nsew signal output
rlabel metal4 s 168238 8124 168298 10880 6 um_iw[162]
port 150 nsew signal output
rlabel metal4 s 167502 8396 167562 10880 6 um_iw[163]
port 151 nsew signal output
rlabel metal4 s 166766 8260 166826 10880 6 um_iw[164]
port 152 nsew signal output
rlabel metal4 s 166030 8396 166090 10880 6 um_iw[165]
port 153 nsew signal output
rlabel metal4 s 165294 8396 165354 10880 6 um_iw[166]
port 154 nsew signal output
rlabel metal4 s 164558 8396 164618 10880 6 um_iw[167]
port 155 nsew signal output
rlabel metal4 s 163822 9756 163882 10880 6 um_iw[168]
port 156 nsew signal output
rlabel metal4 s 163086 8396 163146 10880 6 um_iw[169]
port 157 nsew signal output
rlabel metal4 s 19934 0 19994 2756 6 um_iw[16]
port 158 nsew signal output
rlabel metal4 s 162350 8396 162410 10880 6 um_iw[170]
port 159 nsew signal output
rlabel metal4 s 161614 8532 161674 10880 6 um_iw[171]
port 160 nsew signal output
rlabel metal4 s 160878 8396 160938 10880 6 um_iw[172]
port 161 nsew signal output
rlabel metal4 s 160142 8396 160202 10880 6 um_iw[173]
port 162 nsew signal output
rlabel metal4 s 159406 9756 159466 10880 6 um_iw[174]
port 163 nsew signal output
rlabel metal4 s 158670 9484 158730 10880 6 um_iw[175]
port 164 nsew signal output
rlabel metal4 s 157934 9756 157994 10880 6 um_iw[176]
port 165 nsew signal output
rlabel metal4 s 157198 10300 157258 10880 6 um_iw[177]
port 166 nsew signal output
rlabel metal4 s 156462 9756 156522 10880 6 um_iw[178]
port 167 nsew signal output
rlabel metal4 s 155726 9756 155786 10880 6 um_iw[179]
port 168 nsew signal output
rlabel metal4 s 19198 0 19258 2892 6 um_iw[17]
port 169 nsew signal output
rlabel metal4 s 202370 0 202430 370 6 um_iw[180]
port 170 nsew signal output
rlabel metal4 s 201634 0 201694 370 6 um_iw[181]
port 171 nsew signal output
rlabel metal4 s 200898 0 200958 370 6 um_iw[182]
port 172 nsew signal output
rlabel metal4 s 200162 0 200222 370 6 um_iw[183]
port 173 nsew signal output
rlabel metal4 s 199426 0 199486 370 6 um_iw[184]
port 174 nsew signal output
rlabel metal4 s 198690 0 198750 370 6 um_iw[185]
port 175 nsew signal output
rlabel metal4 s 197954 0 198014 370 6 um_iw[186]
port 176 nsew signal output
rlabel metal4 s 197218 0 197278 370 6 um_iw[187]
port 177 nsew signal output
rlabel metal4 s 196482 0 196542 370 6 um_iw[188]
port 178 nsew signal output
rlabel metal4 s 195746 0 195806 370 6 um_iw[189]
port 179 nsew signal output
rlabel metal4 s 31710 10300 31770 10880 6 um_iw[18]
port 180 nsew signal output
rlabel metal4 s 195010 0 195070 370 6 um_iw[190]
port 181 nsew signal output
rlabel metal4 s 194274 0 194334 370 6 um_iw[191]
port 182 nsew signal output
rlabel metal4 s 193538 0 193598 370 6 um_iw[192]
port 183 nsew signal output
rlabel metal4 s 192802 0 192862 370 6 um_iw[193]
port 184 nsew signal output
rlabel metal4 s 192066 0 192126 370 6 um_iw[194]
port 185 nsew signal output
rlabel metal4 s 191330 0 191390 370 6 um_iw[195]
port 186 nsew signal output
rlabel metal4 s 190594 0 190654 370 6 um_iw[196]
port 187 nsew signal output
rlabel metal4 s 189858 0 189918 370 6 um_iw[197]
port 188 nsew signal output
rlabel metal4 s 202370 10436 202430 10880 6 um_iw[198]
port 189 nsew signal output
rlabel metal4 s 201634 10300 201694 10880 6 um_iw[199]
port 190 nsew signal output
rlabel metal4 s 30974 8668 31034 10880 6 um_iw[19]
port 191 nsew signal output
rlabel metal4 s 30974 0 31034 308 6 um_iw[1]
port 192 nsew signal output
rlabel metal4 s 200898 10436 200958 10880 6 um_iw[200]
port 193 nsew signal output
rlabel metal4 s 200162 10300 200222 10880 6 um_iw[201]
port 194 nsew signal output
rlabel metal4 s 199426 10300 199486 10880 6 um_iw[202]
port 195 nsew signal output
rlabel metal4 s 198690 10436 198750 10880 6 um_iw[203]
port 196 nsew signal output
rlabel metal4 s 197954 10300 198014 10880 6 um_iw[204]
port 197 nsew signal output
rlabel metal4 s 197218 10300 197278 10880 6 um_iw[205]
port 198 nsew signal output
rlabel metal4 s 196482 10300 196542 10880 6 um_iw[206]
port 199 nsew signal output
rlabel metal4 s 195746 10300 195806 10880 6 um_iw[207]
port 200 nsew signal output
rlabel metal4 s 195010 10300 195070 10880 6 um_iw[208]
port 201 nsew signal output
rlabel metal4 s 194274 10300 194334 10880 6 um_iw[209]
port 202 nsew signal output
rlabel metal4 s 30238 8668 30298 10880 6 um_iw[20]
port 203 nsew signal output
rlabel metal4 s 193538 10436 193598 10880 6 um_iw[210]
port 204 nsew signal output
rlabel metal4 s 192802 10300 192862 10880 6 um_iw[211]
port 205 nsew signal output
rlabel metal4 s 192066 10300 192126 10880 6 um_iw[212]
port 206 nsew signal output
rlabel metal4 s 191330 10300 191390 10880 6 um_iw[213]
port 207 nsew signal output
rlabel metal4 s 190594 10436 190654 10880 6 um_iw[214]
port 208 nsew signal output
rlabel metal4 s 189858 10300 189918 10880 6 um_iw[215]
port 209 nsew signal output
rlabel metal4 s 236502 0 236562 1124 6 um_iw[216]
port 210 nsew signal output
rlabel metal4 s 235766 0 235826 2756 6 um_iw[217]
port 211 nsew signal output
rlabel metal4 s 235030 0 235090 444 6 um_iw[218]
port 212 nsew signal output
rlabel metal4 s 234294 0 234354 308 6 um_iw[219]
port 213 nsew signal output
rlabel metal4 s 29502 8668 29562 10880 6 um_iw[21]
port 214 nsew signal output
rlabel metal4 s 233558 0 233618 308 6 um_iw[220]
port 215 nsew signal output
rlabel metal4 s 232822 0 232882 1124 6 um_iw[221]
port 216 nsew signal output
rlabel metal4 s 232086 0 232146 1124 6 um_iw[222]
port 217 nsew signal output
rlabel metal4 s 231350 0 231410 1124 6 um_iw[223]
port 218 nsew signal output
rlabel metal4 s 230614 0 230674 308 6 um_iw[224]
port 219 nsew signal output
rlabel metal4 s 229878 0 229938 308 6 um_iw[225]
port 220 nsew signal output
rlabel metal4 s 229142 0 229202 308 6 um_iw[226]
port 221 nsew signal output
rlabel metal4 s 228406 0 228466 1124 6 um_iw[227]
port 222 nsew signal output
rlabel metal4 s 227670 0 227730 1260 6 um_iw[228]
port 223 nsew signal output
rlabel metal4 s 226934 0 226994 1260 6 um_iw[229]
port 224 nsew signal output
rlabel metal4 s 28766 9484 28826 10880 6 um_iw[22]
port 225 nsew signal output
rlabel metal4 s 226198 0 226258 2756 6 um_iw[230]
port 226 nsew signal output
rlabel metal4 s 225462 0 225522 1396 6 um_iw[231]
port 227 nsew signal output
rlabel metal4 s 224726 0 224786 2756 6 um_iw[232]
port 228 nsew signal output
rlabel metal4 s 223990 0 224050 1396 6 um_iw[233]
port 229 nsew signal output
rlabel metal4 s 236502 8668 236562 10880 6 um_iw[234]
port 230 nsew signal output
rlabel metal4 s 235766 9212 235826 10880 6 um_iw[235]
port 231 nsew signal output
rlabel metal4 s 235030 9756 235090 10880 6 um_iw[236]
port 232 nsew signal output
rlabel metal4 s 234294 9756 234354 10880 6 um_iw[237]
port 233 nsew signal output
rlabel metal4 s 233558 9756 233618 10880 6 um_iw[238]
port 234 nsew signal output
rlabel metal4 s 232822 8668 232882 10880 6 um_iw[239]
port 235 nsew signal output
rlabel metal4 s 28030 8396 28090 10880 6 um_iw[23]
port 236 nsew signal output
rlabel metal4 s 232086 8668 232146 10880 6 um_iw[240]
port 237 nsew signal output
rlabel metal4 s 231350 9756 231410 10880 6 um_iw[241]
port 238 nsew signal output
rlabel metal4 s 230614 8396 230674 10880 6 um_iw[242]
port 239 nsew signal output
rlabel metal4 s 229878 9756 229938 10880 6 um_iw[243]
port 240 nsew signal output
rlabel metal4 s 229142 8668 229202 10880 6 um_iw[244]
port 241 nsew signal output
rlabel metal4 s 228406 9484 228466 10880 6 um_iw[245]
port 242 nsew signal output
rlabel metal4 s 227670 8668 227730 10880 6 um_iw[246]
port 243 nsew signal output
rlabel metal4 s 226934 8668 226994 10880 6 um_iw[247]
port 244 nsew signal output
rlabel metal4 s 226198 8668 226258 10880 6 um_iw[248]
port 245 nsew signal output
rlabel metal4 s 225462 9756 225522 10880 6 um_iw[249]
port 246 nsew signal output
rlabel metal4 s 27294 7852 27354 10880 6 um_iw[24]
port 247 nsew signal output
rlabel metal4 s 224726 8396 224786 10880 6 um_iw[250]
port 248 nsew signal output
rlabel metal4 s 223990 9212 224050 10880 6 um_iw[251]
port 249 nsew signal output
rlabel metal4 s 270634 0 270694 370 6 um_iw[252]
port 250 nsew signal output
rlabel metal4 s 269898 0 269958 580 6 um_iw[253]
port 251 nsew signal output
rlabel metal4 s 269162 0 269222 444 6 um_iw[254]
port 252 nsew signal output
rlabel metal4 s 268426 0 268486 580 6 um_iw[255]
port 253 nsew signal output
rlabel metal4 s 267690 0 267750 580 6 um_iw[256]
port 254 nsew signal output
rlabel metal4 s 266954 0 267014 580 6 um_iw[257]
port 255 nsew signal output
rlabel metal4 s 266218 0 266278 580 6 um_iw[258]
port 256 nsew signal output
rlabel metal4 s 265482 0 265542 580 6 um_iw[259]
port 257 nsew signal output
rlabel metal4 s 26558 8396 26618 10880 6 um_iw[25]
port 258 nsew signal output
rlabel metal4 s 264746 0 264806 370 6 um_iw[260]
port 259 nsew signal output
rlabel metal4 s 264010 0 264070 580 6 um_iw[261]
port 260 nsew signal output
rlabel metal4 s 263274 0 263334 580 6 um_iw[262]
port 261 nsew signal output
rlabel metal4 s 262538 0 262598 580 6 um_iw[263]
port 262 nsew signal output
rlabel metal4 s 261802 0 261862 444 6 um_iw[264]
port 263 nsew signal output
rlabel metal4 s 261066 0 261126 580 6 um_iw[265]
port 264 nsew signal output
rlabel metal4 s 260330 0 260390 580 6 um_iw[266]
port 265 nsew signal output
rlabel metal4 s 259594 0 259654 580 6 um_iw[267]
port 266 nsew signal output
rlabel metal4 s 258858 0 258918 580 6 um_iw[268]
port 267 nsew signal output
rlabel metal4 s 258122 0 258182 642 6 um_iw[269]
port 268 nsew signal output
rlabel metal4 s 25822 9620 25882 10880 6 um_iw[26]
port 269 nsew signal output
rlabel metal4 s 270634 10238 270694 10880 6 um_iw[270]
port 270 nsew signal output
rlabel metal4 s 269898 10238 269958 10880 6 um_iw[271]
port 271 nsew signal output
rlabel metal4 s 269162 10238 269222 10880 6 um_iw[272]
port 272 nsew signal output
rlabel metal4 s 268426 10238 268486 10880 6 um_iw[273]
port 273 nsew signal output
rlabel metal4 s 267690 10238 267750 10880 6 um_iw[274]
port 274 nsew signal output
rlabel metal4 s 266954 10238 267014 10880 6 um_iw[275]
port 275 nsew signal output
rlabel metal4 s 266218 10510 266278 10880 6 um_iw[276]
port 276 nsew signal output
rlabel metal4 s 265482 10300 265542 10880 6 um_iw[277]
port 277 nsew signal output
rlabel metal4 s 264746 10436 264806 10880 6 um_iw[278]
port 278 nsew signal output
rlabel metal4 s 264010 10300 264070 10880 6 um_iw[279]
port 279 nsew signal output
rlabel metal4 s 25086 6900 25146 10880 6 um_iw[27]
port 280 nsew signal output
rlabel metal4 s 263274 10300 263334 10880 6 um_iw[280]
port 281 nsew signal output
rlabel metal4 s 262538 10300 262598 10880 6 um_iw[281]
port 282 nsew signal output
rlabel metal4 s 261802 10300 261862 10880 6 um_iw[282]
port 283 nsew signal output
rlabel metal4 s 261066 10436 261126 10880 6 um_iw[283]
port 284 nsew signal output
rlabel metal4 s 260330 10300 260390 10880 6 um_iw[284]
port 285 nsew signal output
rlabel metal4 s 259594 10300 259654 10880 6 um_iw[285]
port 286 nsew signal output
rlabel metal4 s 258858 10300 258918 10880 6 um_iw[286]
port 287 nsew signal output
rlabel metal4 s 258122 10300 258182 10880 6 um_iw[287]
port 288 nsew signal output
rlabel metal4 s 24350 8668 24410 10880 6 um_iw[28]
port 289 nsew signal output
rlabel metal4 s 23614 6900 23674 10880 6 um_iw[29]
port 290 nsew signal output
rlabel metal4 s 30238 0 30298 580 6 um_iw[2]
port 291 nsew signal output
rlabel metal4 s 22878 6900 22938 10880 6 um_iw[30]
port 292 nsew signal output
rlabel metal4 s 22142 10164 22202 10880 6 um_iw[31]
port 293 nsew signal output
rlabel metal4 s 21406 9892 21466 10880 6 um_iw[32]
port 294 nsew signal output
rlabel metal4 s 20670 10572 20730 10880 6 um_iw[33]
port 295 nsew signal output
rlabel metal4 s 19934 6900 19994 10880 6 um_iw[34]
port 296 nsew signal output
rlabel metal4 s 19198 6900 19258 10880 6 um_iw[35]
port 297 nsew signal output
rlabel metal4 s 65842 0 65902 444 6 um_iw[36]
port 298 nsew signal output
rlabel metal4 s 65106 0 65166 580 6 um_iw[37]
port 299 nsew signal output
rlabel metal4 s 64370 0 64430 580 6 um_iw[38]
port 300 nsew signal output
rlabel metal4 s 63634 0 63694 580 6 um_iw[39]
port 301 nsew signal output
rlabel metal4 s 29502 0 29562 444 6 um_iw[3]
port 302 nsew signal output
rlabel metal4 s 62898 0 62958 580 6 um_iw[40]
port 303 nsew signal output
rlabel metal4 s 62162 0 62222 580 6 um_iw[41]
port 304 nsew signal output
rlabel metal4 s 61426 0 61486 580 6 um_iw[42]
port 305 nsew signal output
rlabel metal4 s 60690 0 60750 580 6 um_iw[43]
port 306 nsew signal output
rlabel metal4 s 59954 0 60014 370 6 um_iw[44]
port 307 nsew signal output
rlabel metal4 s 59218 0 59278 370 6 um_iw[45]
port 308 nsew signal output
rlabel metal4 s 58482 0 58542 580 6 um_iw[46]
port 309 nsew signal output
rlabel metal4 s 57746 0 57806 580 6 um_iw[47]
port 310 nsew signal output
rlabel metal4 s 57010 0 57070 580 6 um_iw[48]
port 311 nsew signal output
rlabel metal4 s 56274 0 56334 580 6 um_iw[49]
port 312 nsew signal output
rlabel metal4 s 28766 0 28826 580 6 um_iw[4]
port 313 nsew signal output
rlabel metal4 s 55538 0 55598 580 6 um_iw[50]
port 314 nsew signal output
rlabel metal4 s 54802 0 54862 580 6 um_iw[51]
port 315 nsew signal output
rlabel metal4 s 54066 0 54126 370 6 um_iw[52]
port 316 nsew signal output
rlabel metal4 s 53330 0 53390 580 6 um_iw[53]
port 317 nsew signal output
rlabel metal4 s 65842 10300 65902 10880 6 um_iw[54]
port 318 nsew signal output
rlabel metal4 s 65106 10300 65166 10880 6 um_iw[55]
port 319 nsew signal output
rlabel metal4 s 64370 10300 64430 10880 6 um_iw[56]
port 320 nsew signal output
rlabel metal4 s 63634 10300 63694 10880 6 um_iw[57]
port 321 nsew signal output
rlabel metal4 s 62898 10300 62958 10880 6 um_iw[58]
port 322 nsew signal output
rlabel metal4 s 62162 10300 62222 10880 6 um_iw[59]
port 323 nsew signal output
rlabel metal4 s 28030 0 28090 444 6 um_iw[5]
port 324 nsew signal output
rlabel metal4 s 61426 10300 61486 10880 6 um_iw[60]
port 325 nsew signal output
rlabel metal4 s 60690 10300 60750 10880 6 um_iw[61]
port 326 nsew signal output
rlabel metal4 s 59954 10300 60014 10880 6 um_iw[62]
port 327 nsew signal output
rlabel metal4 s 59218 10300 59278 10880 6 um_iw[63]
port 328 nsew signal output
rlabel metal4 s 58482 10300 58542 10880 6 um_iw[64]
port 329 nsew signal output
rlabel metal4 s 57746 10300 57806 10880 6 um_iw[65]
port 330 nsew signal output
rlabel metal4 s 57010 10300 57070 10880 6 um_iw[66]
port 331 nsew signal output
rlabel metal4 s 56274 10300 56334 10880 6 um_iw[67]
port 332 nsew signal output
rlabel metal4 s 55538 10300 55598 10880 6 um_iw[68]
port 333 nsew signal output
rlabel metal4 s 54802 10300 54862 10880 6 um_iw[69]
port 334 nsew signal output
rlabel metal4 s 27294 0 27354 1260 6 um_iw[6]
port 335 nsew signal output
rlabel metal4 s 54066 10436 54126 10880 6 um_iw[70]
port 336 nsew signal output
rlabel metal4 s 53330 10300 53390 10880 6 um_iw[71]
port 337 nsew signal output
rlabel metal4 s 99974 0 100034 444 6 um_iw[72]
port 338 nsew signal output
rlabel metal4 s 99238 0 99298 1532 6 um_iw[73]
port 339 nsew signal output
rlabel metal4 s 98502 0 98562 716 6 um_iw[74]
port 340 nsew signal output
rlabel metal4 s 97766 0 97826 716 6 um_iw[75]
port 341 nsew signal output
rlabel metal4 s 97030 0 97090 444 6 um_iw[76]
port 342 nsew signal output
rlabel metal4 s 96294 0 96354 1124 6 um_iw[77]
port 343 nsew signal output
rlabel metal4 s 95558 0 95618 1124 6 um_iw[78]
port 344 nsew signal output
rlabel metal4 s 94822 0 94882 1124 6 um_iw[79]
port 345 nsew signal output
rlabel metal4 s 26558 0 26618 1260 6 um_iw[7]
port 346 nsew signal output
rlabel metal4 s 94086 0 94146 1124 6 um_iw[80]
port 347 nsew signal output
rlabel metal4 s 93350 0 93410 716 6 um_iw[81]
port 348 nsew signal output
rlabel metal4 s 92614 0 92674 308 6 um_iw[82]
port 349 nsew signal output
rlabel metal4 s 91878 0 91938 716 6 um_iw[83]
port 350 nsew signal output
rlabel metal4 s 91142 0 91202 308 6 um_iw[84]
port 351 nsew signal output
rlabel metal4 s 90406 0 90466 716 6 um_iw[85]
port 352 nsew signal output
rlabel metal4 s 89670 0 89730 308 6 um_iw[86]
port 353 nsew signal output
rlabel metal4 s 88934 0 88994 1260 6 um_iw[87]
port 354 nsew signal output
rlabel metal4 s 88198 0 88258 1124 6 um_iw[88]
port 355 nsew signal output
rlabel metal4 s 87462 0 87522 1260 6 um_iw[89]
port 356 nsew signal output
rlabel metal4 s 25822 0 25882 1260 6 um_iw[8]
port 357 nsew signal output
rlabel metal4 s 99974 8668 100034 10880 6 um_iw[90]
port 358 nsew signal output
rlabel metal4 s 99238 8260 99298 10880 6 um_iw[91]
port 359 nsew signal output
rlabel metal4 s 98502 8668 98562 10880 6 um_iw[92]
port 360 nsew signal output
rlabel metal4 s 97766 9756 97826 10880 6 um_iw[93]
port 361 nsew signal output
rlabel metal4 s 97030 8668 97090 10880 6 um_iw[94]
port 362 nsew signal output
rlabel metal4 s 96294 9756 96354 10880 6 um_iw[95]
port 363 nsew signal output
rlabel metal4 s 95558 9756 95618 10880 6 um_iw[96]
port 364 nsew signal output
rlabel metal4 s 94822 8668 94882 10880 6 um_iw[97]
port 365 nsew signal output
rlabel metal4 s 94086 8668 94146 10880 6 um_iw[98]
port 366 nsew signal output
rlabel metal4 s 93350 9756 93410 10880 6 um_iw[99]
port 367 nsew signal output
rlabel metal4 s 25086 0 25146 2756 6 um_iw[9]
port 368 nsew signal output
rlabel metal4 s 798 0 858 1396 6 um_k_zero[0]
port 369 nsew signal output
rlabel metal4 s 171458 0 171518 370 6 um_k_zero[10]
port 370 nsew signal output
rlabel metal4 s 171458 10300 171518 10880 6 um_k_zero[11]
port 371 nsew signal output
rlabel metal4 s 205590 0 205650 370 6 um_k_zero[12]
port 372 nsew signal output
rlabel metal4 s 205590 9620 205650 10880 6 um_k_zero[13]
port 373 nsew signal output
rlabel metal4 s 239722 0 239782 308 6 um_k_zero[14]
port 374 nsew signal output
rlabel metal4 s 239722 10300 239782 10880 6 um_k_zero[15]
port 375 nsew signal output
rlabel metal4 s 798 9212 858 10880 6 um_k_zero[1]
port 376 nsew signal output
rlabel metal4 s 34930 0 34990 308 6 um_k_zero[2]
port 377 nsew signal output
rlabel metal4 s 34930 10300 34990 10880 6 um_k_zero[3]
port 378 nsew signal output
rlabel metal4 s 69062 0 69122 716 6 um_k_zero[4]
port 379 nsew signal output
rlabel metal4 s 69062 9620 69122 10880 6 um_k_zero[5]
port 380 nsew signal output
rlabel metal4 s 103194 0 103254 444 6 um_k_zero[6]
port 381 nsew signal output
rlabel metal4 s 103194 10300 103254 10880 6 um_k_zero[7]
port 382 nsew signal output
rlabel metal4 s 137326 0 137386 1396 6 um_k_zero[8]
port 383 nsew signal output
rlabel metal4 s 137326 9620 137386 10880 6 um_k_zero[9]
port 384 nsew signal output
rlabel metal4 s 18462 0 18522 580 6 um_ow[0]
port 385 nsew signal input
rlabel metal4 s 83782 0 83842 1532 6 um_ow[100]
port 386 nsew signal input
rlabel metal4 s 83046 0 83106 1532 6 um_ow[101]
port 387 nsew signal input
rlabel metal4 s 82310 0 82370 1260 6 um_ow[102]
port 388 nsew signal input
rlabel metal4 s 81574 0 81634 1532 6 um_ow[103]
port 389 nsew signal input
rlabel metal4 s 80838 0 80898 716 6 um_ow[104]
port 390 nsew signal input
rlabel metal4 s 80102 0 80162 1532 6 um_ow[105]
port 391 nsew signal input
rlabel metal4 s 79366 0 79426 1260 6 um_ow[106]
port 392 nsew signal input
rlabel metal4 s 78630 0 78690 716 6 um_ow[107]
port 393 nsew signal input
rlabel metal4 s 77894 0 77954 1260 6 um_ow[108]
port 394 nsew signal input
rlabel metal4 s 77158 0 77218 988 6 um_ow[109]
port 395 nsew signal input
rlabel metal4 s 11102 0 11162 580 6 um_ow[10]
port 396 nsew signal input
rlabel metal4 s 76422 0 76482 1260 6 um_ow[110]
port 397 nsew signal input
rlabel metal4 s 75686 0 75746 988 6 um_ow[111]
port 398 nsew signal input
rlabel metal4 s 74950 0 75010 580 6 um_ow[112]
port 399 nsew signal input
rlabel metal4 s 74214 0 74274 988 6 um_ow[113]
port 400 nsew signal input
rlabel metal4 s 73478 0 73538 1260 6 um_ow[114]
port 401 nsew signal input
rlabel metal4 s 72742 0 72802 580 6 um_ow[115]
port 402 nsew signal input
rlabel metal4 s 72006 0 72066 988 6 um_ow[116]
port 403 nsew signal input
rlabel metal4 s 71270 0 71330 1260 6 um_ow[117]
port 404 nsew signal input
rlabel metal4 s 70534 0 70594 988 6 um_ow[118]
port 405 nsew signal input
rlabel metal4 s 69798 0 69858 716 6 um_ow[119]
port 406 nsew signal input
rlabel metal4 s 10366 0 10426 580 6 um_ow[11]
port 407 nsew signal input
rlabel metal4 s 86726 10572 86786 10880 6 um_ow[120]
port 408 nsew signal input
rlabel metal4 s 85990 9892 86050 10880 6 um_ow[121]
port 409 nsew signal input
rlabel metal4 s 85254 9892 85314 10880 6 um_ow[122]
port 410 nsew signal input
rlabel metal4 s 84518 10572 84578 10880 6 um_ow[123]
port 411 nsew signal input
rlabel metal4 s 83782 10436 83842 10880 6 um_ow[124]
port 412 nsew signal input
rlabel metal4 s 83046 9620 83106 10880 6 um_ow[125]
port 413 nsew signal input
rlabel metal4 s 82310 10436 82370 10880 6 um_ow[126]
port 414 nsew signal input
rlabel metal4 s 81574 9756 81634 10880 6 um_ow[127]
port 415 nsew signal input
rlabel metal4 s 80838 9620 80898 10880 6 um_ow[128]
port 416 nsew signal input
rlabel metal4 s 80102 9076 80162 10880 6 um_ow[129]
port 417 nsew signal input
rlabel metal4 s 9630 0 9690 580 6 um_ow[12]
port 418 nsew signal input
rlabel metal4 s 79366 9756 79426 10880 6 um_ow[130]
port 419 nsew signal input
rlabel metal4 s 78630 9076 78690 10880 6 um_ow[131]
port 420 nsew signal input
rlabel metal4 s 77894 9620 77954 10880 6 um_ow[132]
port 421 nsew signal input
rlabel metal4 s 77158 10436 77218 10880 6 um_ow[133]
port 422 nsew signal input
rlabel metal4 s 76422 9756 76482 10880 6 um_ow[134]
port 423 nsew signal input
rlabel metal4 s 75686 9620 75746 10880 6 um_ow[135]
port 424 nsew signal input
rlabel metal4 s 74950 9076 75010 10880 6 um_ow[136]
port 425 nsew signal input
rlabel metal4 s 74214 10572 74274 10880 6 um_ow[137]
port 426 nsew signal input
rlabel metal4 s 73478 9076 73538 10880 6 um_ow[138]
port 427 nsew signal input
rlabel metal4 s 72742 9620 72802 10880 6 um_ow[139]
port 428 nsew signal input
rlabel metal4 s 8894 0 8954 716 6 um_ow[13]
port 429 nsew signal input
rlabel metal4 s 72006 10436 72066 10880 6 um_ow[140]
port 430 nsew signal input
rlabel metal4 s 71270 10572 71330 10880 6 um_ow[141]
port 431 nsew signal input
rlabel metal4 s 70534 9620 70594 10880 6 um_ow[142]
port 432 nsew signal input
rlabel metal4 s 69798 9076 69858 10880 6 um_ow[143]
port 433 nsew signal input
rlabel metal4 s 120858 0 120918 580 6 um_ow[144]
port 434 nsew signal input
rlabel metal4 s 120122 0 120182 580 6 um_ow[145]
port 435 nsew signal input
rlabel metal4 s 119386 0 119446 580 6 um_ow[146]
port 436 nsew signal input
rlabel metal4 s 118650 0 118710 580 6 um_ow[147]
port 437 nsew signal input
rlabel metal4 s 117914 0 117974 580 6 um_ow[148]
port 438 nsew signal input
rlabel metal4 s 117178 0 117238 370 6 um_ow[149]
port 439 nsew signal input
rlabel metal4 s 8158 0 8218 580 6 um_ow[14]
port 440 nsew signal input
rlabel metal4 s 116442 0 116502 580 6 um_ow[150]
port 441 nsew signal input
rlabel metal4 s 115706 0 115766 580 6 um_ow[151]
port 442 nsew signal input
rlabel metal4 s 114970 0 115030 580 6 um_ow[152]
port 443 nsew signal input
rlabel metal4 s 114234 0 114294 580 6 um_ow[153]
port 444 nsew signal input
rlabel metal4 s 113498 0 113558 308 6 um_ow[154]
port 445 nsew signal input
rlabel metal4 s 112762 0 112822 444 6 um_ow[155]
port 446 nsew signal input
rlabel metal4 s 112026 0 112086 444 6 um_ow[156]
port 447 nsew signal input
rlabel metal4 s 111290 0 111350 444 6 um_ow[157]
port 448 nsew signal input
rlabel metal4 s 110554 0 110614 444 6 um_ow[158]
port 449 nsew signal input
rlabel metal4 s 109818 0 109878 444 6 um_ow[159]
port 450 nsew signal input
rlabel metal4 s 7422 0 7482 716 6 um_ow[15]
port 451 nsew signal input
rlabel metal4 s 109082 0 109142 444 6 um_ow[160]
port 452 nsew signal input
rlabel metal4 s 108346 0 108406 444 6 um_ow[161]
port 453 nsew signal input
rlabel metal4 s 107610 0 107670 444 6 um_ow[162]
port 454 nsew signal input
rlabel metal4 s 106874 0 106934 444 6 um_ow[163]
port 455 nsew signal input
rlabel metal4 s 106138 0 106198 444 6 um_ow[164]
port 456 nsew signal input
rlabel metal4 s 105402 0 105462 444 6 um_ow[165]
port 457 nsew signal input
rlabel metal4 s 104666 0 104726 444 6 um_ow[166]
port 458 nsew signal input
rlabel metal4 s 103930 0 103990 444 6 um_ow[167]
port 459 nsew signal input
rlabel metal4 s 120858 10300 120918 10880 6 um_ow[168]
port 460 nsew signal input
rlabel metal4 s 120122 10300 120182 10880 6 um_ow[169]
port 461 nsew signal input
rlabel metal4 s 6686 0 6746 988 6 um_ow[16]
port 462 nsew signal input
rlabel metal4 s 119386 10300 119446 10880 6 um_ow[170]
port 463 nsew signal input
rlabel metal4 s 118650 10300 118710 10880 6 um_ow[171]
port 464 nsew signal input
rlabel metal4 s 117914 10300 117974 10880 6 um_ow[172]
port 465 nsew signal input
rlabel metal4 s 117178 10300 117238 10880 6 um_ow[173]
port 466 nsew signal input
rlabel metal4 s 116442 10300 116502 10880 6 um_ow[174]
port 467 nsew signal input
rlabel metal4 s 115706 10300 115766 10880 6 um_ow[175]
port 468 nsew signal input
rlabel metal4 s 114970 10300 115030 10880 6 um_ow[176]
port 469 nsew signal input
rlabel metal4 s 114234 10300 114294 10880 6 um_ow[177]
port 470 nsew signal input
rlabel metal4 s 113498 10300 113558 10880 6 um_ow[178]
port 471 nsew signal input
rlabel metal4 s 112762 10300 112822 10880 6 um_ow[179]
port 472 nsew signal input
rlabel metal4 s 5950 0 6010 716 6 um_ow[17]
port 473 nsew signal input
rlabel metal4 s 112026 10300 112086 10880 6 um_ow[180]
port 474 nsew signal input
rlabel metal4 s 111290 10300 111350 10880 6 um_ow[181]
port 475 nsew signal input
rlabel metal4 s 110554 10300 110614 10880 6 um_ow[182]
port 476 nsew signal input
rlabel metal4 s 109818 10300 109878 10880 6 um_ow[183]
port 477 nsew signal input
rlabel metal4 s 109082 10300 109142 10880 6 um_ow[184]
port 478 nsew signal input
rlabel metal4 s 108346 10300 108406 10880 6 um_ow[185]
port 479 nsew signal input
rlabel metal4 s 107610 10300 107670 10880 6 um_ow[186]
port 480 nsew signal input
rlabel metal4 s 106874 10300 106934 10880 6 um_ow[187]
port 481 nsew signal input
rlabel metal4 s 106138 10300 106198 10880 6 um_ow[188]
port 482 nsew signal input
rlabel metal4 s 105402 10300 105462 10880 6 um_ow[189]
port 483 nsew signal input
rlabel metal4 s 5214 0 5274 716 6 um_ow[18]
port 484 nsew signal input
rlabel metal4 s 104666 10300 104726 10880 6 um_ow[190]
port 485 nsew signal input
rlabel metal4 s 103930 10300 103990 10880 6 um_ow[191]
port 486 nsew signal input
rlabel metal4 s 154990 0 155050 1260 6 um_ow[192]
port 487 nsew signal input
rlabel metal4 s 154254 0 154314 716 6 um_ow[193]
port 488 nsew signal input
rlabel metal4 s 153518 0 153578 580 6 um_ow[194]
port 489 nsew signal input
rlabel metal4 s 152782 0 152842 716 6 um_ow[195]
port 490 nsew signal input
rlabel metal4 s 152046 0 152106 716 6 um_ow[196]
port 491 nsew signal input
rlabel metal4 s 151310 0 151370 716 6 um_ow[197]
port 492 nsew signal input
rlabel metal4 s 150574 0 150634 716 6 um_ow[198]
port 493 nsew signal input
rlabel metal4 s 149838 0 149898 988 6 um_ow[199]
port 494 nsew signal input
rlabel metal4 s 4478 0 4538 988 6 um_ow[19]
port 495 nsew signal input
rlabel metal4 s 17726 0 17786 580 6 um_ow[1]
port 496 nsew signal input
rlabel metal4 s 149102 0 149162 716 6 um_ow[200]
port 497 nsew signal input
rlabel metal4 s 148366 0 148426 716 6 um_ow[201]
port 498 nsew signal input
rlabel metal4 s 147630 0 147690 580 6 um_ow[202]
port 499 nsew signal input
rlabel metal4 s 146894 0 146954 716 6 um_ow[203]
port 500 nsew signal input
rlabel metal4 s 146158 0 146218 716 6 um_ow[204]
port 501 nsew signal input
rlabel metal4 s 145422 0 145482 716 6 um_ow[205]
port 502 nsew signal input
rlabel metal4 s 144686 0 144746 1396 6 um_ow[206]
port 503 nsew signal input
rlabel metal4 s 143950 0 144010 716 6 um_ow[207]
port 504 nsew signal input
rlabel metal4 s 143214 0 143274 716 6 um_ow[208]
port 505 nsew signal input
rlabel metal4 s 142478 0 142538 988 6 um_ow[209]
port 506 nsew signal input
rlabel metal4 s 3742 0 3802 580 6 um_ow[20]
port 507 nsew signal input
rlabel metal4 s 141742 0 141802 580 6 um_ow[210]
port 508 nsew signal input
rlabel metal4 s 141006 0 141066 716 6 um_ow[211]
port 509 nsew signal input
rlabel metal4 s 140270 0 140330 1260 6 um_ow[212]
port 510 nsew signal input
rlabel metal4 s 139534 0 139594 444 6 um_ow[213]
port 511 nsew signal input
rlabel metal4 s 138798 0 138858 716 6 um_ow[214]
port 512 nsew signal input
rlabel metal4 s 138062 0 138122 580 6 um_ow[215]
port 513 nsew signal input
rlabel metal4 s 154990 9892 155050 10880 6 um_ow[216]
port 514 nsew signal input
rlabel metal4 s 154254 10164 154314 10880 6 um_ow[217]
port 515 nsew signal input
rlabel metal4 s 153518 10300 153578 10880 6 um_ow[218]
port 516 nsew signal input
rlabel metal4 s 152782 10164 152842 10880 6 um_ow[219]
port 517 nsew signal input
rlabel metal4 s 3006 0 3066 716 6 um_ow[21]
port 518 nsew signal input
rlabel metal4 s 152046 10164 152106 10880 6 um_ow[220]
port 519 nsew signal input
rlabel metal4 s 151310 10164 151370 10880 6 um_ow[221]
port 520 nsew signal input
rlabel metal4 s 150574 10164 150634 10880 6 um_ow[222]
port 521 nsew signal input
rlabel metal4 s 149838 9892 149898 10880 6 um_ow[223]
port 522 nsew signal input
rlabel metal4 s 149102 10164 149162 10880 6 um_ow[224]
port 523 nsew signal input
rlabel metal4 s 148366 10164 148426 10880 6 um_ow[225]
port 524 nsew signal input
rlabel metal4 s 147630 10436 147690 10880 6 um_ow[226]
port 525 nsew signal input
rlabel metal4 s 146894 10164 146954 10880 6 um_ow[227]
port 526 nsew signal input
rlabel metal4 s 146158 10164 146218 10880 6 um_ow[228]
port 527 nsew signal input
rlabel metal4 s 145422 10164 145482 10880 6 um_ow[229]
port 528 nsew signal input
rlabel metal4 s 2270 0 2330 988 6 um_ow[22]
port 529 nsew signal input
rlabel metal4 s 144686 9892 144746 10880 6 um_ow[230]
port 530 nsew signal input
rlabel metal4 s 143950 10164 144010 10880 6 um_ow[231]
port 531 nsew signal input
rlabel metal4 s 143214 10164 143274 10880 6 um_ow[232]
port 532 nsew signal input
rlabel metal4 s 142478 10300 142538 10880 6 um_ow[233]
port 533 nsew signal input
rlabel metal4 s 141742 10164 141802 10880 6 um_ow[234]
port 534 nsew signal input
rlabel metal4 s 141006 10164 141066 10880 6 um_ow[235]
port 535 nsew signal input
rlabel metal4 s 140270 10164 140330 10880 6 um_ow[236]
port 536 nsew signal input
rlabel metal4 s 139534 9892 139594 10880 6 um_ow[237]
port 537 nsew signal input
rlabel metal4 s 138798 10164 138858 10880 6 um_ow[238]
port 538 nsew signal input
rlabel metal4 s 138062 10300 138122 10880 6 um_ow[239]
port 539 nsew signal input
rlabel metal4 s 1534 0 1594 1260 6 um_ow[23]
port 540 nsew signal input
rlabel metal4 s 189122 0 189182 370 6 um_ow[240]
port 541 nsew signal input
rlabel metal4 s 188386 0 188446 370 6 um_ow[241]
port 542 nsew signal input
rlabel metal4 s 187650 0 187710 370 6 um_ow[242]
port 543 nsew signal input
rlabel metal4 s 186914 0 186974 370 6 um_ow[243]
port 544 nsew signal input
rlabel metal4 s 186178 0 186238 370 6 um_ow[244]
port 545 nsew signal input
rlabel metal4 s 185442 0 185502 370 6 um_ow[245]
port 546 nsew signal input
rlabel metal4 s 184706 0 184766 370 6 um_ow[246]
port 547 nsew signal input
rlabel metal4 s 183970 0 184030 370 6 um_ow[247]
port 548 nsew signal input
rlabel metal4 s 183234 0 183294 370 6 um_ow[248]
port 549 nsew signal input
rlabel metal4 s 182498 0 182558 370 6 um_ow[249]
port 550 nsew signal input
rlabel metal4 s 18462 10164 18522 10880 6 um_ow[24]
port 551 nsew signal input
rlabel metal4 s 181762 0 181822 370 6 um_ow[250]
port 552 nsew signal input
rlabel metal4 s 181026 0 181086 370 6 um_ow[251]
port 553 nsew signal input
rlabel metal4 s 180290 0 180350 370 6 um_ow[252]
port 554 nsew signal input
rlabel metal4 s 179554 0 179614 370 6 um_ow[253]
port 555 nsew signal input
rlabel metal4 s 178818 0 178878 370 6 um_ow[254]
port 556 nsew signal input
rlabel metal4 s 178082 0 178142 370 6 um_ow[255]
port 557 nsew signal input
rlabel metal4 s 177346 0 177406 370 6 um_ow[256]
port 558 nsew signal input
rlabel metal4 s 176610 0 176670 370 6 um_ow[257]
port 559 nsew signal input
rlabel metal4 s 175874 0 175934 370 6 um_ow[258]
port 560 nsew signal input
rlabel metal4 s 175138 0 175198 370 6 um_ow[259]
port 561 nsew signal input
rlabel metal4 s 17726 10164 17786 10880 6 um_ow[25]
port 562 nsew signal input
rlabel metal4 s 174402 0 174462 370 6 um_ow[260]
port 563 nsew signal input
rlabel metal4 s 173666 0 173726 370 6 um_ow[261]
port 564 nsew signal input
rlabel metal4 s 172930 0 172990 370 6 um_ow[262]
port 565 nsew signal input
rlabel metal4 s 172194 0 172254 370 6 um_ow[263]
port 566 nsew signal input
rlabel metal4 s 189122 10300 189182 10880 6 um_ow[264]
port 567 nsew signal input
rlabel metal4 s 188386 10300 188446 10880 6 um_ow[265]
port 568 nsew signal input
rlabel metal4 s 187650 10300 187710 10880 6 um_ow[266]
port 569 nsew signal input
rlabel metal4 s 186914 10300 186974 10880 6 um_ow[267]
port 570 nsew signal input
rlabel metal4 s 186178 10300 186238 10880 6 um_ow[268]
port 571 nsew signal input
rlabel metal4 s 185442 10300 185502 10880 6 um_ow[269]
port 572 nsew signal input
rlabel metal4 s 16990 10164 17050 10880 6 um_ow[26]
port 573 nsew signal input
rlabel metal4 s 184706 10300 184766 10880 6 um_ow[270]
port 574 nsew signal input
rlabel metal4 s 183970 10300 184030 10880 6 um_ow[271]
port 575 nsew signal input
rlabel metal4 s 183234 10300 183294 10880 6 um_ow[272]
port 576 nsew signal input
rlabel metal4 s 182498 10300 182558 10880 6 um_ow[273]
port 577 nsew signal input
rlabel metal4 s 181762 10436 181822 10880 6 um_ow[274]
port 578 nsew signal input
rlabel metal4 s 181026 10300 181086 10880 6 um_ow[275]
port 579 nsew signal input
rlabel metal4 s 180290 10300 180350 10880 6 um_ow[276]
port 580 nsew signal input
rlabel metal4 s 179554 10300 179614 10880 6 um_ow[277]
port 581 nsew signal input
rlabel metal4 s 178818 10300 178878 10880 6 um_ow[278]
port 582 nsew signal input
rlabel metal4 s 178082 10300 178142 10880 6 um_ow[279]
port 583 nsew signal input
rlabel metal4 s 16254 10164 16314 10880 6 um_ow[27]
port 584 nsew signal input
rlabel metal4 s 177346 10300 177406 10880 6 um_ow[280]
port 585 nsew signal input
rlabel metal4 s 176610 10300 176670 10880 6 um_ow[281]
port 586 nsew signal input
rlabel metal4 s 175874 10300 175934 10880 6 um_ow[282]
port 587 nsew signal input
rlabel metal4 s 175138 10300 175198 10880 6 um_ow[283]
port 588 nsew signal input
rlabel metal4 s 174402 10300 174462 10880 6 um_ow[284]
port 589 nsew signal input
rlabel metal4 s 173666 10300 173726 10880 6 um_ow[285]
port 590 nsew signal input
rlabel metal4 s 172930 10300 172990 10880 6 um_ow[286]
port 591 nsew signal input
rlabel metal4 s 172194 10300 172254 10880 6 um_ow[287]
port 592 nsew signal input
rlabel metal4 s 223254 0 223314 2756 6 um_ow[288]
port 593 nsew signal input
rlabel metal4 s 222518 0 222578 1260 6 um_ow[289]
port 594 nsew signal input
rlabel metal4 s 15518 10164 15578 10880 6 um_ow[28]
port 595 nsew signal input
rlabel metal4 s 221782 0 221842 308 6 um_ow[290]
port 596 nsew signal input
rlabel metal4 s 221046 0 221106 852 6 um_ow[291]
port 597 nsew signal input
rlabel metal4 s 220310 0 220370 1396 6 um_ow[292]
port 598 nsew signal input
rlabel metal4 s 219574 0 219634 308 6 um_ow[293]
port 599 nsew signal input
rlabel metal4 s 218838 0 218898 308 6 um_ow[294]
port 600 nsew signal input
rlabel metal4 s 218102 0 218162 852 6 um_ow[295]
port 601 nsew signal input
rlabel metal4 s 217366 0 217426 852 6 um_ow[296]
port 602 nsew signal input
rlabel metal4 s 216630 0 216690 1396 6 um_ow[297]
port 603 nsew signal input
rlabel metal4 s 215894 0 215954 852 6 um_ow[298]
port 604 nsew signal input
rlabel metal4 s 215158 0 215218 852 6 um_ow[299]
port 605 nsew signal input
rlabel metal4 s 14782 10164 14842 10880 6 um_ow[29]
port 606 nsew signal input
rlabel metal4 s 16990 0 17050 580 6 um_ow[2]
port 607 nsew signal input
rlabel metal4 s 214422 0 214482 852 6 um_ow[300]
port 608 nsew signal input
rlabel metal4 s 213686 0 213746 852 6 um_ow[301]
port 609 nsew signal input
rlabel metal4 s 212950 0 213010 852 6 um_ow[302]
port 610 nsew signal input
rlabel metal4 s 212214 0 212274 852 6 um_ow[303]
port 611 nsew signal input
rlabel metal4 s 211478 0 211538 988 6 um_ow[304]
port 612 nsew signal input
rlabel metal4 s 210742 0 210802 1260 6 um_ow[305]
port 613 nsew signal input
rlabel metal4 s 210006 0 210066 988 6 um_ow[306]
port 614 nsew signal input
rlabel metal4 s 209270 0 209330 852 6 um_ow[307]
port 615 nsew signal input
rlabel metal4 s 208534 0 208594 852 6 um_ow[308]
port 616 nsew signal input
rlabel metal4 s 207798 0 207858 852 6 um_ow[309]
port 617 nsew signal input
rlabel metal4 s 14046 10164 14106 10880 6 um_ow[30]
port 618 nsew signal input
rlabel metal4 s 207062 0 207122 852 6 um_ow[310]
port 619 nsew signal input
rlabel metal4 s 206326 0 206386 852 6 um_ow[311]
port 620 nsew signal input
rlabel metal4 s 223254 10164 223314 10880 6 um_ow[312]
port 621 nsew signal input
rlabel metal4 s 222518 10300 222578 10880 6 um_ow[313]
port 622 nsew signal input
rlabel metal4 s 221782 10300 221842 10880 6 um_ow[314]
port 623 nsew signal input
rlabel metal4 s 221046 10436 221106 10880 6 um_ow[315]
port 624 nsew signal input
rlabel metal4 s 220310 10300 220370 10880 6 um_ow[316]
port 625 nsew signal input
rlabel metal4 s 219574 10164 219634 10880 6 um_ow[317]
port 626 nsew signal input
rlabel metal4 s 218838 10164 218898 10880 6 um_ow[318]
port 627 nsew signal input
rlabel metal4 s 218102 10572 218162 10880 6 um_ow[319]
port 628 nsew signal input
rlabel metal4 s 13310 9892 13370 10880 6 um_ow[31]
port 629 nsew signal input
rlabel metal4 s 217366 10164 217426 10880 6 um_ow[320]
port 630 nsew signal input
rlabel metal4 s 216630 9892 216690 10880 6 um_ow[321]
port 631 nsew signal input
rlabel metal4 s 215894 10164 215954 10880 6 um_ow[322]
port 632 nsew signal input
rlabel metal4 s 215158 10300 215218 10880 6 um_ow[323]
port 633 nsew signal input
rlabel metal4 s 214422 10164 214482 10880 6 um_ow[324]
port 634 nsew signal input
rlabel metal4 s 213686 10164 213746 10880 6 um_ow[325]
port 635 nsew signal input
rlabel metal4 s 212950 10164 213010 10880 6 um_ow[326]
port 636 nsew signal input
rlabel metal4 s 212214 6900 212274 10880 6 um_ow[327]
port 637 nsew signal input
rlabel metal4 s 211478 10436 211538 10880 6 um_ow[328]
port 638 nsew signal input
rlabel metal4 s 210742 10164 210802 10880 6 um_ow[329]
port 639 nsew signal input
rlabel metal4 s 12574 10164 12634 10880 6 um_ow[32]
port 640 nsew signal input
rlabel metal4 s 210006 10436 210066 10880 6 um_ow[330]
port 641 nsew signal input
rlabel metal4 s 209270 10164 209330 10880 6 um_ow[331]
port 642 nsew signal input
rlabel metal4 s 208534 10164 208594 10880 6 um_ow[332]
port 643 nsew signal input
rlabel metal4 s 207798 10572 207858 10880 6 um_ow[333]
port 644 nsew signal input
rlabel metal4 s 207062 10164 207122 10880 6 um_ow[334]
port 645 nsew signal input
rlabel metal4 s 206326 10164 206386 10880 6 um_ow[335]
port 646 nsew signal input
rlabel metal4 s 257386 0 257446 580 6 um_ow[336]
port 647 nsew signal input
rlabel metal4 s 256650 0 256710 580 6 um_ow[337]
port 648 nsew signal input
rlabel metal4 s 255914 0 255974 580 6 um_ow[338]
port 649 nsew signal input
rlabel metal4 s 255178 0 255238 580 6 um_ow[339]
port 650 nsew signal input
rlabel metal4 s 11838 10164 11898 10880 6 um_ow[33]
port 651 nsew signal input
rlabel metal4 s 254442 0 254502 308 6 um_ow[340]
port 652 nsew signal input
rlabel metal4 s 253706 0 253766 580 6 um_ow[341]
port 653 nsew signal input
rlabel metal4 s 252970 0 253030 580 6 um_ow[342]
port 654 nsew signal input
rlabel metal4 s 252234 0 252294 580 6 um_ow[343]
port 655 nsew signal input
rlabel metal4 s 251498 0 251558 580 6 um_ow[344]
port 656 nsew signal input
rlabel metal4 s 250762 0 250822 370 6 um_ow[345]
port 657 nsew signal input
rlabel metal4 s 250026 0 250086 580 6 um_ow[346]
port 658 nsew signal input
rlabel metal4 s 249290 0 249350 370 6 um_ow[347]
port 659 nsew signal input
rlabel metal4 s 248554 0 248614 444 6 um_ow[348]
port 660 nsew signal input
rlabel metal4 s 247818 0 247878 370 6 um_ow[349]
port 661 nsew signal input
rlabel metal4 s 11102 9892 11162 10880 6 um_ow[34]
port 662 nsew signal input
rlabel metal4 s 247082 0 247142 370 6 um_ow[350]
port 663 nsew signal input
rlabel metal4 s 246346 0 246406 444 6 um_ow[351]
port 664 nsew signal input
rlabel metal4 s 245610 0 245670 444 6 um_ow[352]
port 665 nsew signal input
rlabel metal4 s 244874 0 244934 444 6 um_ow[353]
port 666 nsew signal input
rlabel metal4 s 244138 0 244198 370 6 um_ow[354]
port 667 nsew signal input
rlabel metal4 s 243402 0 243462 444 6 um_ow[355]
port 668 nsew signal input
rlabel metal4 s 242666 0 242726 370 6 um_ow[356]
port 669 nsew signal input
rlabel metal4 s 241930 0 241990 444 6 um_ow[357]
port 670 nsew signal input
rlabel metal4 s 241194 0 241254 444 6 um_ow[358]
port 671 nsew signal input
rlabel metal4 s 240458 0 240518 308 6 um_ow[359]
port 672 nsew signal input
rlabel metal4 s 10366 9892 10426 10880 6 um_ow[35]
port 673 nsew signal input
rlabel metal4 s 257386 10300 257446 10880 6 um_ow[360]
port 674 nsew signal input
rlabel metal4 s 256650 10300 256710 10880 6 um_ow[361]
port 675 nsew signal input
rlabel metal4 s 255914 10300 255974 10880 6 um_ow[362]
port 676 nsew signal input
rlabel metal4 s 255178 10300 255238 10880 6 um_ow[363]
port 677 nsew signal input
rlabel metal4 s 254442 10300 254502 10880 6 um_ow[364]
port 678 nsew signal input
rlabel metal4 s 253706 10300 253766 10880 6 um_ow[365]
port 679 nsew signal input
rlabel metal4 s 252970 10300 253030 10880 6 um_ow[366]
port 680 nsew signal input
rlabel metal4 s 252234 10300 252294 10880 6 um_ow[367]
port 681 nsew signal input
rlabel metal4 s 251498 10300 251558 10880 6 um_ow[368]
port 682 nsew signal input
rlabel metal4 s 250762 10300 250822 10880 6 um_ow[369]
port 683 nsew signal input
rlabel metal4 s 9630 10572 9690 10880 6 um_ow[36]
port 684 nsew signal input
rlabel metal4 s 250026 10300 250086 10880 6 um_ow[370]
port 685 nsew signal input
rlabel metal4 s 249290 10300 249350 10880 6 um_ow[371]
port 686 nsew signal input
rlabel metal4 s 248554 10300 248614 10880 6 um_ow[372]
port 687 nsew signal input
rlabel metal4 s 247818 10300 247878 10880 6 um_ow[373]
port 688 nsew signal input
rlabel metal4 s 247082 10300 247142 10880 6 um_ow[374]
port 689 nsew signal input
rlabel metal4 s 246346 10300 246406 10880 6 um_ow[375]
port 690 nsew signal input
rlabel metal4 s 245610 10300 245670 10880 6 um_ow[376]
port 691 nsew signal input
rlabel metal4 s 244874 10300 244934 10880 6 um_ow[377]
port 692 nsew signal input
rlabel metal4 s 244138 10300 244198 10880 6 um_ow[378]
port 693 nsew signal input
rlabel metal4 s 243402 10300 243462 10880 6 um_ow[379]
port 694 nsew signal input
rlabel metal4 s 8894 10164 8954 10880 6 um_ow[37]
port 695 nsew signal input
rlabel metal4 s 242666 10300 242726 10880 6 um_ow[380]
port 696 nsew signal input
rlabel metal4 s 241930 10300 241990 10880 6 um_ow[381]
port 697 nsew signal input
rlabel metal4 s 241194 10300 241254 10880 6 um_ow[382]
port 698 nsew signal input
rlabel metal4 s 240458 10300 240518 10880 6 um_ow[383]
port 699 nsew signal input
rlabel metal4 s 8158 9892 8218 10880 6 um_ow[38]
port 700 nsew signal input
rlabel metal4 s 7422 10164 7482 10880 6 um_ow[39]
port 701 nsew signal input
rlabel metal4 s 16254 0 16314 1396 6 um_ow[3]
port 702 nsew signal input
rlabel metal4 s 6686 10164 6746 10880 6 um_ow[40]
port 703 nsew signal input
rlabel metal4 s 5950 10164 6010 10880 6 um_ow[41]
port 704 nsew signal input
rlabel metal4 s 5214 10164 5274 10880 6 um_ow[42]
port 705 nsew signal input
rlabel metal4 s 4478 10164 4538 10880 6 um_ow[43]
port 706 nsew signal input
rlabel metal4 s 3742 10164 3802 10880 6 um_ow[44]
port 707 nsew signal input
rlabel metal4 s 3006 9892 3066 10880 6 um_ow[45]
port 708 nsew signal input
rlabel metal4 s 2270 10164 2330 10880 6 um_ow[46]
port 709 nsew signal input
rlabel metal4 s 1534 10164 1594 10880 6 um_ow[47]
port 710 nsew signal input
rlabel metal4 s 52594 0 52654 580 6 um_ow[48]
port 711 nsew signal input
rlabel metal4 s 51858 0 51918 580 6 um_ow[49]
port 712 nsew signal input
rlabel metal4 s 15518 0 15578 716 6 um_ow[4]
port 713 nsew signal input
rlabel metal4 s 51122 0 51182 580 6 um_ow[50]
port 714 nsew signal input
rlabel metal4 s 50386 0 50446 580 6 um_ow[51]
port 715 nsew signal input
rlabel metal4 s 49650 0 49710 580 6 um_ow[52]
port 716 nsew signal input
rlabel metal4 s 48914 0 48974 580 6 um_ow[53]
port 717 nsew signal input
rlabel metal4 s 48178 0 48238 580 6 um_ow[54]
port 718 nsew signal input
rlabel metal4 s 47442 0 47502 580 6 um_ow[55]
port 719 nsew signal input
rlabel metal4 s 46706 0 46766 580 6 um_ow[56]
port 720 nsew signal input
rlabel metal4 s 45970 0 46030 580 6 um_ow[57]
port 721 nsew signal input
rlabel metal4 s 45234 0 45294 580 6 um_ow[58]
port 722 nsew signal input
rlabel metal4 s 44498 0 44558 580 6 um_ow[59]
port 723 nsew signal input
rlabel metal4 s 14782 0 14842 716 6 um_ow[5]
port 724 nsew signal input
rlabel metal4 s 43762 0 43822 580 6 um_ow[60]
port 725 nsew signal input
rlabel metal4 s 43026 0 43086 580 6 um_ow[61]
port 726 nsew signal input
rlabel metal4 s 42290 0 42350 580 6 um_ow[62]
port 727 nsew signal input
rlabel metal4 s 41554 0 41614 580 6 um_ow[63]
port 728 nsew signal input
rlabel metal4 s 40818 0 40878 580 6 um_ow[64]
port 729 nsew signal input
rlabel metal4 s 40082 0 40142 580 6 um_ow[65]
port 730 nsew signal input
rlabel metal4 s 39346 0 39406 308 6 um_ow[66]
port 731 nsew signal input
rlabel metal4 s 38610 0 38670 580 6 um_ow[67]
port 732 nsew signal input
rlabel metal4 s 37874 0 37934 580 6 um_ow[68]
port 733 nsew signal input
rlabel metal4 s 37138 0 37198 580 6 um_ow[69]
port 734 nsew signal input
rlabel metal4 s 14046 0 14106 988 6 um_ow[6]
port 735 nsew signal input
rlabel metal4 s 36402 0 36462 580 6 um_ow[70]
port 736 nsew signal input
rlabel metal4 s 35666 0 35726 580 6 um_ow[71]
port 737 nsew signal input
rlabel metal4 s 52594 10300 52654 10880 6 um_ow[72]
port 738 nsew signal input
rlabel metal4 s 51858 10300 51918 10880 6 um_ow[73]
port 739 nsew signal input
rlabel metal4 s 51122 10300 51182 10880 6 um_ow[74]
port 740 nsew signal input
rlabel metal4 s 50386 10300 50446 10880 6 um_ow[75]
port 741 nsew signal input
rlabel metal4 s 49650 10300 49710 10880 6 um_ow[76]
port 742 nsew signal input
rlabel metal4 s 48914 10300 48974 10880 6 um_ow[77]
port 743 nsew signal input
rlabel metal4 s 48178 10300 48238 10880 6 um_ow[78]
port 744 nsew signal input
rlabel metal4 s 47442 10300 47502 10880 6 um_ow[79]
port 745 nsew signal input
rlabel metal4 s 13310 0 13370 580 6 um_ow[7]
port 746 nsew signal input
rlabel metal4 s 46706 10300 46766 10880 6 um_ow[80]
port 747 nsew signal input
rlabel metal4 s 45970 10300 46030 10880 6 um_ow[81]
port 748 nsew signal input
rlabel metal4 s 45234 10300 45294 10880 6 um_ow[82]
port 749 nsew signal input
rlabel metal4 s 44498 10300 44558 10880 6 um_ow[83]
port 750 nsew signal input
rlabel metal4 s 43762 10300 43822 10880 6 um_ow[84]
port 751 nsew signal input
rlabel metal4 s 43026 10300 43086 10880 6 um_ow[85]
port 752 nsew signal input
rlabel metal4 s 42290 10300 42350 10880 6 um_ow[86]
port 753 nsew signal input
rlabel metal4 s 41554 10300 41614 10880 6 um_ow[87]
port 754 nsew signal input
rlabel metal4 s 40818 10300 40878 10880 6 um_ow[88]
port 755 nsew signal input
rlabel metal4 s 40082 10300 40142 10880 6 um_ow[89]
port 756 nsew signal input
rlabel metal4 s 12574 0 12634 580 6 um_ow[8]
port 757 nsew signal input
rlabel metal4 s 39346 10300 39406 10880 6 um_ow[90]
port 758 nsew signal input
rlabel metal4 s 38610 10300 38670 10880 6 um_ow[91]
port 759 nsew signal input
rlabel metal4 s 37874 10300 37934 10880 6 um_ow[92]
port 760 nsew signal input
rlabel metal4 s 37138 10300 37198 10880 6 um_ow[93]
port 761 nsew signal input
rlabel metal4 s 36402 10300 36462 10880 6 um_ow[94]
port 762 nsew signal input
rlabel metal4 s 35666 10300 35726 10880 6 um_ow[95]
port 763 nsew signal input
rlabel metal4 s 86726 0 86786 716 6 um_ow[96]
port 764 nsew signal input
rlabel metal4 s 85990 0 86050 988 6 um_ow[97]
port 765 nsew signal input
rlabel metal4 s 85254 0 85314 716 6 um_ow[98]
port 766 nsew signal input
rlabel metal4 s 84518 0 84578 716 6 um_ow[99]
port 767 nsew signal input
rlabel metal4 s 11838 0 11898 580 6 um_ow[9]
port 768 nsew signal input
rlabel metal4 s 34742 1040 35062 9840 6 vccd1
port 769 nsew power bidirectional
rlabel metal4 s 102339 1040 102659 9840 6 vccd1
port 769 nsew power bidirectional
rlabel metal4 s 169936 1040 170256 9840 6 vccd1
port 769 nsew power bidirectional
rlabel metal4 s 237533 1040 237853 9840 6 vccd1
port 769 nsew power bidirectional
rlabel metal4 s 68540 1040 68860 9840 6 vssd1
port 770 nsew ground bidirectional
rlabel metal4 s 136137 1040 136457 9840 6 vssd1
port 770 nsew ground bidirectional
rlabel metal4 s 203734 1040 204054 9840 6 vssd1
port 770 nsew ground bidirectional
rlabel metal4 s 271331 1040 271651 9840 6 vssd1
port 770 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 272600 11000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4483126
string GDS_FILE /home/uri/p/tinytapeout-03p5/openlane/tt_mux/runs/23_05_22_20_15/results/signoff/tt_mux.magic.gds
string GDS_START 249434
<< end >>

