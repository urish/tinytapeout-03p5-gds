VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_mux
  CLASS BLOCK ;
  FOREIGN tt_mux ;
  ORIGIN 0.000 0.000 ;
  SIZE 1363.000 BY 55.000 ;
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1360.990 47.790 1362.520 48.090 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1360.070 47.110 1362.520 47.410 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1344.950 46.430 1362.520 46.730 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1340.350 45.750 1362.520 46.050 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1340.810 45.070 1362.520 45.370 ;
    END
  END addr[4]
  PIN k_one
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1360.130 44.390 1362.520 44.690 ;
    END
  END k_one
  PIN k_zero
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1359.150 43.710 1362.520 44.010 ;
    END
  END k_zero
  PIN spine_iw[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1361.520 43.030 1362.520 43.330 ;
    END
  END spine_iw[0]
  PIN spine_iw[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1360.130 36.230 1362.520 36.530 ;
    END
  END spine_iw[10]
  PIN spine_iw[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1312.750 35.550 1362.520 35.850 ;
    END
  END spine_iw[11]
  PIN spine_iw[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1340.350 34.870 1362.520 35.170 ;
    END
  END spine_iw[12]
  PIN spine_iw[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1340.810 34.190 1362.520 34.490 ;
    END
  END spine_iw[13]
  PIN spine_iw[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1360.590 33.510 1362.520 33.810 ;
    END
  END spine_iw[14]
  PIN spine_iw[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1359.670 32.830 1362.520 33.130 ;
    END
  END spine_iw[15]
  PIN spine_iw[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1359.150 32.150 1362.520 32.450 ;
    END
  END spine_iw[16]
  PIN spine_iw[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1360.130 31.470 1362.520 31.770 ;
    END
  END spine_iw[17]
  PIN spine_iw[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1344.950 30.790 1362.520 31.090 ;
    END
  END spine_iw[18]
  PIN spine_iw[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1359.210 30.110 1362.520 30.410 ;
    END
  END spine_iw[19]
  PIN spine_iw[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1353.230 42.350 1362.520 42.650 ;
    END
  END spine_iw[1]
  PIN spine_iw[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1358.750 29.430 1362.520 29.730 ;
    END
  END spine_iw[20]
  PIN spine_iw[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1357.310 28.750 1362.520 29.050 ;
    END
  END spine_iw[21]
  PIN spine_iw[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1356.390 28.070 1362.520 28.370 ;
    END
  END spine_iw[22]
  PIN spine_iw[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1359.210 27.390 1362.520 27.690 ;
    END
  END spine_iw[23]
  PIN spine_iw[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1360.130 26.710 1362.520 27.010 ;
    END
  END spine_iw[24]
  PIN spine_iw[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1344.950 26.030 1362.520 26.330 ;
    END
  END spine_iw[25]
  PIN spine_iw[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1360.130 25.350 1362.520 25.650 ;
    END
  END spine_iw[26]
  PIN spine_iw[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1340.810 24.670 1362.520 24.970 ;
    END
  END spine_iw[27]
  PIN spine_iw[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1344.490 23.990 1362.520 24.290 ;
    END
  END spine_iw[28]
  PIN spine_iw[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1361.050 23.310 1362.520 23.610 ;
    END
  END spine_iw[29]
  PIN spine_iw[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1356.450 41.670 1362.520 41.970 ;
    END
  END spine_iw[2]
  PIN spine_iw[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1361.520 22.630 1362.520 22.930 ;
    END
  END spine_iw[30]
  PIN spine_iw[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1352.770 40.990 1362.520 41.290 ;
    END
  END spine_iw[3]
  PIN spine_iw[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1351.850 40.310 1362.520 40.610 ;
    END
  END spine_iw[4]
  PIN spine_iw[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1350.930 39.630 1362.520 39.930 ;
    END
  END spine_iw[5]
  PIN spine_iw[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1340.350 38.950 1362.520 39.250 ;
    END
  END spine_iw[6]
  PIN spine_iw[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1359.210 38.270 1362.520 38.570 ;
    END
  END spine_iw[7]
  PIN spine_iw[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1359.210 37.590 1362.520 37.890 ;
    END
  END spine_iw[8]
  PIN spine_iw[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1340.350 36.910 1362.520 37.210 ;
    END
  END spine_iw[9]
  PIN spine_ow[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1359.840 21.950 1362.520 22.250 ;
    END
  END spine_ow[0]
  PIN spine_ow[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1311.370 15.150 1362.520 15.450 ;
    END
  END spine_ow[10]
  PIN spine_ow[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1360.130 14.470 1362.520 14.770 ;
    END
  END spine_ow[11]
  PIN spine_ow[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1354.150 13.790 1362.520 14.090 ;
    END
  END spine_ow[12]
  PIN spine_ow[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1336.210 13.110 1362.520 13.410 ;
    END
  END spine_ow[13]
  PIN spine_ow[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1342.650 12.430 1362.520 12.730 ;
    END
  END spine_ow[14]
  PIN spine_ow[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1360.130 11.750 1362.520 12.050 ;
    END
  END spine_ow[15]
  PIN spine_ow[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1359.150 11.070 1362.520 11.370 ;
    END
  END spine_ow[16]
  PIN spine_ow[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1359.210 10.390 1362.520 10.690 ;
    END
  END spine_ow[17]
  PIN spine_ow[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1361.050 9.710 1362.520 10.010 ;
    END
  END spine_ow[18]
  PIN spine_ow[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1350.870 9.030 1362.520 9.330 ;
    END
  END spine_ow[19]
  PIN spine_ow[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1359.150 21.270 1362.520 21.570 ;
    END
  END spine_ow[1]
  PIN spine_ow[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1349.950 8.350 1362.520 8.650 ;
    END
  END spine_ow[20]
  PIN spine_ow[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1345.410 7.670 1362.520 7.970 ;
    END
  END spine_ow[21]
  PIN spine_ow[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1344.490 6.990 1362.520 7.290 ;
    END
  END spine_ow[22]
  PIN spine_ow[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1344.430 6.310 1362.520 6.610 ;
    END
  END spine_ow[23]
  PIN spine_ow[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1359.210 5.630 1362.520 5.930 ;
    END
  END spine_ow[24]
  PIN spine_ow[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1359.150 4.950 1362.520 5.250 ;
    END
  END spine_ow[25]
  PIN spine_ow[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1221.210 20.590 1362.520 20.890 ;
    END
  END spine_ow[2]
  PIN spine_ow[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1356.390 19.910 1362.520 20.210 ;
    END
  END spine_ow[3]
  PIN spine_ow[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1357.310 19.230 1362.520 19.530 ;
    END
  END spine_ow[4]
  PIN spine_ow[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1358.290 18.550 1362.520 18.850 ;
    END
  END spine_ow[5]
  PIN spine_ow[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1339.890 17.870 1362.520 18.170 ;
    END
  END spine_ow[6]
  PIN spine_ow[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1360.130 17.190 1362.520 17.490 ;
    END
  END spine_ow[7]
  PIN spine_ow[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1359.150 16.510 1362.520 16.810 ;
    END
  END spine_ow[8]
  PIN spine_ow[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1359.210 15.830 1362.520 16.130 ;
    END
  END spine_ow[9]
  PIN um_ena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 162.230 0.000 162.530 6.980 ;
    END
  END um_ena[0]
  PIN um_ena[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1015.530 0.000 1015.830 1.850 ;
    END
  END um_ena[10]
  PIN um_ena[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1015.530 51.500 1015.830 54.400 ;
    END
  END um_ena[11]
  PIN um_ena[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1186.190 0.000 1186.490 6.980 ;
    END
  END um_ena[12]
  PIN um_ena[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1186.190 46.060 1186.490 54.400 ;
    END
  END um_ena[13]
  PIN um_ena[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1356.850 0.000 1357.150 1.540 ;
    END
  END um_ena[14]
  PIN um_ena[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1356.850 51.190 1357.150 54.400 ;
    END
  END um_ena[15]
  PIN um_ena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 162.230 48.100 162.530 54.400 ;
    END
  END um_ena[1]
  PIN um_ena[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 332.890 0.000 333.190 2.220 ;
    END
  END um_ena[2]
  PIN um_ena[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 332.890 51.500 333.190 54.400 ;
    END
  END um_ena[3]
  PIN um_ena[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 503.550 0.000 503.850 4.260 ;
    END
  END um_ena[4]
  PIN um_ena[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 503.550 48.780 503.850 54.400 ;
    END
  END um_ena[5]
  PIN um_ena[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 674.210 0.000 674.510 1.850 ;
    END
  END um_ena[6]
  PIN um_ena[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 674.210 51.500 674.510 54.400 ;
    END
  END um_ena[7]
  PIN um_ena[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 844.870 0.000 845.170 2.900 ;
    END
  END um_ena[8]
  PIN um_ena[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 844.870 46.060 845.170 54.400 ;
    END
  END um_ena[9]
  PIN um_iw[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 0.000 158.850 2.220 ;
    END
  END um_iw[0]
  PIN um_iw[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 463.070 41.980 463.370 54.400 ;
    END
  END um_iw[100]
  PIN um_iw[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 459.390 43.340 459.690 54.400 ;
    END
  END um_iw[101]
  PIN um_iw[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 455.710 44.020 456.010 54.400 ;
    END
  END um_iw[102]
  PIN um_iw[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 452.030 43.340 452.330 54.400 ;
    END
  END um_iw[103]
  PIN um_iw[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 448.350 51.500 448.650 54.400 ;
    END
  END um_iw[104]
  PIN um_iw[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 444.670 40.620 444.970 54.400 ;
    END
  END um_iw[105]
  PIN um_iw[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 440.990 46.060 441.290 54.400 ;
    END
  END um_iw[106]
  PIN um_iw[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 437.310 43.340 437.610 54.400 ;
    END
  END um_iw[107]
  PIN um_iw[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 670.530 0.000 670.830 2.900 ;
    END
  END um_iw[108]
  PIN um_iw[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 666.850 0.000 667.150 2.900 ;
    END
  END um_iw[109]
  PIN um_iw[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 0.000 122.050 16.500 ;
    END
  END um_iw[10]
  PIN um_iw[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 663.170 0.000 663.470 2.900 ;
    END
  END um_iw[110]
  PIN um_iw[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 659.490 0.000 659.790 2.900 ;
    END
  END um_iw[111]
  PIN um_iw[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 655.810 0.000 656.110 2.900 ;
    END
  END um_iw[112]
  PIN um_iw[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 652.130 0.000 652.430 1.540 ;
    END
  END um_iw[113]
  PIN um_iw[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 648.450 0.000 648.750 2.900 ;
    END
  END um_iw[114]
  PIN um_iw[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 644.770 0.000 645.070 2.900 ;
    END
  END um_iw[115]
  PIN um_iw[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 641.090 0.000 641.390 1.850 ;
    END
  END um_iw[116]
  PIN um_iw[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 637.410 0.000 637.710 2.900 ;
    END
  END um_iw[117]
  PIN um_iw[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 633.730 0.000 634.030 2.900 ;
    END
  END um_iw[118]
  PIN um_iw[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 630.050 0.000 630.350 2.900 ;
    END
  END um_iw[119]
  PIN um_iw[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 0.000 118.370 2.900 ;
    END
  END um_iw[11]
  PIN um_iw[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 626.370 0.000 626.670 2.900 ;
    END
  END um_iw[120]
  PIN um_iw[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 622.690 0.000 622.990 2.900 ;
    END
  END um_iw[121]
  PIN um_iw[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 619.010 0.000 619.310 2.900 ;
    END
  END um_iw[122]
  PIN um_iw[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 615.330 0.000 615.630 2.900 ;
    END
  END um_iw[123]
  PIN um_iw[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 611.650 0.000 611.950 2.900 ;
    END
  END um_iw[124]
  PIN um_iw[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 607.970 0.000 608.270 2.900 ;
    END
  END um_iw[125]
  PIN um_iw[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 670.530 51.500 670.830 54.400 ;
    END
  END um_iw[126]
  PIN um_iw[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 666.850 51.500 667.150 54.400 ;
    END
  END um_iw[127]
  PIN um_iw[128]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 663.170 51.500 663.470 54.400 ;
    END
  END um_iw[128]
  PIN um_iw[129]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 659.490 51.500 659.790 54.400 ;
    END
  END um_iw[129]
  PIN um_iw[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 0.000 114.690 14.460 ;
    END
  END um_iw[12]
  PIN um_iw[130]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 655.810 51.500 656.110 54.400 ;
    END
  END um_iw[130]
  PIN um_iw[131]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 652.130 51.500 652.430 54.400 ;
    END
  END um_iw[131]
  PIN um_iw[132]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 648.450 51.500 648.750 54.400 ;
    END
  END um_iw[132]
  PIN um_iw[133]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 644.770 51.500 645.070 54.400 ;
    END
  END um_iw[133]
  PIN um_iw[134]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 641.090 52.180 641.390 54.400 ;
    END
  END um_iw[134]
  PIN um_iw[135]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 637.410 51.500 637.710 54.400 ;
    END
  END um_iw[135]
  PIN um_iw[136]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 633.730 51.500 634.030 54.400 ;
    END
  END um_iw[136]
  PIN um_iw[137]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 630.050 51.500 630.350 54.400 ;
    END
  END um_iw[137]
  PIN um_iw[138]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 626.370 52.180 626.670 54.400 ;
    END
  END um_iw[138]
  PIN um_iw[139]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 622.690 51.500 622.990 54.400 ;
    END
  END um_iw[139]
  PIN um_iw[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 0.000 111.010 13.780 ;
    END
  END um_iw[13]
  PIN um_iw[140]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 619.010 51.500 619.310 54.400 ;
    END
  END um_iw[140]
  PIN um_iw[141]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 615.330 51.500 615.630 54.400 ;
    END
  END um_iw[141]
  PIN um_iw[142]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 611.650 51.500 611.950 54.400 ;
    END
  END um_iw[142]
  PIN um_iw[143]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 607.970 51.500 608.270 54.400 ;
    END
  END um_iw[143]
  PIN um_iw[144]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 841.190 0.000 841.490 6.980 ;
    END
  END um_iw[144]
  PIN um_iw[145]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 837.510 0.000 837.810 2.900 ;
    END
  END um_iw[145]
  PIN um_iw[146]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 833.830 0.000 834.130 5.620 ;
    END
  END um_iw[146]
  PIN um_iw[147]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 830.150 0.000 830.450 5.620 ;
    END
  END um_iw[147]
  PIN um_iw[148]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 826.470 0.000 826.770 5.620 ;
    END
  END um_iw[148]
  PIN um_iw[149]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 822.790 0.000 823.090 2.900 ;
    END
  END um_iw[149]
  PIN um_iw[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 0.000 107.330 8.340 ;
    END
  END um_iw[14]
  PIN um_iw[150]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 819.110 0.000 819.410 6.980 ;
    END
  END um_iw[150]
  PIN um_iw[151]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 815.430 0.000 815.730 5.620 ;
    END
  END um_iw[151]
  PIN um_iw[152]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 811.750 0.000 812.050 2.900 ;
    END
  END um_iw[152]
  PIN um_iw[153]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 808.070 0.000 808.370 5.620 ;
    END
  END um_iw[153]
  PIN um_iw[154]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 804.390 0.000 804.690 2.900 ;
    END
  END um_iw[154]
  PIN um_iw[155]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 800.710 0.000 801.010 5.620 ;
    END
  END um_iw[155]
  PIN um_iw[156]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 797.030 0.000 797.330 13.780 ;
    END
  END um_iw[156]
  PIN um_iw[157]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 793.350 0.000 793.650 2.900 ;
    END
  END um_iw[157]
  PIN um_iw[158]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 789.670 0.000 789.970 6.980 ;
    END
  END um_iw[158]
  PIN um_iw[159]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 785.990 0.000 786.290 13.780 ;
    END
  END um_iw[159]
  PIN um_iw[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 0.000 103.650 6.980 ;
    END
  END um_iw[15]
  PIN um_iw[160]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 782.310 0.000 782.610 6.980 ;
    END
  END um_iw[160]
  PIN um_iw[161]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 778.630 0.000 778.930 6.980 ;
    END
  END um_iw[161]
  PIN um_iw[162]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 841.190 40.620 841.490 54.400 ;
    END
  END um_iw[162]
  PIN um_iw[163]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 837.510 41.980 837.810 54.400 ;
    END
  END um_iw[163]
  PIN um_iw[164]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 833.830 41.300 834.130 54.400 ;
    END
  END um_iw[164]
  PIN um_iw[165]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 830.150 41.980 830.450 54.400 ;
    END
  END um_iw[165]
  PIN um_iw[166]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 826.470 41.980 826.770 54.400 ;
    END
  END um_iw[166]
  PIN um_iw[167]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 822.790 41.980 823.090 54.400 ;
    END
  END um_iw[167]
  PIN um_iw[168]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 819.110 48.780 819.410 54.400 ;
    END
  END um_iw[168]
  PIN um_iw[169]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 815.430 41.980 815.730 54.400 ;
    END
  END um_iw[169]
  PIN um_iw[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 0.000 99.970 13.780 ;
    END
  END um_iw[16]
  PIN um_iw[170]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 811.750 41.980 812.050 54.400 ;
    END
  END um_iw[170]
  PIN um_iw[171]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 808.070 42.660 808.370 54.400 ;
    END
  END um_iw[171]
  PIN um_iw[172]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 804.390 41.980 804.690 54.400 ;
    END
  END um_iw[172]
  PIN um_iw[173]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 800.710 41.980 801.010 54.400 ;
    END
  END um_iw[173]
  PIN um_iw[174]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 797.030 48.780 797.330 54.400 ;
    END
  END um_iw[174]
  PIN um_iw[175]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 793.350 47.420 793.650 54.400 ;
    END
  END um_iw[175]
  PIN um_iw[176]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 789.670 48.780 789.970 54.400 ;
    END
  END um_iw[176]
  PIN um_iw[177]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 785.990 51.500 786.290 54.400 ;
    END
  END um_iw[177]
  PIN um_iw[178]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 782.310 48.780 782.610 54.400 ;
    END
  END um_iw[178]
  PIN um_iw[179]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 778.630 48.780 778.930 54.400 ;
    END
  END um_iw[179]
  PIN um_iw[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 0.000 96.290 14.460 ;
    END
  END um_iw[17]
  PIN um_iw[180]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1011.850 0.000 1012.150 1.850 ;
    END
  END um_iw[180]
  PIN um_iw[181]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1008.170 0.000 1008.470 1.850 ;
    END
  END um_iw[181]
  PIN um_iw[182]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1004.490 0.000 1004.790 1.850 ;
    END
  END um_iw[182]
  PIN um_iw[183]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1000.810 0.000 1001.110 1.850 ;
    END
  END um_iw[183]
  PIN um_iw[184]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 997.130 0.000 997.430 1.850 ;
    END
  END um_iw[184]
  PIN um_iw[185]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 993.450 0.000 993.750 1.850 ;
    END
  END um_iw[185]
  PIN um_iw[186]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 989.770 0.000 990.070 1.850 ;
    END
  END um_iw[186]
  PIN um_iw[187]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 986.090 0.000 986.390 1.850 ;
    END
  END um_iw[187]
  PIN um_iw[188]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 982.410 0.000 982.710 1.850 ;
    END
  END um_iw[188]
  PIN um_iw[189]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 978.730 0.000 979.030 1.850 ;
    END
  END um_iw[189]
  PIN um_iw[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 51.500 158.850 54.400 ;
    END
  END um_iw[18]
  PIN um_iw[190]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 975.050 0.000 975.350 1.850 ;
    END
  END um_iw[190]
  PIN um_iw[191]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 971.370 0.000 971.670 1.850 ;
    END
  END um_iw[191]
  PIN um_iw[192]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 967.690 0.000 967.990 1.850 ;
    END
  END um_iw[192]
  PIN um_iw[193]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 964.010 0.000 964.310 1.850 ;
    END
  END um_iw[193]
  PIN um_iw[194]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 960.330 0.000 960.630 1.850 ;
    END
  END um_iw[194]
  PIN um_iw[195]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 956.650 0.000 956.950 1.850 ;
    END
  END um_iw[195]
  PIN um_iw[196]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 952.970 0.000 953.270 1.850 ;
    END
  END um_iw[196]
  PIN um_iw[197]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 949.290 0.000 949.590 1.850 ;
    END
  END um_iw[197]
  PIN um_iw[198]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1011.850 52.180 1012.150 54.400 ;
    END
  END um_iw[198]
  PIN um_iw[199]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1008.170 51.500 1008.470 54.400 ;
    END
  END um_iw[199]
  PIN um_iw[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 43.340 155.170 54.400 ;
    END
  END um_iw[19]
  PIN um_iw[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 0.000 155.170 1.540 ;
    END
  END um_iw[1]
  PIN um_iw[200]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1004.490 52.180 1004.790 54.400 ;
    END
  END um_iw[200]
  PIN um_iw[201]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1000.810 51.500 1001.110 54.400 ;
    END
  END um_iw[201]
  PIN um_iw[202]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 997.130 51.500 997.430 54.400 ;
    END
  END um_iw[202]
  PIN um_iw[203]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 993.450 52.180 993.750 54.400 ;
    END
  END um_iw[203]
  PIN um_iw[204]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 989.770 51.500 990.070 54.400 ;
    END
  END um_iw[204]
  PIN um_iw[205]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 986.090 51.500 986.390 54.400 ;
    END
  END um_iw[205]
  PIN um_iw[206]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 982.410 51.500 982.710 54.400 ;
    END
  END um_iw[206]
  PIN um_iw[207]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 978.730 51.500 979.030 54.400 ;
    END
  END um_iw[207]
  PIN um_iw[208]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 975.050 51.500 975.350 54.400 ;
    END
  END um_iw[208]
  PIN um_iw[209]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 971.370 51.500 971.670 54.400 ;
    END
  END um_iw[209]
  PIN um_iw[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 43.340 151.490 54.400 ;
    END
  END um_iw[20]
  PIN um_iw[210]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 967.690 52.180 967.990 54.400 ;
    END
  END um_iw[210]
  PIN um_iw[211]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 964.010 51.500 964.310 54.400 ;
    END
  END um_iw[211]
  PIN um_iw[212]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 960.330 51.500 960.630 54.400 ;
    END
  END um_iw[212]
  PIN um_iw[213]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 956.650 51.500 956.950 54.400 ;
    END
  END um_iw[213]
  PIN um_iw[214]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 952.970 52.180 953.270 54.400 ;
    END
  END um_iw[214]
  PIN um_iw[215]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 949.290 51.500 949.590 54.400 ;
    END
  END um_iw[215]
  PIN um_iw[216]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1182.510 0.000 1182.810 5.620 ;
    END
  END um_iw[216]
  PIN um_iw[217]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1178.830 0.000 1179.130 13.780 ;
    END
  END um_iw[217]
  PIN um_iw[218]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1175.150 0.000 1175.450 2.220 ;
    END
  END um_iw[218]
  PIN um_iw[219]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1171.470 0.000 1171.770 1.540 ;
    END
  END um_iw[219]
  PIN um_iw[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 43.340 147.810 54.400 ;
    END
  END um_iw[21]
  PIN um_iw[220]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1167.790 0.000 1168.090 1.540 ;
    END
  END um_iw[220]
  PIN um_iw[221]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1164.110 0.000 1164.410 5.620 ;
    END
  END um_iw[221]
  PIN um_iw[222]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1160.430 0.000 1160.730 5.620 ;
    END
  END um_iw[222]
  PIN um_iw[223]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1156.750 0.000 1157.050 5.620 ;
    END
  END um_iw[223]
  PIN um_iw[224]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1153.070 0.000 1153.370 1.540 ;
    END
  END um_iw[224]
  PIN um_iw[225]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1149.390 0.000 1149.690 1.540 ;
    END
  END um_iw[225]
  PIN um_iw[226]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1145.710 0.000 1146.010 1.540 ;
    END
  END um_iw[226]
  PIN um_iw[227]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1142.030 0.000 1142.330 5.620 ;
    END
  END um_iw[227]
  PIN um_iw[228]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1138.350 0.000 1138.650 6.300 ;
    END
  END um_iw[228]
  PIN um_iw[229]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1134.670 0.000 1134.970 6.300 ;
    END
  END um_iw[229]
  PIN um_iw[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 47.420 144.130 54.400 ;
    END
  END um_iw[22]
  PIN um_iw[230]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1130.990 0.000 1131.290 13.780 ;
    END
  END um_iw[230]
  PIN um_iw[231]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1127.310 0.000 1127.610 6.980 ;
    END
  END um_iw[231]
  PIN um_iw[232]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1123.630 0.000 1123.930 13.780 ;
    END
  END um_iw[232]
  PIN um_iw[233]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1119.950 0.000 1120.250 6.980 ;
    END
  END um_iw[233]
  PIN um_iw[234]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1182.510 43.340 1182.810 54.400 ;
    END
  END um_iw[234]
  PIN um_iw[235]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1178.830 46.060 1179.130 54.400 ;
    END
  END um_iw[235]
  PIN um_iw[236]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1175.150 48.780 1175.450 54.400 ;
    END
  END um_iw[236]
  PIN um_iw[237]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1171.470 48.780 1171.770 54.400 ;
    END
  END um_iw[237]
  PIN um_iw[238]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1167.790 48.780 1168.090 54.400 ;
    END
  END um_iw[238]
  PIN um_iw[239]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1164.110 43.340 1164.410 54.400 ;
    END
  END um_iw[239]
  PIN um_iw[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 41.980 140.450 54.400 ;
    END
  END um_iw[23]
  PIN um_iw[240]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1160.430 43.340 1160.730 54.400 ;
    END
  END um_iw[240]
  PIN um_iw[241]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1156.750 48.780 1157.050 54.400 ;
    END
  END um_iw[241]
  PIN um_iw[242]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1153.070 41.980 1153.370 54.400 ;
    END
  END um_iw[242]
  PIN um_iw[243]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1149.390 48.780 1149.690 54.400 ;
    END
  END um_iw[243]
  PIN um_iw[244]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1145.710 43.340 1146.010 54.400 ;
    END
  END um_iw[244]
  PIN um_iw[245]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1142.030 47.420 1142.330 54.400 ;
    END
  END um_iw[245]
  PIN um_iw[246]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1138.350 43.340 1138.650 54.400 ;
    END
  END um_iw[246]
  PIN um_iw[247]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1134.670 43.340 1134.970 54.400 ;
    END
  END um_iw[247]
  PIN um_iw[248]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1130.990 43.340 1131.290 54.400 ;
    END
  END um_iw[248]
  PIN um_iw[249]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1127.310 48.780 1127.610 54.400 ;
    END
  END um_iw[249]
  PIN um_iw[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 39.260 136.770 54.400 ;
    END
  END um_iw[24]
  PIN um_iw[250]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1123.630 41.980 1123.930 54.400 ;
    END
  END um_iw[250]
  PIN um_iw[251]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1119.950 46.060 1120.250 54.400 ;
    END
  END um_iw[251]
  PIN um_iw[252]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1353.170 0.000 1353.470 1.850 ;
    END
  END um_iw[252]
  PIN um_iw[253]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1349.490 0.000 1349.790 2.900 ;
    END
  END um_iw[253]
  PIN um_iw[254]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1345.810 0.000 1346.110 2.220 ;
    END
  END um_iw[254]
  PIN um_iw[255]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1342.130 0.000 1342.430 2.900 ;
    END
  END um_iw[255]
  PIN um_iw[256]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1338.450 0.000 1338.750 2.900 ;
    END
  END um_iw[256]
  PIN um_iw[257]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1334.770 0.000 1335.070 2.900 ;
    END
  END um_iw[257]
  PIN um_iw[258]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1331.090 0.000 1331.390 2.900 ;
    END
  END um_iw[258]
  PIN um_iw[259]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1327.410 0.000 1327.710 2.900 ;
    END
  END um_iw[259]
  PIN um_iw[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 41.980 133.090 54.400 ;
    END
  END um_iw[25]
  PIN um_iw[260]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1323.730 0.000 1324.030 1.850 ;
    END
  END um_iw[260]
  PIN um_iw[261]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1320.050 0.000 1320.350 2.900 ;
    END
  END um_iw[261]
  PIN um_iw[262]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1316.370 0.000 1316.670 2.900 ;
    END
  END um_iw[262]
  PIN um_iw[263]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1312.690 0.000 1312.990 2.900 ;
    END
  END um_iw[263]
  PIN um_iw[264]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1309.010 0.000 1309.310 2.220 ;
    END
  END um_iw[264]
  PIN um_iw[265]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1305.330 0.000 1305.630 2.900 ;
    END
  END um_iw[265]
  PIN um_iw[266]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1301.650 0.000 1301.950 2.900 ;
    END
  END um_iw[266]
  PIN um_iw[267]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1297.970 0.000 1298.270 2.900 ;
    END
  END um_iw[267]
  PIN um_iw[268]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1294.290 0.000 1294.590 2.900 ;
    END
  END um_iw[268]
  PIN um_iw[269]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1290.610 0.000 1290.910 3.210 ;
    END
  END um_iw[269]
  PIN um_iw[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 48.100 129.410 54.400 ;
    END
  END um_iw[26]
  PIN um_iw[270]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1353.170 51.190 1353.470 54.400 ;
    END
  END um_iw[270]
  PIN um_iw[271]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1349.490 51.190 1349.790 54.400 ;
    END
  END um_iw[271]
  PIN um_iw[272]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1345.810 51.190 1346.110 54.400 ;
    END
  END um_iw[272]
  PIN um_iw[273]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1342.130 51.190 1342.430 54.400 ;
    END
  END um_iw[273]
  PIN um_iw[274]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1338.450 51.190 1338.750 54.400 ;
    END
  END um_iw[274]
  PIN um_iw[275]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1334.770 51.190 1335.070 54.400 ;
    END
  END um_iw[275]
  PIN um_iw[276]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1331.090 52.550 1331.390 54.400 ;
    END
  END um_iw[276]
  PIN um_iw[277]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1327.410 51.500 1327.710 54.400 ;
    END
  END um_iw[277]
  PIN um_iw[278]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1323.730 52.180 1324.030 54.400 ;
    END
  END um_iw[278]
  PIN um_iw[279]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1320.050 51.500 1320.350 54.400 ;
    END
  END um_iw[279]
  PIN um_iw[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 34.500 125.730 54.400 ;
    END
  END um_iw[27]
  PIN um_iw[280]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1316.370 51.500 1316.670 54.400 ;
    END
  END um_iw[280]
  PIN um_iw[281]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1312.690 51.500 1312.990 54.400 ;
    END
  END um_iw[281]
  PIN um_iw[282]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1309.010 51.500 1309.310 54.400 ;
    END
  END um_iw[282]
  PIN um_iw[283]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1305.330 52.180 1305.630 54.400 ;
    END
  END um_iw[283]
  PIN um_iw[284]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1301.650 51.500 1301.950 54.400 ;
    END
  END um_iw[284]
  PIN um_iw[285]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1297.970 51.500 1298.270 54.400 ;
    END
  END um_iw[285]
  PIN um_iw[286]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1294.290 51.500 1294.590 54.400 ;
    END
  END um_iw[286]
  PIN um_iw[287]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1290.610 51.500 1290.910 54.400 ;
    END
  END um_iw[287]
  PIN um_iw[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 43.340 122.050 54.400 ;
    END
  END um_iw[28]
  PIN um_iw[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 34.500 118.370 54.400 ;
    END
  END um_iw[29]
  PIN um_iw[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 0.000 151.490 2.900 ;
    END
  END um_iw[2]
  PIN um_iw[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 34.500 114.690 54.400 ;
    END
  END um_iw[30]
  PIN um_iw[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 50.820 111.010 54.400 ;
    END
  END um_iw[31]
  PIN um_iw[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 49.460 107.330 54.400 ;
    END
  END um_iw[32]
  PIN um_iw[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 52.860 103.650 54.400 ;
    END
  END um_iw[33]
  PIN um_iw[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 34.500 99.970 54.400 ;
    END
  END um_iw[34]
  PIN um_iw[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 34.500 96.290 54.400 ;
    END
  END um_iw[35]
  PIN um_iw[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 329.210 0.000 329.510 2.220 ;
    END
  END um_iw[36]
  PIN um_iw[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 325.530 0.000 325.830 2.900 ;
    END
  END um_iw[37]
  PIN um_iw[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 321.850 0.000 322.150 2.900 ;
    END
  END um_iw[38]
  PIN um_iw[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 318.170 0.000 318.470 2.900 ;
    END
  END um_iw[39]
  PIN um_iw[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 0.000 147.810 2.220 ;
    END
  END um_iw[3]
  PIN um_iw[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 314.490 0.000 314.790 2.900 ;
    END
  END um_iw[40]
  PIN um_iw[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 310.810 0.000 311.110 2.900 ;
    END
  END um_iw[41]
  PIN um_iw[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 307.130 0.000 307.430 2.900 ;
    END
  END um_iw[42]
  PIN um_iw[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 303.450 0.000 303.750 2.900 ;
    END
  END um_iw[43]
  PIN um_iw[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 299.770 0.000 300.070 1.850 ;
    END
  END um_iw[44]
  PIN um_iw[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 296.090 0.000 296.390 1.850 ;
    END
  END um_iw[45]
  PIN um_iw[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 292.410 0.000 292.710 2.900 ;
    END
  END um_iw[46]
  PIN um_iw[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 288.730 0.000 289.030 2.900 ;
    END
  END um_iw[47]
  PIN um_iw[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 285.050 0.000 285.350 2.900 ;
    END
  END um_iw[48]
  PIN um_iw[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 281.370 0.000 281.670 2.900 ;
    END
  END um_iw[49]
  PIN um_iw[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 0.000 144.130 2.900 ;
    END
  END um_iw[4]
  PIN um_iw[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 277.690 0.000 277.990 2.900 ;
    END
  END um_iw[50]
  PIN um_iw[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 274.010 0.000 274.310 2.900 ;
    END
  END um_iw[51]
  PIN um_iw[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 270.330 0.000 270.630 1.850 ;
    END
  END um_iw[52]
  PIN um_iw[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 266.650 0.000 266.950 2.900 ;
    END
  END um_iw[53]
  PIN um_iw[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 329.210 51.500 329.510 54.400 ;
    END
  END um_iw[54]
  PIN um_iw[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 325.530 51.500 325.830 54.400 ;
    END
  END um_iw[55]
  PIN um_iw[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 321.850 51.500 322.150 54.400 ;
    END
  END um_iw[56]
  PIN um_iw[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 318.170 51.500 318.470 54.400 ;
    END
  END um_iw[57]
  PIN um_iw[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 314.490 51.500 314.790 54.400 ;
    END
  END um_iw[58]
  PIN um_iw[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 310.810 51.500 311.110 54.400 ;
    END
  END um_iw[59]
  PIN um_iw[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 0.000 140.450 2.220 ;
    END
  END um_iw[5]
  PIN um_iw[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 307.130 51.500 307.430 54.400 ;
    END
  END um_iw[60]
  PIN um_iw[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 303.450 51.500 303.750 54.400 ;
    END
  END um_iw[61]
  PIN um_iw[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 299.770 51.500 300.070 54.400 ;
    END
  END um_iw[62]
  PIN um_iw[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 296.090 51.500 296.390 54.400 ;
    END
  END um_iw[63]
  PIN um_iw[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 292.410 51.500 292.710 54.400 ;
    END
  END um_iw[64]
  PIN um_iw[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 288.730 51.500 289.030 54.400 ;
    END
  END um_iw[65]
  PIN um_iw[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 285.050 51.500 285.350 54.400 ;
    END
  END um_iw[66]
  PIN um_iw[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 281.370 51.500 281.670 54.400 ;
    END
  END um_iw[67]
  PIN um_iw[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 277.690 51.500 277.990 54.400 ;
    END
  END um_iw[68]
  PIN um_iw[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 274.010 51.500 274.310 54.400 ;
    END
  END um_iw[69]
  PIN um_iw[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 0.000 136.770 6.300 ;
    END
  END um_iw[6]
  PIN um_iw[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 270.330 52.180 270.630 54.400 ;
    END
  END um_iw[70]
  PIN um_iw[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 266.650 51.500 266.950 54.400 ;
    END
  END um_iw[71]
  PIN um_iw[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 499.870 0.000 500.170 2.220 ;
    END
  END um_iw[72]
  PIN um_iw[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 496.190 0.000 496.490 7.660 ;
    END
  END um_iw[73]
  PIN um_iw[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 492.510 0.000 492.810 3.580 ;
    END
  END um_iw[74]
  PIN um_iw[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 488.830 0.000 489.130 3.580 ;
    END
  END um_iw[75]
  PIN um_iw[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 485.150 0.000 485.450 2.220 ;
    END
  END um_iw[76]
  PIN um_iw[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 481.470 0.000 481.770 5.620 ;
    END
  END um_iw[77]
  PIN um_iw[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 477.790 0.000 478.090 5.620 ;
    END
  END um_iw[78]
  PIN um_iw[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 474.110 0.000 474.410 5.620 ;
    END
  END um_iw[79]
  PIN um_iw[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 0.000 133.090 6.300 ;
    END
  END um_iw[7]
  PIN um_iw[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 470.430 0.000 470.730 5.620 ;
    END
  END um_iw[80]
  PIN um_iw[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 466.750 0.000 467.050 3.580 ;
    END
  END um_iw[81]
  PIN um_iw[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 463.070 0.000 463.370 1.540 ;
    END
  END um_iw[82]
  PIN um_iw[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 459.390 0.000 459.690 3.580 ;
    END
  END um_iw[83]
  PIN um_iw[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 455.710 0.000 456.010 1.540 ;
    END
  END um_iw[84]
  PIN um_iw[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 452.030 0.000 452.330 3.580 ;
    END
  END um_iw[85]
  PIN um_iw[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 448.350 0.000 448.650 1.540 ;
    END
  END um_iw[86]
  PIN um_iw[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 444.670 0.000 444.970 6.300 ;
    END
  END um_iw[87]
  PIN um_iw[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 440.990 0.000 441.290 5.620 ;
    END
  END um_iw[88]
  PIN um_iw[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 437.310 0.000 437.610 6.300 ;
    END
  END um_iw[89]
  PIN um_iw[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 0.000 129.410 6.300 ;
    END
  END um_iw[8]
  PIN um_iw[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 499.870 43.340 500.170 54.400 ;
    END
  END um_iw[90]
  PIN um_iw[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 496.190 41.300 496.490 54.400 ;
    END
  END um_iw[91]
  PIN um_iw[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 492.510 43.340 492.810 54.400 ;
    END
  END um_iw[92]
  PIN um_iw[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 488.830 48.780 489.130 54.400 ;
    END
  END um_iw[93]
  PIN um_iw[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 485.150 43.340 485.450 54.400 ;
    END
  END um_iw[94]
  PIN um_iw[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 481.470 48.780 481.770 54.400 ;
    END
  END um_iw[95]
  PIN um_iw[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 477.790 48.780 478.090 54.400 ;
    END
  END um_iw[96]
  PIN um_iw[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 474.110 43.340 474.410 54.400 ;
    END
  END um_iw[97]
  PIN um_iw[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 470.430 43.340 470.730 54.400 ;
    END
  END um_iw[98]
  PIN um_iw[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 466.750 48.780 467.050 54.400 ;
    END
  END um_iw[99]
  PIN um_iw[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 0.000 125.730 13.780 ;
    END
  END um_iw[9]
  PIN um_k_zero[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 0.000 4.290 6.980 ;
    END
  END um_k_zero[0]
  PIN um_k_zero[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 857.290 0.000 857.590 1.850 ;
    END
  END um_k_zero[10]
  PIN um_k_zero[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 857.290 51.500 857.590 54.400 ;
    END
  END um_k_zero[11]
  PIN um_k_zero[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1027.950 0.000 1028.250 1.850 ;
    END
  END um_k_zero[12]
  PIN um_k_zero[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1027.950 48.100 1028.250 54.400 ;
    END
  END um_k_zero[13]
  PIN um_k_zero[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1198.610 0.000 1198.910 1.540 ;
    END
  END um_k_zero[14]
  PIN um_k_zero[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1198.610 51.500 1198.910 54.400 ;
    END
  END um_k_zero[15]
  PIN um_k_zero[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 46.060 4.290 54.400 ;
    END
  END um_k_zero[1]
  PIN um_k_zero[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 174.650 0.000 174.950 1.540 ;
    END
  END um_k_zero[2]
  PIN um_k_zero[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 174.650 51.500 174.950 54.400 ;
    END
  END um_k_zero[3]
  PIN um_k_zero[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 345.310 0.000 345.610 3.580 ;
    END
  END um_k_zero[4]
  PIN um_k_zero[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 345.310 48.100 345.610 54.400 ;
    END
  END um_k_zero[5]
  PIN um_k_zero[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 515.970 0.000 516.270 2.220 ;
    END
  END um_k_zero[6]
  PIN um_k_zero[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 515.970 51.500 516.270 54.400 ;
    END
  END um_k_zero[7]
  PIN um_k_zero[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 686.630 0.000 686.930 6.980 ;
    END
  END um_k_zero[8]
  PIN um_k_zero[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 686.630 48.100 686.930 54.400 ;
    END
  END um_k_zero[9]
  PIN um_ow[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 0.000 92.610 2.900 ;
    END
  END um_ow[0]
  PIN um_ow[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 418.910 0.000 419.210 7.660 ;
    END
  END um_ow[100]
  PIN um_ow[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 415.230 0.000 415.530 7.660 ;
    END
  END um_ow[101]
  PIN um_ow[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 411.550 0.000 411.850 6.300 ;
    END
  END um_ow[102]
  PIN um_ow[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 407.870 0.000 408.170 7.660 ;
    END
  END um_ow[103]
  PIN um_ow[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 404.190 0.000 404.490 3.580 ;
    END
  END um_ow[104]
  PIN um_ow[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 400.510 0.000 400.810 7.660 ;
    END
  END um_ow[105]
  PIN um_ow[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 396.830 0.000 397.130 6.300 ;
    END
  END um_ow[106]
  PIN um_ow[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 393.150 0.000 393.450 3.580 ;
    END
  END um_ow[107]
  PIN um_ow[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 389.470 0.000 389.770 6.300 ;
    END
  END um_ow[108]
  PIN um_ow[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 385.790 0.000 386.090 4.940 ;
    END
  END um_ow[109]
  PIN um_ow[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 0.000 55.810 2.900 ;
    END
  END um_ow[10]
  PIN um_ow[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 382.110 0.000 382.410 6.300 ;
    END
  END um_ow[110]
  PIN um_ow[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 378.430 0.000 378.730 4.940 ;
    END
  END um_ow[111]
  PIN um_ow[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 374.750 0.000 375.050 2.900 ;
    END
  END um_ow[112]
  PIN um_ow[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 371.070 0.000 371.370 4.940 ;
    END
  END um_ow[113]
  PIN um_ow[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 367.390 0.000 367.690 6.300 ;
    END
  END um_ow[114]
  PIN um_ow[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 363.710 0.000 364.010 2.900 ;
    END
  END um_ow[115]
  PIN um_ow[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 360.030 0.000 360.330 4.940 ;
    END
  END um_ow[116]
  PIN um_ow[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 356.350 0.000 356.650 6.300 ;
    END
  END um_ow[117]
  PIN um_ow[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 352.670 0.000 352.970 4.940 ;
    END
  END um_ow[118]
  PIN um_ow[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 348.990 0.000 349.290 3.580 ;
    END
  END um_ow[119]
  PIN um_ow[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 0.000 52.130 2.900 ;
    END
  END um_ow[11]
  PIN um_ow[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 433.630 52.860 433.930 54.400 ;
    END
  END um_ow[120]
  PIN um_ow[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 429.950 49.460 430.250 54.400 ;
    END
  END um_ow[121]
  PIN um_ow[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 426.270 49.460 426.570 54.400 ;
    END
  END um_ow[122]
  PIN um_ow[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 422.590 52.860 422.890 54.400 ;
    END
  END um_ow[123]
  PIN um_ow[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 418.910 52.180 419.210 54.400 ;
    END
  END um_ow[124]
  PIN um_ow[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 415.230 48.100 415.530 54.400 ;
    END
  END um_ow[125]
  PIN um_ow[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 411.550 52.180 411.850 54.400 ;
    END
  END um_ow[126]
  PIN um_ow[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 407.870 48.780 408.170 54.400 ;
    END
  END um_ow[127]
  PIN um_ow[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 404.190 48.100 404.490 54.400 ;
    END
  END um_ow[128]
  PIN um_ow[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 400.510 45.380 400.810 54.400 ;
    END
  END um_ow[129]
  PIN um_ow[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 0.000 48.450 2.900 ;
    END
  END um_ow[12]
  PIN um_ow[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 396.830 48.780 397.130 54.400 ;
    END
  END um_ow[130]
  PIN um_ow[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 393.150 45.380 393.450 54.400 ;
    END
  END um_ow[131]
  PIN um_ow[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 389.470 48.100 389.770 54.400 ;
    END
  END um_ow[132]
  PIN um_ow[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 385.790 52.180 386.090 54.400 ;
    END
  END um_ow[133]
  PIN um_ow[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 382.110 48.780 382.410 54.400 ;
    END
  END um_ow[134]
  PIN um_ow[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 378.430 48.100 378.730 54.400 ;
    END
  END um_ow[135]
  PIN um_ow[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 374.750 45.380 375.050 54.400 ;
    END
  END um_ow[136]
  PIN um_ow[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 371.070 52.860 371.370 54.400 ;
    END
  END um_ow[137]
  PIN um_ow[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 367.390 45.380 367.690 54.400 ;
    END
  END um_ow[138]
  PIN um_ow[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 363.710 48.100 364.010 54.400 ;
    END
  END um_ow[139]
  PIN um_ow[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 0.000 44.770 3.580 ;
    END
  END um_ow[13]
  PIN um_ow[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 360.030 52.180 360.330 54.400 ;
    END
  END um_ow[140]
  PIN um_ow[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 356.350 52.860 356.650 54.400 ;
    END
  END um_ow[141]
  PIN um_ow[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 352.670 48.100 352.970 54.400 ;
    END
  END um_ow[142]
  PIN um_ow[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 348.990 45.380 349.290 54.400 ;
    END
  END um_ow[143]
  PIN um_ow[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 604.290 0.000 604.590 2.900 ;
    END
  END um_ow[144]
  PIN um_ow[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 600.610 0.000 600.910 2.900 ;
    END
  END um_ow[145]
  PIN um_ow[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 596.930 0.000 597.230 2.900 ;
    END
  END um_ow[146]
  PIN um_ow[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 593.250 0.000 593.550 2.900 ;
    END
  END um_ow[147]
  PIN um_ow[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 589.570 0.000 589.870 2.900 ;
    END
  END um_ow[148]
  PIN um_ow[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 585.890 0.000 586.190 1.850 ;
    END
  END um_ow[149]
  PIN um_ow[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 0.000 41.090 2.900 ;
    END
  END um_ow[14]
  PIN um_ow[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 582.210 0.000 582.510 2.900 ;
    END
  END um_ow[150]
  PIN um_ow[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 578.530 0.000 578.830 2.900 ;
    END
  END um_ow[151]
  PIN um_ow[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 574.850 0.000 575.150 2.900 ;
    END
  END um_ow[152]
  PIN um_ow[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 571.170 0.000 571.470 2.900 ;
    END
  END um_ow[153]
  PIN um_ow[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 567.490 0.000 567.790 1.540 ;
    END
  END um_ow[154]
  PIN um_ow[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 563.810 0.000 564.110 2.220 ;
    END
  END um_ow[155]
  PIN um_ow[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 560.130 0.000 560.430 2.220 ;
    END
  END um_ow[156]
  PIN um_ow[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 556.450 0.000 556.750 2.220 ;
    END
  END um_ow[157]
  PIN um_ow[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 552.770 0.000 553.070 2.220 ;
    END
  END um_ow[158]
  PIN um_ow[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 549.090 0.000 549.390 2.220 ;
    END
  END um_ow[159]
  PIN um_ow[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 0.000 37.410 3.580 ;
    END
  END um_ow[15]
  PIN um_ow[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 545.410 0.000 545.710 2.220 ;
    END
  END um_ow[160]
  PIN um_ow[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 541.730 0.000 542.030 2.220 ;
    END
  END um_ow[161]
  PIN um_ow[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 538.050 0.000 538.350 2.220 ;
    END
  END um_ow[162]
  PIN um_ow[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 534.370 0.000 534.670 2.220 ;
    END
  END um_ow[163]
  PIN um_ow[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 530.690 0.000 530.990 2.220 ;
    END
  END um_ow[164]
  PIN um_ow[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 527.010 0.000 527.310 2.220 ;
    END
  END um_ow[165]
  PIN um_ow[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 523.330 0.000 523.630 2.220 ;
    END
  END um_ow[166]
  PIN um_ow[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 519.650 0.000 519.950 2.220 ;
    END
  END um_ow[167]
  PIN um_ow[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 604.290 51.500 604.590 54.400 ;
    END
  END um_ow[168]
  PIN um_ow[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 600.610 51.500 600.910 54.400 ;
    END
  END um_ow[169]
  PIN um_ow[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 0.000 33.730 4.940 ;
    END
  END um_ow[16]
  PIN um_ow[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 596.930 51.500 597.230 54.400 ;
    END
  END um_ow[170]
  PIN um_ow[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 593.250 51.500 593.550 54.400 ;
    END
  END um_ow[171]
  PIN um_ow[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 589.570 51.500 589.870 54.400 ;
    END
  END um_ow[172]
  PIN um_ow[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 585.890 51.500 586.190 54.400 ;
    END
  END um_ow[173]
  PIN um_ow[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 582.210 51.500 582.510 54.400 ;
    END
  END um_ow[174]
  PIN um_ow[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 578.530 51.500 578.830 54.400 ;
    END
  END um_ow[175]
  PIN um_ow[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 574.850 51.500 575.150 54.400 ;
    END
  END um_ow[176]
  PIN um_ow[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 571.170 51.500 571.470 54.400 ;
    END
  END um_ow[177]
  PIN um_ow[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 567.490 51.500 567.790 54.400 ;
    END
  END um_ow[178]
  PIN um_ow[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 563.810 51.500 564.110 54.400 ;
    END
  END um_ow[179]
  PIN um_ow[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 0.000 30.050 3.580 ;
    END
  END um_ow[17]
  PIN um_ow[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 560.130 51.500 560.430 54.400 ;
    END
  END um_ow[180]
  PIN um_ow[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 556.450 51.500 556.750 54.400 ;
    END
  END um_ow[181]
  PIN um_ow[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 552.770 51.500 553.070 54.400 ;
    END
  END um_ow[182]
  PIN um_ow[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 549.090 51.500 549.390 54.400 ;
    END
  END um_ow[183]
  PIN um_ow[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 545.410 51.500 545.710 54.400 ;
    END
  END um_ow[184]
  PIN um_ow[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 541.730 51.500 542.030 54.400 ;
    END
  END um_ow[185]
  PIN um_ow[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 538.050 51.500 538.350 54.400 ;
    END
  END um_ow[186]
  PIN um_ow[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 534.370 51.500 534.670 54.400 ;
    END
  END um_ow[187]
  PIN um_ow[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 530.690 51.500 530.990 54.400 ;
    END
  END um_ow[188]
  PIN um_ow[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 527.010 51.500 527.310 54.400 ;
    END
  END um_ow[189]
  PIN um_ow[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 0.000 26.370 3.580 ;
    END
  END um_ow[18]
  PIN um_ow[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 523.330 51.500 523.630 54.400 ;
    END
  END um_ow[190]
  PIN um_ow[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 519.650 51.500 519.950 54.400 ;
    END
  END um_ow[191]
  PIN um_ow[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 774.950 0.000 775.250 6.300 ;
    END
  END um_ow[192]
  PIN um_ow[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 771.270 0.000 771.570 3.580 ;
    END
  END um_ow[193]
  PIN um_ow[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 767.590 0.000 767.890 2.900 ;
    END
  END um_ow[194]
  PIN um_ow[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 763.910 0.000 764.210 3.580 ;
    END
  END um_ow[195]
  PIN um_ow[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 760.230 0.000 760.530 3.580 ;
    END
  END um_ow[196]
  PIN um_ow[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 756.550 0.000 756.850 3.580 ;
    END
  END um_ow[197]
  PIN um_ow[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 752.870 0.000 753.170 3.580 ;
    END
  END um_ow[198]
  PIN um_ow[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 749.190 0.000 749.490 4.940 ;
    END
  END um_ow[199]
  PIN um_ow[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 0.000 22.690 4.940 ;
    END
  END um_ow[19]
  PIN um_ow[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 0.000 88.930 2.900 ;
    END
  END um_ow[1]
  PIN um_ow[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 745.510 0.000 745.810 3.580 ;
    END
  END um_ow[200]
  PIN um_ow[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 741.830 0.000 742.130 3.580 ;
    END
  END um_ow[201]
  PIN um_ow[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 738.150 0.000 738.450 2.900 ;
    END
  END um_ow[202]
  PIN um_ow[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 734.470 0.000 734.770 3.580 ;
    END
  END um_ow[203]
  PIN um_ow[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 730.790 0.000 731.090 3.580 ;
    END
  END um_ow[204]
  PIN um_ow[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 727.110 0.000 727.410 3.580 ;
    END
  END um_ow[205]
  PIN um_ow[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 723.430 0.000 723.730 6.980 ;
    END
  END um_ow[206]
  PIN um_ow[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 719.750 0.000 720.050 3.580 ;
    END
  END um_ow[207]
  PIN um_ow[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 716.070 0.000 716.370 3.580 ;
    END
  END um_ow[208]
  PIN um_ow[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 712.390 0.000 712.690 4.940 ;
    END
  END um_ow[209]
  PIN um_ow[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 0.000 19.010 2.900 ;
    END
  END um_ow[20]
  PIN um_ow[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 708.710 0.000 709.010 2.900 ;
    END
  END um_ow[210]
  PIN um_ow[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 705.030 0.000 705.330 3.580 ;
    END
  END um_ow[211]
  PIN um_ow[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 701.350 0.000 701.650 6.300 ;
    END
  END um_ow[212]
  PIN um_ow[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 697.670 0.000 697.970 2.220 ;
    END
  END um_ow[213]
  PIN um_ow[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 693.990 0.000 694.290 3.580 ;
    END
  END um_ow[214]
  PIN um_ow[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 690.310 0.000 690.610 2.900 ;
    END
  END um_ow[215]
  PIN um_ow[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 774.950 49.460 775.250 54.400 ;
    END
  END um_ow[216]
  PIN um_ow[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 771.270 50.820 771.570 54.400 ;
    END
  END um_ow[217]
  PIN um_ow[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 767.590 51.500 767.890 54.400 ;
    END
  END um_ow[218]
  PIN um_ow[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 763.910 50.820 764.210 54.400 ;
    END
  END um_ow[219]
  PIN um_ow[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 0.000 15.330 3.580 ;
    END
  END um_ow[21]
  PIN um_ow[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 760.230 50.820 760.530 54.400 ;
    END
  END um_ow[220]
  PIN um_ow[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 756.550 50.820 756.850 54.400 ;
    END
  END um_ow[221]
  PIN um_ow[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 752.870 50.820 753.170 54.400 ;
    END
  END um_ow[222]
  PIN um_ow[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 749.190 49.460 749.490 54.400 ;
    END
  END um_ow[223]
  PIN um_ow[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 745.510 50.820 745.810 54.400 ;
    END
  END um_ow[224]
  PIN um_ow[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 741.830 50.820 742.130 54.400 ;
    END
  END um_ow[225]
  PIN um_ow[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 738.150 52.180 738.450 54.400 ;
    END
  END um_ow[226]
  PIN um_ow[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 734.470 50.820 734.770 54.400 ;
    END
  END um_ow[227]
  PIN um_ow[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 730.790 50.820 731.090 54.400 ;
    END
  END um_ow[228]
  PIN um_ow[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 727.110 50.820 727.410 54.400 ;
    END
  END um_ow[229]
  PIN um_ow[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 0.000 11.650 4.940 ;
    END
  END um_ow[22]
  PIN um_ow[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 723.430 49.460 723.730 54.400 ;
    END
  END um_ow[230]
  PIN um_ow[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 719.750 50.820 720.050 54.400 ;
    END
  END um_ow[231]
  PIN um_ow[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 716.070 50.820 716.370 54.400 ;
    END
  END um_ow[232]
  PIN um_ow[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 712.390 51.500 712.690 54.400 ;
    END
  END um_ow[233]
  PIN um_ow[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 708.710 50.820 709.010 54.400 ;
    END
  END um_ow[234]
  PIN um_ow[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 705.030 50.820 705.330 54.400 ;
    END
  END um_ow[235]
  PIN um_ow[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 701.350 50.820 701.650 54.400 ;
    END
  END um_ow[236]
  PIN um_ow[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 697.670 49.460 697.970 54.400 ;
    END
  END um_ow[237]
  PIN um_ow[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 693.990 50.820 694.290 54.400 ;
    END
  END um_ow[238]
  PIN um_ow[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 690.310 51.500 690.610 54.400 ;
    END
  END um_ow[239]
  PIN um_ow[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 0.000 7.970 6.300 ;
    END
  END um_ow[23]
  PIN um_ow[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 945.610 0.000 945.910 1.850 ;
    END
  END um_ow[240]
  PIN um_ow[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 941.930 0.000 942.230 1.850 ;
    END
  END um_ow[241]
  PIN um_ow[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 938.250 0.000 938.550 1.850 ;
    END
  END um_ow[242]
  PIN um_ow[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 934.570 0.000 934.870 1.850 ;
    END
  END um_ow[243]
  PIN um_ow[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 930.890 0.000 931.190 1.850 ;
    END
  END um_ow[244]
  PIN um_ow[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 927.210 0.000 927.510 1.850 ;
    END
  END um_ow[245]
  PIN um_ow[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 923.530 0.000 923.830 1.850 ;
    END
  END um_ow[246]
  PIN um_ow[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 919.850 0.000 920.150 1.850 ;
    END
  END um_ow[247]
  PIN um_ow[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 916.170 0.000 916.470 1.850 ;
    END
  END um_ow[248]
  PIN um_ow[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 912.490 0.000 912.790 1.850 ;
    END
  END um_ow[249]
  PIN um_ow[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 50.820 92.610 54.400 ;
    END
  END um_ow[24]
  PIN um_ow[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 908.810 0.000 909.110 1.850 ;
    END
  END um_ow[250]
  PIN um_ow[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 905.130 0.000 905.430 1.850 ;
    END
  END um_ow[251]
  PIN um_ow[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 901.450 0.000 901.750 1.850 ;
    END
  END um_ow[252]
  PIN um_ow[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 897.770 0.000 898.070 1.850 ;
    END
  END um_ow[253]
  PIN um_ow[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 894.090 0.000 894.390 1.850 ;
    END
  END um_ow[254]
  PIN um_ow[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 890.410 0.000 890.710 1.850 ;
    END
  END um_ow[255]
  PIN um_ow[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 886.730 0.000 887.030 1.850 ;
    END
  END um_ow[256]
  PIN um_ow[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 883.050 0.000 883.350 1.850 ;
    END
  END um_ow[257]
  PIN um_ow[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 879.370 0.000 879.670 1.850 ;
    END
  END um_ow[258]
  PIN um_ow[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 875.690 0.000 875.990 1.850 ;
    END
  END um_ow[259]
  PIN um_ow[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 50.820 88.930 54.400 ;
    END
  END um_ow[25]
  PIN um_ow[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 872.010 0.000 872.310 1.850 ;
    END
  END um_ow[260]
  PIN um_ow[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 868.330 0.000 868.630 1.850 ;
    END
  END um_ow[261]
  PIN um_ow[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 864.650 0.000 864.950 1.850 ;
    END
  END um_ow[262]
  PIN um_ow[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 860.970 0.000 861.270 1.850 ;
    END
  END um_ow[263]
  PIN um_ow[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 945.610 51.500 945.910 54.400 ;
    END
  END um_ow[264]
  PIN um_ow[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 941.930 51.500 942.230 54.400 ;
    END
  END um_ow[265]
  PIN um_ow[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 938.250 51.500 938.550 54.400 ;
    END
  END um_ow[266]
  PIN um_ow[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 934.570 51.500 934.870 54.400 ;
    END
  END um_ow[267]
  PIN um_ow[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 930.890 51.500 931.190 54.400 ;
    END
  END um_ow[268]
  PIN um_ow[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 927.210 51.500 927.510 54.400 ;
    END
  END um_ow[269]
  PIN um_ow[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 50.820 85.250 54.400 ;
    END
  END um_ow[26]
  PIN um_ow[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 923.530 51.500 923.830 54.400 ;
    END
  END um_ow[270]
  PIN um_ow[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 919.850 51.500 920.150 54.400 ;
    END
  END um_ow[271]
  PIN um_ow[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 916.170 51.500 916.470 54.400 ;
    END
  END um_ow[272]
  PIN um_ow[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 912.490 51.500 912.790 54.400 ;
    END
  END um_ow[273]
  PIN um_ow[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 908.810 52.180 909.110 54.400 ;
    END
  END um_ow[274]
  PIN um_ow[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 905.130 51.500 905.430 54.400 ;
    END
  END um_ow[275]
  PIN um_ow[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 901.450 51.500 901.750 54.400 ;
    END
  END um_ow[276]
  PIN um_ow[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 897.770 51.500 898.070 54.400 ;
    END
  END um_ow[277]
  PIN um_ow[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 894.090 51.500 894.390 54.400 ;
    END
  END um_ow[278]
  PIN um_ow[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 890.410 51.500 890.710 54.400 ;
    END
  END um_ow[279]
  PIN um_ow[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 50.820 81.570 54.400 ;
    END
  END um_ow[27]
  PIN um_ow[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 886.730 51.500 887.030 54.400 ;
    END
  END um_ow[280]
  PIN um_ow[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 883.050 51.500 883.350 54.400 ;
    END
  END um_ow[281]
  PIN um_ow[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 879.370 51.500 879.670 54.400 ;
    END
  END um_ow[282]
  PIN um_ow[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 875.690 51.500 875.990 54.400 ;
    END
  END um_ow[283]
  PIN um_ow[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 872.010 51.500 872.310 54.400 ;
    END
  END um_ow[284]
  PIN um_ow[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 868.330 51.500 868.630 54.400 ;
    END
  END um_ow[285]
  PIN um_ow[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 864.650 51.500 864.950 54.400 ;
    END
  END um_ow[286]
  PIN um_ow[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 860.970 51.500 861.270 54.400 ;
    END
  END um_ow[287]
  PIN um_ow[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1116.270 0.000 1116.570 13.780 ;
    END
  END um_ow[288]
  PIN um_ow[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1112.590 0.000 1112.890 6.300 ;
    END
  END um_ow[289]
  PIN um_ow[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 50.820 77.890 54.400 ;
    END
  END um_ow[28]
  PIN um_ow[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1108.910 0.000 1109.210 1.540 ;
    END
  END um_ow[290]
  PIN um_ow[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1105.230 0.000 1105.530 4.260 ;
    END
  END um_ow[291]
  PIN um_ow[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1101.550 0.000 1101.850 6.980 ;
    END
  END um_ow[292]
  PIN um_ow[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1097.870 0.000 1098.170 1.540 ;
    END
  END um_ow[293]
  PIN um_ow[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1094.190 0.000 1094.490 1.540 ;
    END
  END um_ow[294]
  PIN um_ow[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1090.510 0.000 1090.810 4.260 ;
    END
  END um_ow[295]
  PIN um_ow[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1086.830 0.000 1087.130 4.260 ;
    END
  END um_ow[296]
  PIN um_ow[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1083.150 0.000 1083.450 6.980 ;
    END
  END um_ow[297]
  PIN um_ow[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1079.470 0.000 1079.770 4.260 ;
    END
  END um_ow[298]
  PIN um_ow[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1075.790 0.000 1076.090 4.260 ;
    END
  END um_ow[299]
  PIN um_ow[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 50.820 74.210 54.400 ;
    END
  END um_ow[29]
  PIN um_ow[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 0.000 85.250 2.900 ;
    END
  END um_ow[2]
  PIN um_ow[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1072.110 0.000 1072.410 4.260 ;
    END
  END um_ow[300]
  PIN um_ow[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1068.430 0.000 1068.730 4.260 ;
    END
  END um_ow[301]
  PIN um_ow[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1064.750 0.000 1065.050 4.260 ;
    END
  END um_ow[302]
  PIN um_ow[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1061.070 0.000 1061.370 4.260 ;
    END
  END um_ow[303]
  PIN um_ow[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1057.390 0.000 1057.690 4.940 ;
    END
  END um_ow[304]
  PIN um_ow[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1053.710 0.000 1054.010 6.300 ;
    END
  END um_ow[305]
  PIN um_ow[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1050.030 0.000 1050.330 4.940 ;
    END
  END um_ow[306]
  PIN um_ow[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1046.350 0.000 1046.650 4.260 ;
    END
  END um_ow[307]
  PIN um_ow[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1042.670 0.000 1042.970 4.260 ;
    END
  END um_ow[308]
  PIN um_ow[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1038.990 0.000 1039.290 4.260 ;
    END
  END um_ow[309]
  PIN um_ow[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 50.820 70.530 54.400 ;
    END
  END um_ow[30]
  PIN um_ow[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1035.310 0.000 1035.610 4.260 ;
    END
  END um_ow[310]
  PIN um_ow[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1031.630 0.000 1031.930 4.260 ;
    END
  END um_ow[311]
  PIN um_ow[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1116.270 50.820 1116.570 54.400 ;
    END
  END um_ow[312]
  PIN um_ow[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1112.590 51.500 1112.890 54.400 ;
    END
  END um_ow[313]
  PIN um_ow[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1108.910 51.500 1109.210 54.400 ;
    END
  END um_ow[314]
  PIN um_ow[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1105.230 52.180 1105.530 54.400 ;
    END
  END um_ow[315]
  PIN um_ow[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1101.550 51.500 1101.850 54.400 ;
    END
  END um_ow[316]
  PIN um_ow[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1097.870 50.820 1098.170 54.400 ;
    END
  END um_ow[317]
  PIN um_ow[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1094.190 50.820 1094.490 54.400 ;
    END
  END um_ow[318]
  PIN um_ow[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1090.510 52.860 1090.810 54.400 ;
    END
  END um_ow[319]
  PIN um_ow[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 49.460 66.850 54.400 ;
    END
  END um_ow[31]
  PIN um_ow[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1086.830 50.820 1087.130 54.400 ;
    END
  END um_ow[320]
  PIN um_ow[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1083.150 49.460 1083.450 54.400 ;
    END
  END um_ow[321]
  PIN um_ow[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1079.470 50.820 1079.770 54.400 ;
    END
  END um_ow[322]
  PIN um_ow[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1075.790 51.500 1076.090 54.400 ;
    END
  END um_ow[323]
  PIN um_ow[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1072.110 50.820 1072.410 54.400 ;
    END
  END um_ow[324]
  PIN um_ow[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1068.430 50.820 1068.730 54.400 ;
    END
  END um_ow[325]
  PIN um_ow[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1064.750 50.820 1065.050 54.400 ;
    END
  END um_ow[326]
  PIN um_ow[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1061.070 34.500 1061.370 54.400 ;
    END
  END um_ow[327]
  PIN um_ow[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1057.390 52.180 1057.690 54.400 ;
    END
  END um_ow[328]
  PIN um_ow[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1053.710 50.820 1054.010 54.400 ;
    END
  END um_ow[329]
  PIN um_ow[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 50.820 63.170 54.400 ;
    END
  END um_ow[32]
  PIN um_ow[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1050.030 52.180 1050.330 54.400 ;
    END
  END um_ow[330]
  PIN um_ow[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1046.350 50.820 1046.650 54.400 ;
    END
  END um_ow[331]
  PIN um_ow[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1042.670 50.820 1042.970 54.400 ;
    END
  END um_ow[332]
  PIN um_ow[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1038.990 52.860 1039.290 54.400 ;
    END
  END um_ow[333]
  PIN um_ow[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1035.310 50.820 1035.610 54.400 ;
    END
  END um_ow[334]
  PIN um_ow[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1031.630 50.820 1031.930 54.400 ;
    END
  END um_ow[335]
  PIN um_ow[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1286.930 0.000 1287.230 2.900 ;
    END
  END um_ow[336]
  PIN um_ow[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1283.250 0.000 1283.550 2.900 ;
    END
  END um_ow[337]
  PIN um_ow[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1279.570 0.000 1279.870 2.900 ;
    END
  END um_ow[338]
  PIN um_ow[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1275.890 0.000 1276.190 2.900 ;
    END
  END um_ow[339]
  PIN um_ow[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 50.820 59.490 54.400 ;
    END
  END um_ow[33]
  PIN um_ow[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1272.210 0.000 1272.510 1.540 ;
    END
  END um_ow[340]
  PIN um_ow[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1268.530 0.000 1268.830 2.900 ;
    END
  END um_ow[341]
  PIN um_ow[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1264.850 0.000 1265.150 2.900 ;
    END
  END um_ow[342]
  PIN um_ow[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1261.170 0.000 1261.470 2.900 ;
    END
  END um_ow[343]
  PIN um_ow[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1257.490 0.000 1257.790 2.900 ;
    END
  END um_ow[344]
  PIN um_ow[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1253.810 0.000 1254.110 1.850 ;
    END
  END um_ow[345]
  PIN um_ow[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1250.130 0.000 1250.430 2.900 ;
    END
  END um_ow[346]
  PIN um_ow[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1246.450 0.000 1246.750 1.850 ;
    END
  END um_ow[347]
  PIN um_ow[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1242.770 0.000 1243.070 2.220 ;
    END
  END um_ow[348]
  PIN um_ow[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1239.090 0.000 1239.390 1.850 ;
    END
  END um_ow[349]
  PIN um_ow[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 49.460 55.810 54.400 ;
    END
  END um_ow[34]
  PIN um_ow[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1235.410 0.000 1235.710 1.850 ;
    END
  END um_ow[350]
  PIN um_ow[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1231.730 0.000 1232.030 2.220 ;
    END
  END um_ow[351]
  PIN um_ow[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1228.050 0.000 1228.350 2.220 ;
    END
  END um_ow[352]
  PIN um_ow[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1224.370 0.000 1224.670 2.220 ;
    END
  END um_ow[353]
  PIN um_ow[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1220.690 0.000 1220.990 1.850 ;
    END
  END um_ow[354]
  PIN um_ow[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1217.010 0.000 1217.310 2.220 ;
    END
  END um_ow[355]
  PIN um_ow[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1213.330 0.000 1213.630 1.850 ;
    END
  END um_ow[356]
  PIN um_ow[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1209.650 0.000 1209.950 2.220 ;
    END
  END um_ow[357]
  PIN um_ow[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1205.970 0.000 1206.270 2.220 ;
    END
  END um_ow[358]
  PIN um_ow[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1202.290 0.000 1202.590 1.540 ;
    END
  END um_ow[359]
  PIN um_ow[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 49.460 52.130 54.400 ;
    END
  END um_ow[35]
  PIN um_ow[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1286.930 51.500 1287.230 54.400 ;
    END
  END um_ow[360]
  PIN um_ow[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1283.250 51.500 1283.550 54.400 ;
    END
  END um_ow[361]
  PIN um_ow[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1279.570 51.500 1279.870 54.400 ;
    END
  END um_ow[362]
  PIN um_ow[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1275.890 51.500 1276.190 54.400 ;
    END
  END um_ow[363]
  PIN um_ow[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1272.210 51.500 1272.510 54.400 ;
    END
  END um_ow[364]
  PIN um_ow[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1268.530 51.500 1268.830 54.400 ;
    END
  END um_ow[365]
  PIN um_ow[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1264.850 51.500 1265.150 54.400 ;
    END
  END um_ow[366]
  PIN um_ow[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1261.170 51.500 1261.470 54.400 ;
    END
  END um_ow[367]
  PIN um_ow[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1257.490 51.500 1257.790 54.400 ;
    END
  END um_ow[368]
  PIN um_ow[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1253.810 51.500 1254.110 54.400 ;
    END
  END um_ow[369]
  PIN um_ow[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 52.860 48.450 54.400 ;
    END
  END um_ow[36]
  PIN um_ow[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1250.130 51.500 1250.430 54.400 ;
    END
  END um_ow[370]
  PIN um_ow[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1246.450 51.500 1246.750 54.400 ;
    END
  END um_ow[371]
  PIN um_ow[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1242.770 51.500 1243.070 54.400 ;
    END
  END um_ow[372]
  PIN um_ow[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1239.090 51.500 1239.390 54.400 ;
    END
  END um_ow[373]
  PIN um_ow[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1235.410 51.500 1235.710 54.400 ;
    END
  END um_ow[374]
  PIN um_ow[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1231.730 51.500 1232.030 54.400 ;
    END
  END um_ow[375]
  PIN um_ow[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1228.050 51.500 1228.350 54.400 ;
    END
  END um_ow[376]
  PIN um_ow[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1224.370 51.500 1224.670 54.400 ;
    END
  END um_ow[377]
  PIN um_ow[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1220.690 51.500 1220.990 54.400 ;
    END
  END um_ow[378]
  PIN um_ow[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1217.010 51.500 1217.310 54.400 ;
    END
  END um_ow[379]
  PIN um_ow[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 50.820 44.770 54.400 ;
    END
  END um_ow[37]
  PIN um_ow[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1213.330 51.500 1213.630 54.400 ;
    END
  END um_ow[380]
  PIN um_ow[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1209.650 51.500 1209.950 54.400 ;
    END
  END um_ow[381]
  PIN um_ow[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1205.970 51.500 1206.270 54.400 ;
    END
  END um_ow[382]
  PIN um_ow[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1202.290 51.500 1202.590 54.400 ;
    END
  END um_ow[383]
  PIN um_ow[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 49.460 41.090 54.400 ;
    END
  END um_ow[38]
  PIN um_ow[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 50.820 37.410 54.400 ;
    END
  END um_ow[39]
  PIN um_ow[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 0.000 81.570 6.980 ;
    END
  END um_ow[3]
  PIN um_ow[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 50.820 33.730 54.400 ;
    END
  END um_ow[40]
  PIN um_ow[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 50.820 30.050 54.400 ;
    END
  END um_ow[41]
  PIN um_ow[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 50.820 26.370 54.400 ;
    END
  END um_ow[42]
  PIN um_ow[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 50.820 22.690 54.400 ;
    END
  END um_ow[43]
  PIN um_ow[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 50.820 19.010 54.400 ;
    END
  END um_ow[44]
  PIN um_ow[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 49.460 15.330 54.400 ;
    END
  END um_ow[45]
  PIN um_ow[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 50.820 11.650 54.400 ;
    END
  END um_ow[46]
  PIN um_ow[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 50.820 7.970 54.400 ;
    END
  END um_ow[47]
  PIN um_ow[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 262.970 0.000 263.270 2.900 ;
    END
  END um_ow[48]
  PIN um_ow[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 259.290 0.000 259.590 2.900 ;
    END
  END um_ow[49]
  PIN um_ow[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 0.000 77.890 3.580 ;
    END
  END um_ow[4]
  PIN um_ow[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 255.610 0.000 255.910 2.900 ;
    END
  END um_ow[50]
  PIN um_ow[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 251.930 0.000 252.230 2.900 ;
    END
  END um_ow[51]
  PIN um_ow[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 248.250 0.000 248.550 2.900 ;
    END
  END um_ow[52]
  PIN um_ow[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 244.570 0.000 244.870 2.900 ;
    END
  END um_ow[53]
  PIN um_ow[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 240.890 0.000 241.190 2.900 ;
    END
  END um_ow[54]
  PIN um_ow[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 237.210 0.000 237.510 2.900 ;
    END
  END um_ow[55]
  PIN um_ow[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 233.530 0.000 233.830 2.900 ;
    END
  END um_ow[56]
  PIN um_ow[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 229.850 0.000 230.150 2.900 ;
    END
  END um_ow[57]
  PIN um_ow[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 226.170 0.000 226.470 2.900 ;
    END
  END um_ow[58]
  PIN um_ow[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 222.490 0.000 222.790 2.900 ;
    END
  END um_ow[59]
  PIN um_ow[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 0.000 74.210 3.580 ;
    END
  END um_ow[5]
  PIN um_ow[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 218.810 0.000 219.110 2.900 ;
    END
  END um_ow[60]
  PIN um_ow[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 215.130 0.000 215.430 2.900 ;
    END
  END um_ow[61]
  PIN um_ow[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 211.450 0.000 211.750 2.900 ;
    END
  END um_ow[62]
  PIN um_ow[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 207.770 0.000 208.070 2.900 ;
    END
  END um_ow[63]
  PIN um_ow[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 204.090 0.000 204.390 2.900 ;
    END
  END um_ow[64]
  PIN um_ow[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 200.410 0.000 200.710 2.900 ;
    END
  END um_ow[65]
  PIN um_ow[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 196.730 0.000 197.030 1.540 ;
    END
  END um_ow[66]
  PIN um_ow[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 193.050 0.000 193.350 2.900 ;
    END
  END um_ow[67]
  PIN um_ow[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 189.370 0.000 189.670 2.900 ;
    END
  END um_ow[68]
  PIN um_ow[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 185.690 0.000 185.990 2.900 ;
    END
  END um_ow[69]
  PIN um_ow[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 0.000 70.530 4.940 ;
    END
  END um_ow[6]
  PIN um_ow[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 182.010 0.000 182.310 2.900 ;
    END
  END um_ow[70]
  PIN um_ow[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 178.330 0.000 178.630 2.900 ;
    END
  END um_ow[71]
  PIN um_ow[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 262.970 51.500 263.270 54.400 ;
    END
  END um_ow[72]
  PIN um_ow[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 259.290 51.500 259.590 54.400 ;
    END
  END um_ow[73]
  PIN um_ow[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 255.610 51.500 255.910 54.400 ;
    END
  END um_ow[74]
  PIN um_ow[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 251.930 51.500 252.230 54.400 ;
    END
  END um_ow[75]
  PIN um_ow[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 248.250 51.500 248.550 54.400 ;
    END
  END um_ow[76]
  PIN um_ow[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 244.570 51.500 244.870 54.400 ;
    END
  END um_ow[77]
  PIN um_ow[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 240.890 51.500 241.190 54.400 ;
    END
  END um_ow[78]
  PIN um_ow[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 237.210 51.500 237.510 54.400 ;
    END
  END um_ow[79]
  PIN um_ow[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 0.000 66.850 2.900 ;
    END
  END um_ow[7]
  PIN um_ow[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 233.530 51.500 233.830 54.400 ;
    END
  END um_ow[80]
  PIN um_ow[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 229.850 51.500 230.150 54.400 ;
    END
  END um_ow[81]
  PIN um_ow[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 226.170 51.500 226.470 54.400 ;
    END
  END um_ow[82]
  PIN um_ow[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 222.490 51.500 222.790 54.400 ;
    END
  END um_ow[83]
  PIN um_ow[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 218.810 51.500 219.110 54.400 ;
    END
  END um_ow[84]
  PIN um_ow[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 215.130 51.500 215.430 54.400 ;
    END
  END um_ow[85]
  PIN um_ow[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 211.450 51.500 211.750 54.400 ;
    END
  END um_ow[86]
  PIN um_ow[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 207.770 51.500 208.070 54.400 ;
    END
  END um_ow[87]
  PIN um_ow[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 204.090 51.500 204.390 54.400 ;
    END
  END um_ow[88]
  PIN um_ow[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 200.410 51.500 200.710 54.400 ;
    END
  END um_ow[89]
  PIN um_ow[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 0.000 63.170 2.900 ;
    END
  END um_ow[8]
  PIN um_ow[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 196.730 51.500 197.030 54.400 ;
    END
  END um_ow[90]
  PIN um_ow[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 193.050 51.500 193.350 54.400 ;
    END
  END um_ow[91]
  PIN um_ow[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 189.370 51.500 189.670 54.400 ;
    END
  END um_ow[92]
  PIN um_ow[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 185.690 51.500 185.990 54.400 ;
    END
  END um_ow[93]
  PIN um_ow[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 182.010 51.500 182.310 54.400 ;
    END
  END um_ow[94]
  PIN um_ow[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 178.330 51.500 178.630 54.400 ;
    END
  END um_ow[95]
  PIN um_ow[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 433.630 0.000 433.930 3.580 ;
    END
  END um_ow[96]
  PIN um_ow[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 429.950 0.000 430.250 4.940 ;
    END
  END um_ow[97]
  PIN um_ow[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 426.270 0.000 426.570 3.580 ;
    END
  END um_ow[98]
  PIN um_ow[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 422.590 0.000 422.890 3.580 ;
    END
  END um_ow[99]
  PIN um_ow[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 0.000 59.490 2.900 ;
    END
  END um_ow[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 173.710 5.200 175.310 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 511.695 5.200 513.295 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 849.680 5.200 851.280 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1187.665 5.200 1189.265 49.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 342.700 5.200 344.300 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 680.685 5.200 682.285 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1018.670 5.200 1020.270 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1356.655 5.200 1358.255 49.200 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 1357.460 49.045 ;
      LAYER met1 ;
        RECT 4.210 1.060 1361.070 54.360 ;
      LAYER met2 ;
        RECT 4.230 0.155 1361.050 54.390 ;
      LAYER met3 ;
        RECT 3.750 48.490 1362.210 54.225 ;
        RECT 3.750 47.810 1360.590 48.490 ;
        RECT 3.750 47.130 1359.670 47.810 ;
        RECT 3.750 46.450 1344.550 47.130 ;
        RECT 3.750 45.350 1339.950 46.450 ;
        RECT 3.750 44.670 1340.410 45.350 ;
        RECT 3.750 44.410 1359.730 44.670 ;
        RECT 3.750 43.310 1358.750 44.410 ;
        RECT 3.750 43.050 1361.120 43.310 ;
        RECT 3.750 41.950 1352.830 43.050 ;
        RECT 3.750 41.690 1356.050 41.950 ;
        RECT 3.750 41.010 1352.370 41.690 ;
        RECT 3.750 40.330 1351.450 41.010 ;
        RECT 3.750 39.650 1350.530 40.330 ;
        RECT 3.750 38.550 1339.950 39.650 ;
        RECT 3.750 37.610 1358.810 38.550 ;
        RECT 3.750 36.510 1339.950 37.610 ;
        RECT 3.750 36.250 1359.730 36.510 ;
        RECT 3.750 35.150 1312.350 36.250 ;
        RECT 3.750 34.470 1339.950 35.150 ;
        RECT 3.750 33.790 1340.410 34.470 ;
        RECT 3.750 33.530 1360.190 33.790 ;
        RECT 3.750 32.850 1359.270 33.530 ;
        RECT 3.750 31.750 1358.750 32.850 ;
        RECT 3.750 31.490 1359.730 31.750 ;
        RECT 3.750 30.390 1344.550 31.490 ;
        RECT 3.750 30.130 1358.810 30.390 ;
        RECT 3.750 29.450 1358.350 30.130 ;
        RECT 3.750 28.770 1356.910 29.450 ;
        RECT 3.750 27.670 1355.990 28.770 ;
        RECT 3.750 26.990 1358.810 27.670 ;
        RECT 3.750 26.730 1359.730 26.990 ;
        RECT 3.750 25.630 1344.550 26.730 ;
        RECT 3.750 25.370 1359.730 25.630 ;
        RECT 3.750 24.270 1340.410 25.370 ;
        RECT 3.750 23.590 1344.090 24.270 ;
        RECT 3.750 22.910 1360.650 23.590 ;
        RECT 3.750 22.650 1361.120 22.910 ;
        RECT 3.750 21.970 1359.440 22.650 ;
        RECT 3.750 21.290 1358.750 21.970 ;
        RECT 3.750 20.190 1220.810 21.290 ;
        RECT 3.750 19.510 1355.990 20.190 ;
        RECT 3.750 18.830 1356.910 19.510 ;
        RECT 3.750 18.570 1357.890 18.830 ;
        RECT 3.750 17.470 1339.490 18.570 ;
        RECT 3.750 17.210 1359.730 17.470 ;
        RECT 3.750 16.110 1358.750 17.210 ;
        RECT 3.750 15.850 1358.810 16.110 ;
        RECT 3.750 14.750 1310.970 15.850 ;
        RECT 3.750 14.490 1359.730 14.750 ;
        RECT 3.750 13.810 1353.750 14.490 ;
        RECT 3.750 12.710 1335.810 13.810 ;
        RECT 3.750 12.030 1342.250 12.710 ;
        RECT 3.750 11.770 1359.730 12.030 ;
        RECT 3.750 10.670 1358.750 11.770 ;
        RECT 3.750 9.990 1358.810 10.670 ;
        RECT 3.750 9.730 1360.650 9.990 ;
        RECT 3.750 9.050 1350.470 9.730 ;
        RECT 3.750 8.370 1349.550 9.050 ;
        RECT 3.750 7.690 1345.010 8.370 ;
        RECT 3.750 7.010 1344.090 7.690 ;
        RECT 3.750 5.910 1344.030 7.010 ;
        RECT 3.750 5.650 1358.810 5.910 ;
        RECT 3.750 4.550 1358.750 5.650 ;
        RECT 3.750 0.175 1362.210 4.550 ;
      LAYER met4 ;
        RECT 4.690 50.420 7.270 52.865 ;
        RECT 8.370 50.420 10.950 52.865 ;
        RECT 12.050 50.420 14.630 52.865 ;
        RECT 4.690 49.060 14.630 50.420 ;
        RECT 15.730 50.420 18.310 52.865 ;
        RECT 19.410 50.420 21.990 52.865 ;
        RECT 23.090 50.420 25.670 52.865 ;
        RECT 26.770 50.420 29.350 52.865 ;
        RECT 30.450 50.420 33.030 52.865 ;
        RECT 34.130 50.420 36.710 52.865 ;
        RECT 37.810 50.420 40.390 52.865 ;
        RECT 15.730 49.060 40.390 50.420 ;
        RECT 41.490 50.420 44.070 52.865 ;
        RECT 45.170 52.460 47.750 52.865 ;
        RECT 48.850 52.460 51.430 52.865 ;
        RECT 45.170 50.420 51.430 52.460 ;
        RECT 41.490 49.060 51.430 50.420 ;
        RECT 52.530 49.060 55.110 52.865 ;
        RECT 56.210 50.420 58.790 52.865 ;
        RECT 59.890 50.420 62.470 52.865 ;
        RECT 63.570 50.420 66.150 52.865 ;
        RECT 56.210 49.060 66.150 50.420 ;
        RECT 67.250 50.420 69.830 52.865 ;
        RECT 70.930 50.420 73.510 52.865 ;
        RECT 74.610 50.420 77.190 52.865 ;
        RECT 78.290 50.420 80.870 52.865 ;
        RECT 81.970 50.420 84.550 52.865 ;
        RECT 85.650 50.420 88.230 52.865 ;
        RECT 89.330 50.420 91.910 52.865 ;
        RECT 93.010 50.420 95.590 52.865 ;
        RECT 67.250 49.060 95.590 50.420 ;
        RECT 4.690 45.660 95.590 49.060 ;
        RECT 3.975 34.100 95.590 45.660 ;
        RECT 96.690 34.100 99.270 52.865 ;
        RECT 100.370 52.460 102.950 52.865 ;
        RECT 104.050 52.460 106.630 52.865 ;
        RECT 100.370 49.060 106.630 52.460 ;
        RECT 107.730 50.420 110.310 52.865 ;
        RECT 111.410 50.420 113.990 52.865 ;
        RECT 107.730 49.060 113.990 50.420 ;
        RECT 100.370 34.100 113.990 49.060 ;
        RECT 115.090 34.100 117.670 52.865 ;
        RECT 118.770 42.940 121.350 52.865 ;
        RECT 122.450 42.940 125.030 52.865 ;
        RECT 118.770 34.100 125.030 42.940 ;
        RECT 126.130 47.700 128.710 52.865 ;
        RECT 129.810 47.700 132.390 52.865 ;
        RECT 126.130 41.580 132.390 47.700 ;
        RECT 133.490 41.580 136.070 52.865 ;
        RECT 126.130 38.860 136.070 41.580 ;
        RECT 137.170 41.580 139.750 52.865 ;
        RECT 140.850 47.020 143.430 52.865 ;
        RECT 144.530 47.020 147.110 52.865 ;
        RECT 140.850 42.940 147.110 47.020 ;
        RECT 148.210 42.940 150.790 52.865 ;
        RECT 151.890 42.940 154.470 52.865 ;
        RECT 155.570 51.100 158.150 52.865 ;
        RECT 159.250 51.100 161.830 52.865 ;
        RECT 155.570 47.700 161.830 51.100 ;
        RECT 162.930 51.100 174.250 52.865 ;
        RECT 175.350 51.100 177.930 52.865 ;
        RECT 179.030 51.100 181.610 52.865 ;
        RECT 182.710 51.100 185.290 52.865 ;
        RECT 186.390 51.100 188.970 52.865 ;
        RECT 190.070 51.100 192.650 52.865 ;
        RECT 193.750 51.100 196.330 52.865 ;
        RECT 197.430 51.100 200.010 52.865 ;
        RECT 201.110 51.100 203.690 52.865 ;
        RECT 204.790 51.100 207.370 52.865 ;
        RECT 208.470 51.100 211.050 52.865 ;
        RECT 212.150 51.100 214.730 52.865 ;
        RECT 215.830 51.100 218.410 52.865 ;
        RECT 219.510 51.100 222.090 52.865 ;
        RECT 223.190 51.100 225.770 52.865 ;
        RECT 226.870 51.100 229.450 52.865 ;
        RECT 230.550 51.100 233.130 52.865 ;
        RECT 234.230 51.100 236.810 52.865 ;
        RECT 237.910 51.100 240.490 52.865 ;
        RECT 241.590 51.100 244.170 52.865 ;
        RECT 245.270 51.100 247.850 52.865 ;
        RECT 248.950 51.100 251.530 52.865 ;
        RECT 252.630 51.100 255.210 52.865 ;
        RECT 256.310 51.100 258.890 52.865 ;
        RECT 259.990 51.100 262.570 52.865 ;
        RECT 263.670 51.100 266.250 52.865 ;
        RECT 267.350 51.780 269.930 52.865 ;
        RECT 271.030 51.780 273.610 52.865 ;
        RECT 267.350 51.100 273.610 51.780 ;
        RECT 274.710 51.100 277.290 52.865 ;
        RECT 278.390 51.100 280.970 52.865 ;
        RECT 282.070 51.100 284.650 52.865 ;
        RECT 285.750 51.100 288.330 52.865 ;
        RECT 289.430 51.100 292.010 52.865 ;
        RECT 293.110 51.100 295.690 52.865 ;
        RECT 296.790 51.100 299.370 52.865 ;
        RECT 300.470 51.100 303.050 52.865 ;
        RECT 304.150 51.100 306.730 52.865 ;
        RECT 307.830 51.100 310.410 52.865 ;
        RECT 311.510 51.100 314.090 52.865 ;
        RECT 315.190 51.100 317.770 52.865 ;
        RECT 318.870 51.100 321.450 52.865 ;
        RECT 322.550 51.100 325.130 52.865 ;
        RECT 326.230 51.100 328.810 52.865 ;
        RECT 329.910 51.100 332.490 52.865 ;
        RECT 333.590 51.100 344.910 52.865 ;
        RECT 162.930 49.600 344.910 51.100 ;
        RECT 162.930 47.700 173.310 49.600 ;
        RECT 155.570 42.940 173.310 47.700 ;
        RECT 140.850 41.580 173.310 42.940 ;
        RECT 137.170 38.860 173.310 41.580 ;
        RECT 126.130 34.100 173.310 38.860 ;
        RECT 3.975 16.900 173.310 34.100 ;
        RECT 3.975 14.860 121.350 16.900 ;
        RECT 3.975 7.380 95.590 14.860 ;
        RECT 4.690 6.700 80.870 7.380 ;
        RECT 4.690 1.535 7.270 6.700 ;
        RECT 8.370 5.340 80.870 6.700 ;
        RECT 8.370 1.535 10.950 5.340 ;
        RECT 12.050 3.980 21.990 5.340 ;
        RECT 12.050 1.535 14.630 3.980 ;
        RECT 15.730 3.300 21.990 3.980 ;
        RECT 15.730 1.535 18.310 3.300 ;
        RECT 19.410 1.535 21.990 3.300 ;
        RECT 23.090 3.980 33.030 5.340 ;
        RECT 23.090 1.535 25.670 3.980 ;
        RECT 26.770 1.535 29.350 3.980 ;
        RECT 30.450 1.535 33.030 3.980 ;
        RECT 34.130 3.980 69.830 5.340 ;
        RECT 34.130 1.535 36.710 3.980 ;
        RECT 37.810 3.300 44.070 3.980 ;
        RECT 37.810 1.535 40.390 3.300 ;
        RECT 41.490 1.535 44.070 3.300 ;
        RECT 45.170 3.300 69.830 3.980 ;
        RECT 45.170 1.535 47.750 3.300 ;
        RECT 48.850 1.535 51.430 3.300 ;
        RECT 52.530 1.535 55.110 3.300 ;
        RECT 56.210 1.535 58.790 3.300 ;
        RECT 59.890 1.535 62.470 3.300 ;
        RECT 63.570 1.535 66.150 3.300 ;
        RECT 67.250 1.535 69.830 3.300 ;
        RECT 70.930 3.980 80.870 5.340 ;
        RECT 70.930 1.535 73.510 3.980 ;
        RECT 74.610 1.535 77.190 3.980 ;
        RECT 78.290 1.535 80.870 3.980 ;
        RECT 81.970 3.300 95.590 7.380 ;
        RECT 81.970 1.535 84.550 3.300 ;
        RECT 85.650 1.535 88.230 3.300 ;
        RECT 89.330 1.535 91.910 3.300 ;
        RECT 93.010 1.535 95.590 3.300 ;
        RECT 96.690 14.180 113.990 14.860 ;
        RECT 96.690 1.535 99.270 14.180 ;
        RECT 100.370 8.740 110.310 14.180 ;
        RECT 100.370 7.380 106.630 8.740 ;
        RECT 100.370 1.535 102.950 7.380 ;
        RECT 104.050 1.535 106.630 7.380 ;
        RECT 107.730 1.535 110.310 8.740 ;
        RECT 111.410 1.535 113.990 14.180 ;
        RECT 115.090 3.300 121.350 14.860 ;
        RECT 115.090 1.535 117.670 3.300 ;
        RECT 118.770 1.535 121.350 3.300 ;
        RECT 122.450 14.180 173.310 16.900 ;
        RECT 122.450 1.535 125.030 14.180 ;
        RECT 126.130 7.380 173.310 14.180 ;
        RECT 126.130 6.700 161.830 7.380 ;
        RECT 126.130 1.535 128.710 6.700 ;
        RECT 129.810 1.535 132.390 6.700 ;
        RECT 133.490 1.535 136.070 6.700 ;
        RECT 137.170 3.300 161.830 6.700 ;
        RECT 137.170 2.620 143.430 3.300 ;
        RECT 137.170 1.535 139.750 2.620 ;
        RECT 140.850 1.535 143.430 2.620 ;
        RECT 144.530 2.620 150.790 3.300 ;
        RECT 144.530 1.535 147.110 2.620 ;
        RECT 148.210 1.535 150.790 2.620 ;
        RECT 151.890 2.620 161.830 3.300 ;
        RECT 151.890 1.940 158.150 2.620 ;
        RECT 151.890 1.535 154.470 1.940 ;
        RECT 155.570 1.535 158.150 1.940 ;
        RECT 159.250 1.535 161.830 2.620 ;
        RECT 162.930 4.800 173.310 7.380 ;
        RECT 175.710 4.800 342.300 49.600 ;
        RECT 344.700 47.700 344.910 49.600 ;
        RECT 346.010 47.700 348.590 52.865 ;
        RECT 344.700 44.980 348.590 47.700 ;
        RECT 349.690 47.700 352.270 52.865 ;
        RECT 353.370 52.460 355.950 52.865 ;
        RECT 357.050 52.460 359.630 52.865 ;
        RECT 353.370 51.780 359.630 52.460 ;
        RECT 360.730 51.780 363.310 52.865 ;
        RECT 353.370 47.700 363.310 51.780 ;
        RECT 364.410 47.700 366.990 52.865 ;
        RECT 349.690 44.980 366.990 47.700 ;
        RECT 368.090 52.460 370.670 52.865 ;
        RECT 371.770 52.460 374.350 52.865 ;
        RECT 368.090 44.980 374.350 52.460 ;
        RECT 375.450 47.700 378.030 52.865 ;
        RECT 379.130 48.380 381.710 52.865 ;
        RECT 382.810 51.780 385.390 52.865 ;
        RECT 386.490 51.780 389.070 52.865 ;
        RECT 382.810 48.380 389.070 51.780 ;
        RECT 379.130 47.700 389.070 48.380 ;
        RECT 390.170 47.700 392.750 52.865 ;
        RECT 375.450 44.980 392.750 47.700 ;
        RECT 393.850 48.380 396.430 52.865 ;
        RECT 397.530 48.380 400.110 52.865 ;
        RECT 393.850 44.980 400.110 48.380 ;
        RECT 401.210 47.700 403.790 52.865 ;
        RECT 404.890 48.380 407.470 52.865 ;
        RECT 408.570 51.780 411.150 52.865 ;
        RECT 412.250 51.780 414.830 52.865 ;
        RECT 408.570 48.380 414.830 51.780 ;
        RECT 404.890 47.700 414.830 48.380 ;
        RECT 415.930 51.780 418.510 52.865 ;
        RECT 419.610 52.460 422.190 52.865 ;
        RECT 423.290 52.460 425.870 52.865 ;
        RECT 419.610 51.780 425.870 52.460 ;
        RECT 415.930 49.060 425.870 51.780 ;
        RECT 426.970 49.060 429.550 52.865 ;
        RECT 430.650 52.460 433.230 52.865 ;
        RECT 434.330 52.460 436.910 52.865 ;
        RECT 430.650 49.060 436.910 52.460 ;
        RECT 415.930 47.700 436.910 49.060 ;
        RECT 401.210 44.980 436.910 47.700 ;
        RECT 344.700 42.940 436.910 44.980 ;
        RECT 438.010 45.660 440.590 52.865 ;
        RECT 441.690 45.660 444.270 52.865 ;
        RECT 438.010 42.940 444.270 45.660 ;
        RECT 344.700 40.220 444.270 42.940 ;
        RECT 445.370 51.100 447.950 52.865 ;
        RECT 449.050 51.100 451.630 52.865 ;
        RECT 445.370 42.940 451.630 51.100 ;
        RECT 452.730 43.620 455.310 52.865 ;
        RECT 456.410 43.620 458.990 52.865 ;
        RECT 452.730 42.940 458.990 43.620 ;
        RECT 460.090 42.940 462.670 52.865 ;
        RECT 445.370 41.580 462.670 42.940 ;
        RECT 463.770 48.380 466.350 52.865 ;
        RECT 467.450 48.380 470.030 52.865 ;
        RECT 463.770 42.940 470.030 48.380 ;
        RECT 471.130 42.940 473.710 52.865 ;
        RECT 474.810 48.380 477.390 52.865 ;
        RECT 478.490 48.380 481.070 52.865 ;
        RECT 482.170 48.380 484.750 52.865 ;
        RECT 474.810 42.940 484.750 48.380 ;
        RECT 485.850 48.380 488.430 52.865 ;
        RECT 489.530 48.380 492.110 52.865 ;
        RECT 485.850 42.940 492.110 48.380 ;
        RECT 493.210 42.940 495.790 52.865 ;
        RECT 463.770 41.580 495.790 42.940 ;
        RECT 445.370 40.900 495.790 41.580 ;
        RECT 496.890 42.940 499.470 52.865 ;
        RECT 500.570 48.380 503.150 52.865 ;
        RECT 504.250 51.100 515.570 52.865 ;
        RECT 516.670 51.100 519.250 52.865 ;
        RECT 520.350 51.100 522.930 52.865 ;
        RECT 524.030 51.100 526.610 52.865 ;
        RECT 527.710 51.100 530.290 52.865 ;
        RECT 531.390 51.100 533.970 52.865 ;
        RECT 535.070 51.100 537.650 52.865 ;
        RECT 538.750 51.100 541.330 52.865 ;
        RECT 542.430 51.100 545.010 52.865 ;
        RECT 546.110 51.100 548.690 52.865 ;
        RECT 549.790 51.100 552.370 52.865 ;
        RECT 553.470 51.100 556.050 52.865 ;
        RECT 557.150 51.100 559.730 52.865 ;
        RECT 560.830 51.100 563.410 52.865 ;
        RECT 564.510 51.100 567.090 52.865 ;
        RECT 568.190 51.100 570.770 52.865 ;
        RECT 571.870 51.100 574.450 52.865 ;
        RECT 575.550 51.100 578.130 52.865 ;
        RECT 579.230 51.100 581.810 52.865 ;
        RECT 582.910 51.100 585.490 52.865 ;
        RECT 586.590 51.100 589.170 52.865 ;
        RECT 590.270 51.100 592.850 52.865 ;
        RECT 593.950 51.100 596.530 52.865 ;
        RECT 597.630 51.100 600.210 52.865 ;
        RECT 601.310 51.100 603.890 52.865 ;
        RECT 604.990 51.100 607.570 52.865 ;
        RECT 608.670 51.100 611.250 52.865 ;
        RECT 612.350 51.100 614.930 52.865 ;
        RECT 616.030 51.100 618.610 52.865 ;
        RECT 619.710 51.100 622.290 52.865 ;
        RECT 623.390 51.780 625.970 52.865 ;
        RECT 627.070 51.780 629.650 52.865 ;
        RECT 623.390 51.100 629.650 51.780 ;
        RECT 630.750 51.100 633.330 52.865 ;
        RECT 634.430 51.100 637.010 52.865 ;
        RECT 638.110 51.780 640.690 52.865 ;
        RECT 641.790 51.780 644.370 52.865 ;
        RECT 638.110 51.100 644.370 51.780 ;
        RECT 645.470 51.100 648.050 52.865 ;
        RECT 649.150 51.100 651.730 52.865 ;
        RECT 652.830 51.100 655.410 52.865 ;
        RECT 656.510 51.100 659.090 52.865 ;
        RECT 660.190 51.100 662.770 52.865 ;
        RECT 663.870 51.100 666.450 52.865 ;
        RECT 667.550 51.100 670.130 52.865 ;
        RECT 671.230 51.100 673.810 52.865 ;
        RECT 674.910 51.100 686.230 52.865 ;
        RECT 504.250 49.600 686.230 51.100 ;
        RECT 504.250 48.380 511.295 49.600 ;
        RECT 500.570 42.940 511.295 48.380 ;
        RECT 496.890 40.900 511.295 42.940 ;
        RECT 445.370 40.220 511.295 40.900 ;
        RECT 344.700 8.060 511.295 40.220 ;
        RECT 344.700 6.700 400.110 8.060 ;
        RECT 344.700 5.340 355.950 6.700 ;
        RECT 344.700 4.800 352.270 5.340 ;
        RECT 162.930 3.980 352.270 4.800 ;
        RECT 162.930 3.300 344.910 3.980 ;
        RECT 162.930 1.940 177.930 3.300 ;
        RECT 162.930 1.535 174.250 1.940 ;
        RECT 175.350 1.535 177.930 1.940 ;
        RECT 179.030 1.535 181.610 3.300 ;
        RECT 182.710 1.535 185.290 3.300 ;
        RECT 186.390 1.535 188.970 3.300 ;
        RECT 190.070 1.535 192.650 3.300 ;
        RECT 193.750 1.940 200.010 3.300 ;
        RECT 193.750 1.535 196.330 1.940 ;
        RECT 197.430 1.535 200.010 1.940 ;
        RECT 201.110 1.535 203.690 3.300 ;
        RECT 204.790 1.535 207.370 3.300 ;
        RECT 208.470 1.535 211.050 3.300 ;
        RECT 212.150 1.535 214.730 3.300 ;
        RECT 215.830 1.535 218.410 3.300 ;
        RECT 219.510 1.535 222.090 3.300 ;
        RECT 223.190 1.535 225.770 3.300 ;
        RECT 226.870 1.535 229.450 3.300 ;
        RECT 230.550 1.535 233.130 3.300 ;
        RECT 234.230 1.535 236.810 3.300 ;
        RECT 237.910 1.535 240.490 3.300 ;
        RECT 241.590 1.535 244.170 3.300 ;
        RECT 245.270 1.535 247.850 3.300 ;
        RECT 248.950 1.535 251.530 3.300 ;
        RECT 252.630 1.535 255.210 3.300 ;
        RECT 256.310 1.535 258.890 3.300 ;
        RECT 259.990 1.535 262.570 3.300 ;
        RECT 263.670 1.535 266.250 3.300 ;
        RECT 267.350 2.250 273.610 3.300 ;
        RECT 267.350 1.535 269.930 2.250 ;
        RECT 271.030 1.535 273.610 2.250 ;
        RECT 274.710 1.535 277.290 3.300 ;
        RECT 278.390 1.535 280.970 3.300 ;
        RECT 282.070 1.535 284.650 3.300 ;
        RECT 285.750 1.535 288.330 3.300 ;
        RECT 289.430 1.535 292.010 3.300 ;
        RECT 293.110 2.250 303.050 3.300 ;
        RECT 293.110 1.535 295.690 2.250 ;
        RECT 296.790 1.535 299.370 2.250 ;
        RECT 300.470 1.535 303.050 2.250 ;
        RECT 304.150 1.535 306.730 3.300 ;
        RECT 307.830 1.535 310.410 3.300 ;
        RECT 311.510 1.535 314.090 3.300 ;
        RECT 315.190 1.535 317.770 3.300 ;
        RECT 318.870 1.535 321.450 3.300 ;
        RECT 322.550 1.535 325.130 3.300 ;
        RECT 326.230 2.620 344.910 3.300 ;
        RECT 326.230 1.535 328.810 2.620 ;
        RECT 329.910 1.535 332.490 2.620 ;
        RECT 333.590 1.535 344.910 2.620 ;
        RECT 346.010 1.535 348.590 3.980 ;
        RECT 349.690 1.535 352.270 3.980 ;
        RECT 353.370 1.535 355.950 5.340 ;
        RECT 357.050 5.340 366.990 6.700 ;
        RECT 357.050 1.535 359.630 5.340 ;
        RECT 360.730 3.300 366.990 5.340 ;
        RECT 360.730 1.535 363.310 3.300 ;
        RECT 364.410 1.535 366.990 3.300 ;
        RECT 368.090 5.340 381.710 6.700 ;
        RECT 368.090 1.535 370.670 5.340 ;
        RECT 371.770 3.300 378.030 5.340 ;
        RECT 371.770 1.535 374.350 3.300 ;
        RECT 375.450 1.535 378.030 3.300 ;
        RECT 379.130 1.535 381.710 5.340 ;
        RECT 382.810 5.340 389.070 6.700 ;
        RECT 382.810 1.535 385.390 5.340 ;
        RECT 386.490 1.535 389.070 5.340 ;
        RECT 390.170 3.980 396.430 6.700 ;
        RECT 390.170 1.535 392.750 3.980 ;
        RECT 393.850 1.535 396.430 3.980 ;
        RECT 397.530 1.535 400.110 6.700 ;
        RECT 401.210 3.980 407.470 8.060 ;
        RECT 401.210 1.535 403.790 3.980 ;
        RECT 404.890 1.535 407.470 3.980 ;
        RECT 408.570 6.700 414.830 8.060 ;
        RECT 408.570 1.535 411.150 6.700 ;
        RECT 412.250 1.535 414.830 6.700 ;
        RECT 415.930 1.535 418.510 8.060 ;
        RECT 419.610 6.700 495.790 8.060 ;
        RECT 419.610 5.340 436.910 6.700 ;
        RECT 419.610 3.980 429.550 5.340 ;
        RECT 419.610 1.535 422.190 3.980 ;
        RECT 423.290 1.535 425.870 3.980 ;
        RECT 426.970 1.535 429.550 3.980 ;
        RECT 430.650 3.980 436.910 5.340 ;
        RECT 430.650 1.535 433.230 3.980 ;
        RECT 434.330 1.535 436.910 3.980 ;
        RECT 438.010 6.020 444.270 6.700 ;
        RECT 438.010 1.535 440.590 6.020 ;
        RECT 441.690 1.535 444.270 6.020 ;
        RECT 445.370 6.020 495.790 6.700 ;
        RECT 445.370 3.980 470.030 6.020 ;
        RECT 445.370 1.940 451.630 3.980 ;
        RECT 445.370 1.535 447.950 1.940 ;
        RECT 449.050 1.535 451.630 1.940 ;
        RECT 452.730 1.940 458.990 3.980 ;
        RECT 452.730 1.535 455.310 1.940 ;
        RECT 456.410 1.535 458.990 1.940 ;
        RECT 460.090 1.940 466.350 3.980 ;
        RECT 460.090 1.535 462.670 1.940 ;
        RECT 463.770 1.535 466.350 1.940 ;
        RECT 467.450 1.535 470.030 3.980 ;
        RECT 471.130 1.535 473.710 6.020 ;
        RECT 474.810 1.535 477.390 6.020 ;
        RECT 478.490 1.535 481.070 6.020 ;
        RECT 482.170 3.980 495.790 6.020 ;
        RECT 482.170 2.620 488.430 3.980 ;
        RECT 482.170 1.535 484.750 2.620 ;
        RECT 485.850 1.535 488.430 2.620 ;
        RECT 489.530 1.535 492.110 3.980 ;
        RECT 493.210 1.535 495.790 3.980 ;
        RECT 496.890 4.800 511.295 8.060 ;
        RECT 513.695 4.800 680.285 49.600 ;
        RECT 682.685 47.700 686.230 49.600 ;
        RECT 687.330 51.100 689.910 52.865 ;
        RECT 691.010 51.100 693.590 52.865 ;
        RECT 687.330 50.420 693.590 51.100 ;
        RECT 694.690 50.420 697.270 52.865 ;
        RECT 687.330 49.060 697.270 50.420 ;
        RECT 698.370 50.420 700.950 52.865 ;
        RECT 702.050 50.420 704.630 52.865 ;
        RECT 705.730 50.420 708.310 52.865 ;
        RECT 709.410 51.100 711.990 52.865 ;
        RECT 713.090 51.100 715.670 52.865 ;
        RECT 709.410 50.420 715.670 51.100 ;
        RECT 716.770 50.420 719.350 52.865 ;
        RECT 720.450 50.420 723.030 52.865 ;
        RECT 698.370 49.060 723.030 50.420 ;
        RECT 724.130 50.420 726.710 52.865 ;
        RECT 727.810 50.420 730.390 52.865 ;
        RECT 731.490 50.420 734.070 52.865 ;
        RECT 735.170 51.780 737.750 52.865 ;
        RECT 738.850 51.780 741.430 52.865 ;
        RECT 735.170 50.420 741.430 51.780 ;
        RECT 742.530 50.420 745.110 52.865 ;
        RECT 746.210 50.420 748.790 52.865 ;
        RECT 724.130 49.060 748.790 50.420 ;
        RECT 749.890 50.420 752.470 52.865 ;
        RECT 753.570 50.420 756.150 52.865 ;
        RECT 757.250 50.420 759.830 52.865 ;
        RECT 760.930 50.420 763.510 52.865 ;
        RECT 764.610 51.100 767.190 52.865 ;
        RECT 768.290 51.100 770.870 52.865 ;
        RECT 764.610 50.420 770.870 51.100 ;
        RECT 771.970 50.420 774.550 52.865 ;
        RECT 749.890 49.060 774.550 50.420 ;
        RECT 775.650 49.060 778.230 52.865 ;
        RECT 687.330 48.380 778.230 49.060 ;
        RECT 779.330 48.380 781.910 52.865 ;
        RECT 783.010 51.100 785.590 52.865 ;
        RECT 786.690 51.100 789.270 52.865 ;
        RECT 783.010 48.380 789.270 51.100 ;
        RECT 790.370 48.380 792.950 52.865 ;
        RECT 687.330 47.700 792.950 48.380 ;
        RECT 682.685 47.020 792.950 47.700 ;
        RECT 794.050 48.380 796.630 52.865 ;
        RECT 797.730 48.380 800.310 52.865 ;
        RECT 794.050 47.020 800.310 48.380 ;
        RECT 682.685 41.580 800.310 47.020 ;
        RECT 801.410 41.580 803.990 52.865 ;
        RECT 805.090 42.260 807.670 52.865 ;
        RECT 808.770 42.260 811.350 52.865 ;
        RECT 805.090 41.580 811.350 42.260 ;
        RECT 812.450 41.580 815.030 52.865 ;
        RECT 816.130 48.380 818.710 52.865 ;
        RECT 819.810 48.380 822.390 52.865 ;
        RECT 816.130 41.580 822.390 48.380 ;
        RECT 823.490 41.580 826.070 52.865 ;
        RECT 827.170 41.580 829.750 52.865 ;
        RECT 830.850 41.580 833.430 52.865 ;
        RECT 682.685 40.900 833.430 41.580 ;
        RECT 834.530 41.580 837.110 52.865 ;
        RECT 838.210 41.580 840.790 52.865 ;
        RECT 834.530 40.900 840.790 41.580 ;
        RECT 682.685 40.220 840.790 40.900 ;
        RECT 841.890 45.660 844.470 52.865 ;
        RECT 845.570 51.100 856.890 52.865 ;
        RECT 857.990 51.100 860.570 52.865 ;
        RECT 861.670 51.100 864.250 52.865 ;
        RECT 865.350 51.100 867.930 52.865 ;
        RECT 869.030 51.100 871.610 52.865 ;
        RECT 872.710 51.100 875.290 52.865 ;
        RECT 876.390 51.100 878.970 52.865 ;
        RECT 880.070 51.100 882.650 52.865 ;
        RECT 883.750 51.100 886.330 52.865 ;
        RECT 887.430 51.100 890.010 52.865 ;
        RECT 891.110 51.100 893.690 52.865 ;
        RECT 894.790 51.100 897.370 52.865 ;
        RECT 898.470 51.100 901.050 52.865 ;
        RECT 902.150 51.100 904.730 52.865 ;
        RECT 905.830 51.780 908.410 52.865 ;
        RECT 909.510 51.780 912.090 52.865 ;
        RECT 905.830 51.100 912.090 51.780 ;
        RECT 913.190 51.100 915.770 52.865 ;
        RECT 916.870 51.100 919.450 52.865 ;
        RECT 920.550 51.100 923.130 52.865 ;
        RECT 924.230 51.100 926.810 52.865 ;
        RECT 927.910 51.100 930.490 52.865 ;
        RECT 931.590 51.100 934.170 52.865 ;
        RECT 935.270 51.100 937.850 52.865 ;
        RECT 938.950 51.100 941.530 52.865 ;
        RECT 942.630 51.100 945.210 52.865 ;
        RECT 946.310 51.100 948.890 52.865 ;
        RECT 949.990 51.780 952.570 52.865 ;
        RECT 953.670 51.780 956.250 52.865 ;
        RECT 949.990 51.100 956.250 51.780 ;
        RECT 957.350 51.100 959.930 52.865 ;
        RECT 961.030 51.100 963.610 52.865 ;
        RECT 964.710 51.780 967.290 52.865 ;
        RECT 968.390 51.780 970.970 52.865 ;
        RECT 964.710 51.100 970.970 51.780 ;
        RECT 972.070 51.100 974.650 52.865 ;
        RECT 975.750 51.100 978.330 52.865 ;
        RECT 979.430 51.100 982.010 52.865 ;
        RECT 983.110 51.100 985.690 52.865 ;
        RECT 986.790 51.100 989.370 52.865 ;
        RECT 990.470 51.780 993.050 52.865 ;
        RECT 994.150 51.780 996.730 52.865 ;
        RECT 990.470 51.100 996.730 51.780 ;
        RECT 997.830 51.100 1000.410 52.865 ;
        RECT 1001.510 51.780 1004.090 52.865 ;
        RECT 1005.190 51.780 1007.770 52.865 ;
        RECT 1001.510 51.100 1007.770 51.780 ;
        RECT 1008.870 51.780 1011.450 52.865 ;
        RECT 1012.550 51.780 1015.130 52.865 ;
        RECT 1008.870 51.100 1015.130 51.780 ;
        RECT 1016.230 51.100 1027.550 52.865 ;
        RECT 845.570 49.600 1027.550 51.100 ;
        RECT 845.570 45.660 849.280 49.600 ;
        RECT 841.890 40.220 849.280 45.660 ;
        RECT 682.685 14.180 849.280 40.220 ;
        RECT 682.685 7.380 785.590 14.180 ;
        RECT 682.685 4.800 686.230 7.380 ;
        RECT 496.890 4.660 686.230 4.800 ;
        RECT 496.890 2.620 503.150 4.660 ;
        RECT 496.890 1.535 499.470 2.620 ;
        RECT 500.570 1.535 503.150 2.620 ;
        RECT 504.250 3.300 686.230 4.660 ;
        RECT 504.250 2.620 570.770 3.300 ;
        RECT 504.250 1.535 515.570 2.620 ;
        RECT 516.670 1.535 519.250 2.620 ;
        RECT 520.350 1.535 522.930 2.620 ;
        RECT 524.030 1.535 526.610 2.620 ;
        RECT 527.710 1.535 530.290 2.620 ;
        RECT 531.390 1.535 533.970 2.620 ;
        RECT 535.070 1.535 537.650 2.620 ;
        RECT 538.750 1.535 541.330 2.620 ;
        RECT 542.430 1.535 545.010 2.620 ;
        RECT 546.110 1.535 548.690 2.620 ;
        RECT 549.790 1.535 552.370 2.620 ;
        RECT 553.470 1.535 556.050 2.620 ;
        RECT 557.150 1.535 559.730 2.620 ;
        RECT 560.830 1.535 563.410 2.620 ;
        RECT 564.510 1.940 570.770 2.620 ;
        RECT 564.510 1.535 567.090 1.940 ;
        RECT 568.190 1.535 570.770 1.940 ;
        RECT 571.870 1.535 574.450 3.300 ;
        RECT 575.550 1.535 578.130 3.300 ;
        RECT 579.230 1.535 581.810 3.300 ;
        RECT 582.910 2.250 589.170 3.300 ;
        RECT 582.910 1.535 585.490 2.250 ;
        RECT 586.590 1.535 589.170 2.250 ;
        RECT 590.270 1.535 592.850 3.300 ;
        RECT 593.950 1.535 596.530 3.300 ;
        RECT 597.630 1.535 600.210 3.300 ;
        RECT 601.310 1.535 603.890 3.300 ;
        RECT 604.990 1.535 607.570 3.300 ;
        RECT 608.670 1.535 611.250 3.300 ;
        RECT 612.350 1.535 614.930 3.300 ;
        RECT 616.030 1.535 618.610 3.300 ;
        RECT 619.710 1.535 622.290 3.300 ;
        RECT 623.390 1.535 625.970 3.300 ;
        RECT 627.070 1.535 629.650 3.300 ;
        RECT 630.750 1.535 633.330 3.300 ;
        RECT 634.430 1.535 637.010 3.300 ;
        RECT 638.110 2.250 644.370 3.300 ;
        RECT 638.110 1.535 640.690 2.250 ;
        RECT 641.790 1.535 644.370 2.250 ;
        RECT 645.470 1.535 648.050 3.300 ;
        RECT 649.150 1.940 655.410 3.300 ;
        RECT 649.150 1.535 651.730 1.940 ;
        RECT 652.830 1.535 655.410 1.940 ;
        RECT 656.510 1.535 659.090 3.300 ;
        RECT 660.190 1.535 662.770 3.300 ;
        RECT 663.870 1.535 666.450 3.300 ;
        RECT 667.550 1.535 670.130 3.300 ;
        RECT 671.230 2.250 686.230 3.300 ;
        RECT 671.230 1.535 673.810 2.250 ;
        RECT 674.910 1.535 686.230 2.250 ;
        RECT 687.330 6.700 723.030 7.380 ;
        RECT 687.330 3.980 700.950 6.700 ;
        RECT 687.330 3.300 693.590 3.980 ;
        RECT 687.330 1.535 689.910 3.300 ;
        RECT 691.010 1.535 693.590 3.300 ;
        RECT 694.690 2.620 700.950 3.980 ;
        RECT 694.690 1.535 697.270 2.620 ;
        RECT 698.370 1.535 700.950 2.620 ;
        RECT 702.050 5.340 723.030 6.700 ;
        RECT 702.050 3.980 711.990 5.340 ;
        RECT 702.050 1.535 704.630 3.980 ;
        RECT 705.730 3.300 711.990 3.980 ;
        RECT 705.730 1.535 708.310 3.300 ;
        RECT 709.410 1.535 711.990 3.300 ;
        RECT 713.090 3.980 723.030 5.340 ;
        RECT 713.090 1.535 715.670 3.980 ;
        RECT 716.770 1.535 719.350 3.980 ;
        RECT 720.450 1.535 723.030 3.980 ;
        RECT 724.130 6.700 778.230 7.380 ;
        RECT 724.130 5.340 774.550 6.700 ;
        RECT 724.130 3.980 748.790 5.340 ;
        RECT 724.130 1.535 726.710 3.980 ;
        RECT 727.810 1.535 730.390 3.980 ;
        RECT 731.490 1.535 734.070 3.980 ;
        RECT 735.170 3.300 741.430 3.980 ;
        RECT 735.170 1.535 737.750 3.300 ;
        RECT 738.850 1.535 741.430 3.300 ;
        RECT 742.530 1.535 745.110 3.980 ;
        RECT 746.210 1.535 748.790 3.980 ;
        RECT 749.890 3.980 774.550 5.340 ;
        RECT 749.890 1.535 752.470 3.980 ;
        RECT 753.570 1.535 756.150 3.980 ;
        RECT 757.250 1.535 759.830 3.980 ;
        RECT 760.930 1.535 763.510 3.980 ;
        RECT 764.610 3.300 770.870 3.980 ;
        RECT 764.610 1.535 767.190 3.300 ;
        RECT 768.290 1.535 770.870 3.300 ;
        RECT 771.970 1.535 774.550 3.980 ;
        RECT 775.650 1.535 778.230 6.700 ;
        RECT 779.330 1.535 781.910 7.380 ;
        RECT 783.010 1.535 785.590 7.380 ;
        RECT 786.690 7.380 796.630 14.180 ;
        RECT 786.690 1.535 789.270 7.380 ;
        RECT 790.370 3.300 796.630 7.380 ;
        RECT 790.370 1.535 792.950 3.300 ;
        RECT 794.050 1.535 796.630 3.300 ;
        RECT 797.730 7.380 849.280 14.180 ;
        RECT 797.730 6.020 818.710 7.380 ;
        RECT 797.730 1.535 800.310 6.020 ;
        RECT 801.410 3.300 807.670 6.020 ;
        RECT 801.410 1.535 803.990 3.300 ;
        RECT 805.090 1.535 807.670 3.300 ;
        RECT 808.770 3.300 815.030 6.020 ;
        RECT 808.770 1.535 811.350 3.300 ;
        RECT 812.450 1.535 815.030 3.300 ;
        RECT 816.130 1.535 818.710 6.020 ;
        RECT 819.810 6.020 840.790 7.380 ;
        RECT 819.810 3.300 826.070 6.020 ;
        RECT 819.810 1.535 822.390 3.300 ;
        RECT 823.490 1.535 826.070 3.300 ;
        RECT 827.170 1.535 829.750 6.020 ;
        RECT 830.850 1.535 833.430 6.020 ;
        RECT 834.530 3.300 840.790 6.020 ;
        RECT 834.530 1.535 837.110 3.300 ;
        RECT 838.210 1.535 840.790 3.300 ;
        RECT 841.890 4.800 849.280 7.380 ;
        RECT 851.680 4.800 1018.270 49.600 ;
        RECT 1020.670 47.700 1027.550 49.600 ;
        RECT 1028.650 50.420 1031.230 52.865 ;
        RECT 1032.330 50.420 1034.910 52.865 ;
        RECT 1036.010 52.460 1038.590 52.865 ;
        RECT 1039.690 52.460 1042.270 52.865 ;
        RECT 1036.010 50.420 1042.270 52.460 ;
        RECT 1043.370 50.420 1045.950 52.865 ;
        RECT 1047.050 51.780 1049.630 52.865 ;
        RECT 1050.730 51.780 1053.310 52.865 ;
        RECT 1047.050 50.420 1053.310 51.780 ;
        RECT 1054.410 51.780 1056.990 52.865 ;
        RECT 1058.090 51.780 1060.670 52.865 ;
        RECT 1054.410 50.420 1060.670 51.780 ;
        RECT 1028.650 47.700 1060.670 50.420 ;
        RECT 1020.670 34.100 1060.670 47.700 ;
        RECT 1061.770 50.420 1064.350 52.865 ;
        RECT 1065.450 50.420 1068.030 52.865 ;
        RECT 1069.130 50.420 1071.710 52.865 ;
        RECT 1072.810 51.100 1075.390 52.865 ;
        RECT 1076.490 51.100 1079.070 52.865 ;
        RECT 1072.810 50.420 1079.070 51.100 ;
        RECT 1080.170 50.420 1082.750 52.865 ;
        RECT 1061.770 49.060 1082.750 50.420 ;
        RECT 1083.850 50.420 1086.430 52.865 ;
        RECT 1087.530 52.460 1090.110 52.865 ;
        RECT 1091.210 52.460 1093.790 52.865 ;
        RECT 1087.530 50.420 1093.790 52.460 ;
        RECT 1094.890 50.420 1097.470 52.865 ;
        RECT 1098.570 51.100 1101.150 52.865 ;
        RECT 1102.250 51.780 1104.830 52.865 ;
        RECT 1105.930 51.780 1108.510 52.865 ;
        RECT 1102.250 51.100 1108.510 51.780 ;
        RECT 1109.610 51.100 1112.190 52.865 ;
        RECT 1113.290 51.100 1115.870 52.865 ;
        RECT 1098.570 50.420 1115.870 51.100 ;
        RECT 1116.970 50.420 1119.550 52.865 ;
        RECT 1083.850 49.060 1119.550 50.420 ;
        RECT 1061.770 45.660 1119.550 49.060 ;
        RECT 1120.650 45.660 1123.230 52.865 ;
        RECT 1061.770 41.580 1123.230 45.660 ;
        RECT 1124.330 48.380 1126.910 52.865 ;
        RECT 1128.010 48.380 1130.590 52.865 ;
        RECT 1124.330 42.940 1130.590 48.380 ;
        RECT 1131.690 42.940 1134.270 52.865 ;
        RECT 1135.370 42.940 1137.950 52.865 ;
        RECT 1139.050 47.020 1141.630 52.865 ;
        RECT 1142.730 47.020 1145.310 52.865 ;
        RECT 1139.050 42.940 1145.310 47.020 ;
        RECT 1146.410 48.380 1148.990 52.865 ;
        RECT 1150.090 48.380 1152.670 52.865 ;
        RECT 1146.410 42.940 1152.670 48.380 ;
        RECT 1124.330 41.580 1152.670 42.940 ;
        RECT 1153.770 48.380 1156.350 52.865 ;
        RECT 1157.450 48.380 1160.030 52.865 ;
        RECT 1153.770 42.940 1160.030 48.380 ;
        RECT 1161.130 42.940 1163.710 52.865 ;
        RECT 1164.810 48.380 1167.390 52.865 ;
        RECT 1168.490 48.380 1171.070 52.865 ;
        RECT 1172.170 48.380 1174.750 52.865 ;
        RECT 1175.850 48.380 1178.430 52.865 ;
        RECT 1164.810 45.660 1178.430 48.380 ;
        RECT 1179.530 45.660 1182.110 52.865 ;
        RECT 1164.810 42.940 1182.110 45.660 ;
        RECT 1183.210 45.660 1185.790 52.865 ;
        RECT 1186.890 51.100 1198.210 52.865 ;
        RECT 1199.310 51.100 1201.890 52.865 ;
        RECT 1202.990 51.100 1205.570 52.865 ;
        RECT 1206.670 51.100 1209.250 52.865 ;
        RECT 1210.350 51.100 1212.930 52.865 ;
        RECT 1214.030 51.100 1216.610 52.865 ;
        RECT 1217.710 51.100 1220.290 52.865 ;
        RECT 1221.390 51.100 1223.970 52.865 ;
        RECT 1225.070 51.100 1227.650 52.865 ;
        RECT 1228.750 51.100 1231.330 52.865 ;
        RECT 1232.430 51.100 1235.010 52.865 ;
        RECT 1236.110 51.100 1238.690 52.865 ;
        RECT 1239.790 51.100 1242.370 52.865 ;
        RECT 1243.470 51.100 1246.050 52.865 ;
        RECT 1247.150 51.100 1249.730 52.865 ;
        RECT 1250.830 51.100 1253.410 52.865 ;
        RECT 1254.510 51.100 1257.090 52.865 ;
        RECT 1258.190 51.100 1260.770 52.865 ;
        RECT 1261.870 51.100 1264.450 52.865 ;
        RECT 1265.550 51.100 1268.130 52.865 ;
        RECT 1269.230 51.100 1271.810 52.865 ;
        RECT 1272.910 51.100 1275.490 52.865 ;
        RECT 1276.590 51.100 1279.170 52.865 ;
        RECT 1280.270 51.100 1282.850 52.865 ;
        RECT 1283.950 51.100 1286.530 52.865 ;
        RECT 1287.630 51.100 1290.210 52.865 ;
        RECT 1291.310 51.100 1293.890 52.865 ;
        RECT 1294.990 51.100 1297.570 52.865 ;
        RECT 1298.670 51.100 1301.250 52.865 ;
        RECT 1302.350 51.780 1304.930 52.865 ;
        RECT 1306.030 51.780 1308.610 52.865 ;
        RECT 1302.350 51.100 1308.610 51.780 ;
        RECT 1309.710 51.100 1312.290 52.865 ;
        RECT 1313.390 51.100 1315.970 52.865 ;
        RECT 1317.070 51.100 1319.650 52.865 ;
        RECT 1320.750 51.780 1323.330 52.865 ;
        RECT 1324.430 51.780 1327.010 52.865 ;
        RECT 1320.750 51.100 1327.010 51.780 ;
        RECT 1328.110 52.150 1330.690 52.865 ;
        RECT 1331.790 52.150 1334.370 52.865 ;
        RECT 1328.110 51.100 1334.370 52.150 ;
        RECT 1186.890 50.790 1334.370 51.100 ;
        RECT 1335.470 50.790 1338.050 52.865 ;
        RECT 1339.150 50.790 1341.730 52.865 ;
        RECT 1342.830 50.790 1345.410 52.865 ;
        RECT 1346.510 50.790 1349.090 52.865 ;
        RECT 1350.190 50.790 1352.770 52.865 ;
        RECT 1353.870 50.790 1356.450 52.865 ;
        RECT 1186.890 49.600 1357.165 50.790 ;
        RECT 1186.890 45.660 1187.265 49.600 ;
        RECT 1183.210 42.940 1187.265 45.660 ;
        RECT 1153.770 41.580 1187.265 42.940 ;
        RECT 1061.770 34.100 1187.265 41.580 ;
        RECT 1020.670 14.180 1187.265 34.100 ;
        RECT 1020.670 7.380 1115.870 14.180 ;
        RECT 1020.670 6.700 1082.750 7.380 ;
        RECT 1020.670 5.340 1053.310 6.700 ;
        RECT 1020.670 4.800 1049.630 5.340 ;
        RECT 841.890 4.660 1049.630 4.800 ;
        RECT 841.890 3.300 1031.230 4.660 ;
        RECT 841.890 1.535 844.470 3.300 ;
        RECT 845.570 2.250 1031.230 3.300 ;
        RECT 845.570 1.535 856.890 2.250 ;
        RECT 857.990 1.535 860.570 2.250 ;
        RECT 861.670 1.535 864.250 2.250 ;
        RECT 865.350 1.535 867.930 2.250 ;
        RECT 869.030 1.535 871.610 2.250 ;
        RECT 872.710 1.535 875.290 2.250 ;
        RECT 876.390 1.535 878.970 2.250 ;
        RECT 880.070 1.535 882.650 2.250 ;
        RECT 883.750 1.535 886.330 2.250 ;
        RECT 887.430 1.535 890.010 2.250 ;
        RECT 891.110 1.535 893.690 2.250 ;
        RECT 894.790 1.535 897.370 2.250 ;
        RECT 898.470 1.535 901.050 2.250 ;
        RECT 902.150 1.535 904.730 2.250 ;
        RECT 905.830 1.535 908.410 2.250 ;
        RECT 909.510 1.535 912.090 2.250 ;
        RECT 913.190 1.535 915.770 2.250 ;
        RECT 916.870 1.535 919.450 2.250 ;
        RECT 920.550 1.535 923.130 2.250 ;
        RECT 924.230 1.535 926.810 2.250 ;
        RECT 927.910 1.535 930.490 2.250 ;
        RECT 931.590 1.535 934.170 2.250 ;
        RECT 935.270 1.535 937.850 2.250 ;
        RECT 938.950 1.535 941.530 2.250 ;
        RECT 942.630 1.535 945.210 2.250 ;
        RECT 946.310 1.535 948.890 2.250 ;
        RECT 949.990 1.535 952.570 2.250 ;
        RECT 953.670 1.535 956.250 2.250 ;
        RECT 957.350 1.535 959.930 2.250 ;
        RECT 961.030 1.535 963.610 2.250 ;
        RECT 964.710 1.535 967.290 2.250 ;
        RECT 968.390 1.535 970.970 2.250 ;
        RECT 972.070 1.535 974.650 2.250 ;
        RECT 975.750 1.535 978.330 2.250 ;
        RECT 979.430 1.535 982.010 2.250 ;
        RECT 983.110 1.535 985.690 2.250 ;
        RECT 986.790 1.535 989.370 2.250 ;
        RECT 990.470 1.535 993.050 2.250 ;
        RECT 994.150 1.535 996.730 2.250 ;
        RECT 997.830 1.535 1000.410 2.250 ;
        RECT 1001.510 1.535 1004.090 2.250 ;
        RECT 1005.190 1.535 1007.770 2.250 ;
        RECT 1008.870 1.535 1011.450 2.250 ;
        RECT 1012.550 1.535 1015.130 2.250 ;
        RECT 1016.230 1.535 1027.550 2.250 ;
        RECT 1028.650 1.535 1031.230 2.250 ;
        RECT 1032.330 1.535 1034.910 4.660 ;
        RECT 1036.010 1.535 1038.590 4.660 ;
        RECT 1039.690 1.535 1042.270 4.660 ;
        RECT 1043.370 1.535 1045.950 4.660 ;
        RECT 1047.050 1.535 1049.630 4.660 ;
        RECT 1050.730 1.535 1053.310 5.340 ;
        RECT 1054.410 5.340 1082.750 6.700 ;
        RECT 1054.410 1.535 1056.990 5.340 ;
        RECT 1058.090 4.660 1082.750 5.340 ;
        RECT 1058.090 1.535 1060.670 4.660 ;
        RECT 1061.770 1.535 1064.350 4.660 ;
        RECT 1065.450 1.535 1068.030 4.660 ;
        RECT 1069.130 1.535 1071.710 4.660 ;
        RECT 1072.810 1.535 1075.390 4.660 ;
        RECT 1076.490 1.535 1079.070 4.660 ;
        RECT 1080.170 1.535 1082.750 4.660 ;
        RECT 1083.850 4.660 1101.150 7.380 ;
        RECT 1083.850 1.535 1086.430 4.660 ;
        RECT 1087.530 1.535 1090.110 4.660 ;
        RECT 1091.210 1.940 1101.150 4.660 ;
        RECT 1091.210 1.535 1093.790 1.940 ;
        RECT 1094.890 1.535 1097.470 1.940 ;
        RECT 1098.570 1.535 1101.150 1.940 ;
        RECT 1102.250 6.700 1115.870 7.380 ;
        RECT 1102.250 4.660 1112.190 6.700 ;
        RECT 1102.250 1.535 1104.830 4.660 ;
        RECT 1105.930 1.940 1112.190 4.660 ;
        RECT 1105.930 1.535 1108.510 1.940 ;
        RECT 1109.610 1.535 1112.190 1.940 ;
        RECT 1113.290 1.535 1115.870 6.700 ;
        RECT 1116.970 7.380 1123.230 14.180 ;
        RECT 1116.970 1.535 1119.550 7.380 ;
        RECT 1120.650 1.535 1123.230 7.380 ;
        RECT 1124.330 7.380 1130.590 14.180 ;
        RECT 1124.330 1.535 1126.910 7.380 ;
        RECT 1128.010 1.535 1130.590 7.380 ;
        RECT 1131.690 6.700 1178.430 14.180 ;
        RECT 1131.690 1.535 1134.270 6.700 ;
        RECT 1135.370 1.535 1137.950 6.700 ;
        RECT 1139.050 6.020 1178.430 6.700 ;
        RECT 1139.050 1.535 1141.630 6.020 ;
        RECT 1142.730 1.940 1156.350 6.020 ;
        RECT 1142.730 1.535 1145.310 1.940 ;
        RECT 1146.410 1.535 1148.990 1.940 ;
        RECT 1150.090 1.535 1152.670 1.940 ;
        RECT 1153.770 1.535 1156.350 1.940 ;
        RECT 1157.450 1.535 1160.030 6.020 ;
        RECT 1161.130 1.535 1163.710 6.020 ;
        RECT 1164.810 2.620 1178.430 6.020 ;
        RECT 1164.810 1.940 1174.750 2.620 ;
        RECT 1164.810 1.535 1167.390 1.940 ;
        RECT 1168.490 1.535 1171.070 1.940 ;
        RECT 1172.170 1.535 1174.750 1.940 ;
        RECT 1175.850 1.535 1178.430 2.620 ;
        RECT 1179.530 7.380 1187.265 14.180 ;
        RECT 1179.530 6.020 1185.790 7.380 ;
        RECT 1179.530 1.535 1182.110 6.020 ;
        RECT 1183.210 1.535 1185.790 6.020 ;
        RECT 1186.890 4.800 1187.265 7.380 ;
        RECT 1189.665 4.800 1356.255 49.600 ;
        RECT 1186.890 3.610 1357.165 4.800 ;
        RECT 1186.890 3.300 1290.210 3.610 ;
        RECT 1186.890 2.620 1249.730 3.300 ;
        RECT 1186.890 1.940 1205.570 2.620 ;
        RECT 1186.890 1.535 1198.210 1.940 ;
        RECT 1199.310 1.535 1201.890 1.940 ;
        RECT 1202.990 1.535 1205.570 1.940 ;
        RECT 1206.670 1.535 1209.250 2.620 ;
        RECT 1210.350 2.250 1216.610 2.620 ;
        RECT 1210.350 1.535 1212.930 2.250 ;
        RECT 1214.030 1.535 1216.610 2.250 ;
        RECT 1217.710 2.250 1223.970 2.620 ;
        RECT 1217.710 1.535 1220.290 2.250 ;
        RECT 1221.390 1.535 1223.970 2.250 ;
        RECT 1225.070 1.535 1227.650 2.620 ;
        RECT 1228.750 1.535 1231.330 2.620 ;
        RECT 1232.430 2.250 1242.370 2.620 ;
        RECT 1232.430 1.535 1235.010 2.250 ;
        RECT 1236.110 1.535 1238.690 2.250 ;
        RECT 1239.790 1.535 1242.370 2.250 ;
        RECT 1243.470 2.250 1249.730 2.620 ;
        RECT 1243.470 1.535 1246.050 2.250 ;
        RECT 1247.150 1.535 1249.730 2.250 ;
        RECT 1250.830 2.250 1257.090 3.300 ;
        RECT 1250.830 1.535 1253.410 2.250 ;
        RECT 1254.510 1.535 1257.090 2.250 ;
        RECT 1258.190 1.535 1260.770 3.300 ;
        RECT 1261.870 1.535 1264.450 3.300 ;
        RECT 1265.550 1.535 1268.130 3.300 ;
        RECT 1269.230 1.940 1275.490 3.300 ;
        RECT 1269.230 1.535 1271.810 1.940 ;
        RECT 1272.910 1.535 1275.490 1.940 ;
        RECT 1276.590 1.535 1279.170 3.300 ;
        RECT 1280.270 1.535 1282.850 3.300 ;
        RECT 1283.950 1.535 1286.530 3.300 ;
        RECT 1287.630 1.535 1290.210 3.300 ;
        RECT 1291.310 3.300 1357.165 3.610 ;
        RECT 1291.310 1.535 1293.890 3.300 ;
        RECT 1294.990 1.535 1297.570 3.300 ;
        RECT 1298.670 1.535 1301.250 3.300 ;
        RECT 1302.350 1.535 1304.930 3.300 ;
        RECT 1306.030 2.620 1312.290 3.300 ;
        RECT 1306.030 1.535 1308.610 2.620 ;
        RECT 1309.710 1.535 1312.290 2.620 ;
        RECT 1313.390 1.535 1315.970 3.300 ;
        RECT 1317.070 1.535 1319.650 3.300 ;
        RECT 1320.750 2.250 1327.010 3.300 ;
        RECT 1320.750 1.535 1323.330 2.250 ;
        RECT 1324.430 1.535 1327.010 2.250 ;
        RECT 1328.110 1.535 1330.690 3.300 ;
        RECT 1331.790 1.535 1334.370 3.300 ;
        RECT 1335.470 1.535 1338.050 3.300 ;
        RECT 1339.150 1.535 1341.730 3.300 ;
        RECT 1342.830 2.620 1349.090 3.300 ;
        RECT 1342.830 1.535 1345.410 2.620 ;
        RECT 1346.510 1.535 1349.090 2.620 ;
        RECT 1350.190 2.250 1357.165 3.300 ;
        RECT 1350.190 1.535 1352.770 2.250 ;
        RECT 1353.870 1.940 1357.165 2.250 ;
        RECT 1353.870 1.535 1356.450 1.940 ;
  END
END tt_mux
END LIBRARY

