* NGSPICE file created from tt_mux.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

.subckt tt_mux addr[0] addr[1] addr[2] addr[3] addr[4] k_one k_zero spine_iw[0] spine_iw[10]
+ spine_iw[11] spine_iw[12] spine_iw[13] spine_iw[14] spine_iw[15] spine_iw[16] spine_iw[17]
+ spine_iw[18] spine_iw[19] spine_iw[1] spine_iw[20] spine_iw[21] spine_iw[22] spine_iw[23]
+ spine_iw[24] spine_iw[25] spine_iw[26] spine_iw[27] spine_iw[28] spine_iw[29] spine_iw[2]
+ spine_iw[30] spine_iw[3] spine_iw[4] spine_iw[5] spine_iw[6] spine_iw[7] spine_iw[8]
+ spine_iw[9] spine_ow[0] spine_ow[10] spine_ow[11] spine_ow[12] spine_ow[13] spine_ow[14]
+ spine_ow[15] spine_ow[16] spine_ow[17] spine_ow[18] spine_ow[19] spine_ow[1] spine_ow[20]
+ spine_ow[21] spine_ow[22] spine_ow[23] spine_ow[24] spine_ow[25] spine_ow[2] spine_ow[3]
+ spine_ow[4] spine_ow[5] spine_ow[6] spine_ow[7] spine_ow[8] spine_ow[9] um_ena[0]
+ um_ena[10] um_ena[11] um_ena[12] um_ena[13] um_ena[14] um_ena[15] um_ena[1] um_ena[2]
+ um_ena[3] um_ena[4] um_ena[5] um_ena[6] um_ena[7] um_ena[8] um_ena[9] um_iw[0] um_iw[100]
+ um_iw[101] um_iw[102] um_iw[103] um_iw[104] um_iw[105] um_iw[106] um_iw[107] um_iw[108]
+ um_iw[109] um_iw[10] um_iw[110] um_iw[111] um_iw[112] um_iw[113] um_iw[114] um_iw[115]
+ um_iw[116] um_iw[117] um_iw[118] um_iw[119] um_iw[11] um_iw[120] um_iw[121] um_iw[122]
+ um_iw[123] um_iw[124] um_iw[125] um_iw[126] um_iw[127] um_iw[128] um_iw[129] um_iw[12]
+ um_iw[130] um_iw[131] um_iw[132] um_iw[133] um_iw[134] um_iw[135] um_iw[136] um_iw[137]
+ um_iw[138] um_iw[139] um_iw[13] um_iw[140] um_iw[141] um_iw[142] um_iw[143] um_iw[144]
+ um_iw[145] um_iw[146] um_iw[147] um_iw[148] um_iw[149] um_iw[14] um_iw[150] um_iw[151]
+ um_iw[152] um_iw[153] um_iw[154] um_iw[155] um_iw[156] um_iw[157] um_iw[158] um_iw[159]
+ um_iw[15] um_iw[160] um_iw[161] um_iw[162] um_iw[163] um_iw[164] um_iw[165] um_iw[166]
+ um_iw[167] um_iw[168] um_iw[169] um_iw[16] um_iw[170] um_iw[171] um_iw[172] um_iw[173]
+ um_iw[174] um_iw[175] um_iw[176] um_iw[177] um_iw[178] um_iw[179] um_iw[17] um_iw[180]
+ um_iw[181] um_iw[182] um_iw[183] um_iw[184] um_iw[185] um_iw[186] um_iw[187] um_iw[188]
+ um_iw[189] um_iw[18] um_iw[190] um_iw[191] um_iw[192] um_iw[193] um_iw[194] um_iw[195]
+ um_iw[196] um_iw[197] um_iw[198] um_iw[199] um_iw[19] um_iw[1] um_iw[200] um_iw[201]
+ um_iw[202] um_iw[203] um_iw[204] um_iw[205] um_iw[206] um_iw[207] um_iw[208] um_iw[209]
+ um_iw[20] um_iw[210] um_iw[211] um_iw[212] um_iw[213] um_iw[214] um_iw[215] um_iw[216]
+ um_iw[217] um_iw[218] um_iw[219] um_iw[21] um_iw[220] um_iw[221] um_iw[222] um_iw[223]
+ um_iw[224] um_iw[225] um_iw[226] um_iw[227] um_iw[228] um_iw[229] um_iw[22] um_iw[230]
+ um_iw[231] um_iw[232] um_iw[233] um_iw[234] um_iw[235] um_iw[236] um_iw[237] um_iw[238]
+ um_iw[239] um_iw[23] um_iw[240] um_iw[241] um_iw[242] um_iw[243] um_iw[244] um_iw[245]
+ um_iw[246] um_iw[247] um_iw[248] um_iw[249] um_iw[24] um_iw[250] um_iw[251] um_iw[252]
+ um_iw[253] um_iw[254] um_iw[255] um_iw[256] um_iw[257] um_iw[258] um_iw[259] um_iw[25]
+ um_iw[260] um_iw[261] um_iw[262] um_iw[263] um_iw[264] um_iw[265] um_iw[266] um_iw[267]
+ um_iw[268] um_iw[269] um_iw[26] um_iw[270] um_iw[271] um_iw[272] um_iw[273] um_iw[274]
+ um_iw[275] um_iw[276] um_iw[277] um_iw[278] um_iw[279] um_iw[27] um_iw[280] um_iw[281]
+ um_iw[282] um_iw[283] um_iw[284] um_iw[285] um_iw[286] um_iw[287] um_iw[28] um_iw[29]
+ um_iw[2] um_iw[30] um_iw[31] um_iw[32] um_iw[33] um_iw[34] um_iw[35] um_iw[36] um_iw[37]
+ um_iw[38] um_iw[39] um_iw[3] um_iw[40] um_iw[41] um_iw[42] um_iw[43] um_iw[44] um_iw[45]
+ um_iw[46] um_iw[47] um_iw[48] um_iw[49] um_iw[4] um_iw[50] um_iw[51] um_iw[52] um_iw[53]
+ um_iw[54] um_iw[55] um_iw[56] um_iw[57] um_iw[58] um_iw[59] um_iw[5] um_iw[60] um_iw[61]
+ um_iw[62] um_iw[63] um_iw[64] um_iw[65] um_iw[66] um_iw[67] um_iw[68] um_iw[69]
+ um_iw[6] um_iw[70] um_iw[71] um_iw[72] um_iw[73] um_iw[74] um_iw[75] um_iw[76] um_iw[77]
+ um_iw[78] um_iw[79] um_iw[7] um_iw[80] um_iw[81] um_iw[82] um_iw[83] um_iw[84] um_iw[85]
+ um_iw[86] um_iw[87] um_iw[88] um_iw[89] um_iw[8] um_iw[90] um_iw[91] um_iw[92] um_iw[93]
+ um_iw[94] um_iw[95] um_iw[96] um_iw[97] um_iw[98] um_iw[99] um_iw[9] um_k_zero[0]
+ um_k_zero[10] um_k_zero[11] um_k_zero[12] um_k_zero[13] um_k_zero[14] um_k_zero[15]
+ um_k_zero[1] um_k_zero[2] um_k_zero[3] um_k_zero[4] um_k_zero[5] um_k_zero[6] um_k_zero[7]
+ um_k_zero[8] um_k_zero[9] um_ow[0] um_ow[100] um_ow[101] um_ow[102] um_ow[103] um_ow[104]
+ um_ow[105] um_ow[106] um_ow[107] um_ow[108] um_ow[109] um_ow[10] um_ow[110] um_ow[111]
+ um_ow[112] um_ow[113] um_ow[114] um_ow[115] um_ow[116] um_ow[117] um_ow[118] um_ow[119]
+ um_ow[11] um_ow[120] um_ow[121] um_ow[122] um_ow[123] um_ow[124] um_ow[125] um_ow[126]
+ um_ow[127] um_ow[128] um_ow[129] um_ow[12] um_ow[130] um_ow[131] um_ow[132] um_ow[133]
+ um_ow[134] um_ow[135] um_ow[136] um_ow[137] um_ow[138] um_ow[139] um_ow[13] um_ow[140]
+ um_ow[141] um_ow[142] um_ow[143] um_ow[144] um_ow[145] um_ow[146] um_ow[147] um_ow[148]
+ um_ow[149] um_ow[14] um_ow[150] um_ow[151] um_ow[152] um_ow[153] um_ow[154] um_ow[155]
+ um_ow[156] um_ow[157] um_ow[158] um_ow[159] um_ow[15] um_ow[160] um_ow[161] um_ow[162]
+ um_ow[163] um_ow[164] um_ow[165] um_ow[166] um_ow[167] um_ow[168] um_ow[169] um_ow[16]
+ um_ow[170] um_ow[171] um_ow[172] um_ow[173] um_ow[174] um_ow[175] um_ow[176] um_ow[177]
+ um_ow[178] um_ow[179] um_ow[17] um_ow[180] um_ow[181] um_ow[182] um_ow[183] um_ow[184]
+ um_ow[185] um_ow[186] um_ow[187] um_ow[188] um_ow[189] um_ow[18] um_ow[190] um_ow[191]
+ um_ow[192] um_ow[193] um_ow[194] um_ow[195] um_ow[196] um_ow[197] um_ow[198] um_ow[199]
+ um_ow[19] um_ow[1] um_ow[200] um_ow[201] um_ow[202] um_ow[203] um_ow[204] um_ow[205]
+ um_ow[206] um_ow[207] um_ow[208] um_ow[209] um_ow[20] um_ow[210] um_ow[211] um_ow[212]
+ um_ow[213] um_ow[214] um_ow[215] um_ow[216] um_ow[217] um_ow[218] um_ow[219] um_ow[21]
+ um_ow[220] um_ow[221] um_ow[222] um_ow[223] um_ow[224] um_ow[225] um_ow[226] um_ow[227]
+ um_ow[228] um_ow[229] um_ow[22] um_ow[230] um_ow[231] um_ow[232] um_ow[233] um_ow[234]
+ um_ow[235] um_ow[236] um_ow[237] um_ow[238] um_ow[239] um_ow[23] um_ow[240] um_ow[241]
+ um_ow[242] um_ow[243] um_ow[244] um_ow[245] um_ow[246] um_ow[247] um_ow[248] um_ow[249]
+ um_ow[24] um_ow[250] um_ow[251] um_ow[252] um_ow[253] um_ow[254] um_ow[255] um_ow[256]
+ um_ow[257] um_ow[258] um_ow[259] um_ow[25] um_ow[260] um_ow[261] um_ow[262] um_ow[263]
+ um_ow[264] um_ow[265] um_ow[266] um_ow[267] um_ow[268] um_ow[269] um_ow[26] um_ow[270]
+ um_ow[271] um_ow[272] um_ow[273] um_ow[274] um_ow[275] um_ow[276] um_ow[277] um_ow[278]
+ um_ow[279] um_ow[27] um_ow[280] um_ow[281] um_ow[282] um_ow[283] um_ow[284] um_ow[285]
+ um_ow[286] um_ow[287] um_ow[288] um_ow[289] um_ow[28] um_ow[290] um_ow[291] um_ow[292]
+ um_ow[293] um_ow[294] um_ow[295] um_ow[296] um_ow[297] um_ow[298] um_ow[299] um_ow[29]
+ um_ow[2] um_ow[300] um_ow[301] um_ow[302] um_ow[303] um_ow[304] um_ow[305] um_ow[306]
+ um_ow[307] um_ow[308] um_ow[309] um_ow[30] um_ow[310] um_ow[311] um_ow[312] um_ow[313]
+ um_ow[314] um_ow[315] um_ow[316] um_ow[317] um_ow[318] um_ow[319] um_ow[31] um_ow[320]
+ um_ow[321] um_ow[322] um_ow[323] um_ow[324] um_ow[325] um_ow[326] um_ow[327] um_ow[328]
+ um_ow[329] um_ow[32] um_ow[330] um_ow[331] um_ow[332] um_ow[333] um_ow[334] um_ow[335]
+ um_ow[336] um_ow[337] um_ow[338] um_ow[339] um_ow[33] um_ow[340] um_ow[341] um_ow[342]
+ um_ow[343] um_ow[344] um_ow[345] um_ow[346] um_ow[347] um_ow[348] um_ow[349] um_ow[34]
+ um_ow[350] um_ow[351] um_ow[352] um_ow[353] um_ow[354] um_ow[355] um_ow[356] um_ow[357]
+ um_ow[358] um_ow[359] um_ow[35] um_ow[360] um_ow[361] um_ow[362] um_ow[363] um_ow[364]
+ um_ow[365] um_ow[366] um_ow[367] um_ow[368] um_ow[369] um_ow[36] um_ow[370] um_ow[371]
+ um_ow[372] um_ow[373] um_ow[374] um_ow[375] um_ow[376] um_ow[377] um_ow[378] um_ow[379]
+ um_ow[37] um_ow[380] um_ow[381] um_ow[382] um_ow[383] um_ow[38] um_ow[39] um_ow[3]
+ um_ow[40] um_ow[41] um_ow[42] um_ow[43] um_ow[44] um_ow[45] um_ow[46] um_ow[47]
+ um_ow[48] um_ow[49] um_ow[4] um_ow[50] um_ow[51] um_ow[52] um_ow[53] um_ow[54] um_ow[55]
+ um_ow[56] um_ow[57] um_ow[58] um_ow[59] um_ow[5] um_ow[60] um_ow[61] um_ow[62] um_ow[63]
+ um_ow[64] um_ow[65] um_ow[66] um_ow[67] um_ow[68] um_ow[69] um_ow[6] um_ow[70] um_ow[71]
+ um_ow[72] um_ow[73] um_ow[74] um_ow[75] um_ow[76] um_ow[77] um_ow[78] um_ow[79]
+ um_ow[7] um_ow[80] um_ow[81] um_ow[82] um_ow[83] um_ow[84] um_ow[85] um_ow[86] um_ow[87]
+ um_ow[88] um_ow[89] um_ow[8] um_ow[90] um_ow[91] um_ow[92] um_ow[93] um_ow[94] um_ow[95]
+ um_ow[96] um_ow[97] um_ow[98] um_ow[99] um_ow[9] vccd1 vssd1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_2673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[4\].zbuf_bot_iw_I\[10\].genblk1.cell0_I net507 col\[4\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[4\].zbuf_bot_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_224 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_213 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_202 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_432_ col\[7\].zbuf_bot_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[255] sky130_fd_sc_hd__buf_2
XANTENNA_246 col\[0\].genblk1.tbuf_spine_ow_I\[17\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_257 col\[0\].genblk1.tbuf_spine_ow_I\[2\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_235 _013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_2183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_268 col\[0\].genblk1.tbuf_spine_ow_I\[2\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_279 col\[0\].genblk1.tbuf_spine_ow_I\[3\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_2093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_363_ col\[5\].zbuf_bot_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[186] sky130_fd_sc_hd__buf_2
XFILLER_0_7_1493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_294_ col\[3\].zbuf_bot_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[117] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_2879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.mux4_I\[17\].cell0_I net263 net289 net316 net342 net472 net458 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[17\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_11_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_2233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_2289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_415_ col\[6\].zbuf_top_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[238] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_346_ col\[4\].zbuf_top_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[169] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_277_ col\[2\].zbuf_top_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[100] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[0\].zbuf_bot_iw_I\[5\].genblk1.cell0_I net483 col\[0\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[0\].zbuf_bot_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[4\].genblk1.mux4_I\[8\].cell0_I net147 net173 net199 net226 net468 net454 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[8\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_14_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].zbuf_bot_iw_I\[0\].genblk1.cell0_I net509 col\[2\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[2\].zbuf_bot_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XFILLER_0_15_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_200_ col\[0\].zbuf_top_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[23] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_2085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_062_ _009_ vssd1 vssd1 vccd1 vccd1 tbuf_row_ena_I.t sky130_fd_sc_hd__clkbuf_1
Xfanout480 col\[0\].zbuf_bot_iw_I\[7\].a vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_4
Xfanout491 col\[0\].zbuf_bot_iw_I\[1\].a vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__buf_8
Xcol\[0\].genblk1.mux4_I\[6\].cell0_I net385 net268 net368 net394 net462 net448 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[6\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_329_ col\[4\].zbuf_bot_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[152] sky130_fd_sc_hd__buf_2
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_2462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[3\].zbuf_top_iw_I\[17\].genblk1.cell0_I net493 net427 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_2237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[3\].zbuf_bot_iw_I\[8\].genblk1.cell0_I net477 col\[3\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[3\].zbuf_bot_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_1989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[5\].zbuf_bot_iw_I\[3\].genblk1.cell0_I net488 col\[5\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[5\].zbuf_bot_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput301 um_ow[33] vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_2
Xinput312 um_ow[34] vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__clkbuf_2
Xinput334 um_ow[36] vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput345 um_ow[37] vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__clkbuf_2
Xinput323 um_ow[35] vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__clkbuf_2
Xinput356 um_ow[43] vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__clkbuf_2
Xinput378 um_ow[63] vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_1
Xinput367 um_ow[53] vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__clkbuf_1
Xinput389 um_ow[73] vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_2001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.tbuf_spine_ow_I\[21\].cell0_I col\[4\].genblk1.mux4_I\[21\].x net438
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[21\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_10_2854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_5 col\[0\].genblk1.tbuf_spine_ow_I\[0\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_2811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_2866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[5\].zbuf_top_iw_I\[16\].genblk1.cell0_I net496 net423 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[16\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_iw_I\[7\].genblk1.cell0_I net479 net432 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.mux4_I\[9\].cell0_I net41 net67 net94 net120 net466 net452 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[9\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_7_2365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[3\].zbuf_top_iw_I\[2\].genblk1.cell0_I net489 net428 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[0\].genblk1.tbuf_spine_ow_I\[17\].cell0_I col\[0\].genblk1.mux4_I\[17\].x net445
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[17\].z sky130_fd_sc_hd__ebufn_8
Xinput120 um_ow[177] vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__clkbuf_1
Xinput131 um_ow[187] vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__clkbuf_1
Xinput142 um_ow[197] vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_1
Xinput153 um_ow[206] vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__clkbuf_1
Xinput175 um_ow[226] vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_1
Xinput186 um_ow[236] vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_1
Xinput164 um_ow[216] vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_1
Xinput197 um_ow[246] vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__dlymetal6s2s_1
Xtbuf_spine_ow_I\[15\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[15\].z net511 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[15\].z sky130_fd_sc_hd__ebufn_1
XFILLER_0_15_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].genblk1.mux4_I\[12\].cell0_I net44 net71 net97 net124 net465 net451 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[12\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_15_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xzbuf_bus_sel_I\[4\].genblk1.cell0_I net30 net516 vssd1 vssd1 vccd1 vccd1 zbuf_bus_sel_I\[4\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_10_2673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_2641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_225 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_214 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_203 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_247 col\[0\].genblk1.tbuf_spine_ow_I\[18\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_431_ col\[7\].zbuf_bot_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[254] sky130_fd_sc_hd__buf_2
XFILLER_0_3_2015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_258 col\[0\].genblk1.tbuf_spine_ow_I\[2\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_236 col\[0\].genblk1.tbuf_spine_ow_I\[10\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_362_ col\[5\].zbuf_bot_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[185] sky130_fd_sc_hd__buf_2
XANTENNA_269 col\[0\].genblk1.tbuf_spine_ow_I\[2\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_293_ col\[3\].zbuf_bot_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[116] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_top_iw_I\[15\].genblk1.cell0_I net498 net419 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[4\].genblk1.mux4_I\[22\].cell0_I net162 net188 net215 net241 net469 net455 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[22\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_14_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[6\].zbuf_top_iw_I\[5\].genblk1.cell0_I net484 net422 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_414_ col\[6\].zbuf_top_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[237] sky130_fd_sc_hd__buf_2
X_345_ col\[4\].zbuf_top_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[168] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_276_ col\[2\].zbuf_top_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[99] sky130_fd_sc_hd__buf_2
XFILLER_0_14_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_2909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_2554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_2029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_061_ _003_ _006_ _008_ vssd1 vssd1 vccd1 vccd1 _009_ sky130_fd_sc_hd__and3_1
Xfanout481 col\[0\].zbuf_bot_iw_I\[6\].a vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__buf_6
Xfanout470 net474 vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__clkbuf_4
Xfanout492 col\[0\].zbuf_bot_iw_I\[1\].a vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__clkbuf_4
Xcol\[4\].genblk1.tbuf_spine_ow_I\[1\].cell0_I col\[4\].genblk1.mux4_I\[1\].x net439
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[1\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_6_2920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_328_ col\[4\].zbuf_bot_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[151] sky130_fd_sc_hd__buf_2
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_259_ col\[2\].zbuf_bot_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[82] sky130_fd_sc_hd__buf_2
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].genblk1.tbuf_spine_ow_I\[10\].cell0_I col\[2\].genblk1.mux4_I\[10\].x net442
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[10\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_2205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_2249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xzbuf_bus_ena_I.genblk1.cell0_I net16 net516 vssd1 vssd1 vccd1 vccd1 zbuf_bus_ena_I.genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_2_2603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_2750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput302 um_ow[340] vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput335 um_ow[370] vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput324 um_ow[360] vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput313 um_ow[350] vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput346 um_ow[380] vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput357 um_ow[44] vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__clkbuf_2
Xinput379 um_ow[64] vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__clkbuf_1
Xinput368 um_ow[54] vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_2013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_6 col\[0\].genblk1.tbuf_spine_ow_I\[0\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[0\].zbuf_top_iw_I\[16\].genblk1.cell0_I net495 net433 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_2709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_2580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[3\].zbuf_bot_ena_I.genblk1.cell0_I net542 col\[3\].zbuf_bot_ena_I.e vssd1 vssd1
+ vccd1 vccd1 col\[3\].zbuf_bot_ena_I.z sky130_fd_sc_hd__and2_1
XFILLER_0_14_1520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput110 um_ow[168] vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_1
Xinput121 um_ow[178] vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_1
Xinput132 um_ow[188] vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_1
Xinput143 um_ow[198] vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_1
Xinput154 um_ow[207] vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__clkbuf_1
Xinput165 um_ow[217] vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_1
Xinput176 um_ow[227] vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_1
Xinput187 um_ow[237] vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_1
Xinput198 um_ow[247] vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_15_2029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtbuf_spine_ow_I\[19\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[19\].z net511 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[19\].z sky130_fd_sc_hd__ebufn_1
Xcol\[2\].genblk1.mux4_I\[16\].cell0_I net49 net75 net102 net128 net464 net450 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[16\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_13_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_2641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_2685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[1\].zbuf_bot_iw_I\[0\].genblk1.cell0_I net509 col\[1\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[1\].zbuf_bot_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_2653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_2697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_2252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[14\].genblk1.cell1_I zbuf_bus_iw_I\[14\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[14\].a sky130_fd_sc_hd__buf_6
XFILLER_0_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_204 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_2141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_215 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_226 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_248 col\[0\].genblk1.tbuf_spine_ow_I\[18\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_430_ col\[7\].zbuf_bot_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[253] sky130_fd_sc_hd__buf_2
XANTENNA_237 col\[0\].genblk1.tbuf_spine_ow_I\[17\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_259 col\[0\].genblk1.tbuf_spine_ow_I\[2\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_361_ col\[5\].zbuf_bot_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[184] sky130_fd_sc_hd__buf_2
XFILLER_0_7_2185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[2\].zbuf_top_iw_I\[15\].genblk1.cell0_I net497 net429 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_292_ col\[3\].zbuf_bot_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[115] sky130_fd_sc_hd__buf_2
XFILLER_0_1_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].genblk1.tbuf_spine_ow_I\[0\].cell0_I col\[0\].genblk1.mux4_I\[0\].x net444
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[0\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_8_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].zbuf_bot_iw_I\[17\].genblk1.cell0_I net494 col\[6\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[6\].zbuf_bot_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_1513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_413_ col\[6\].zbuf_top_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[236] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xzbuf_bus_iw_I\[1\].genblk1.cell1_I zbuf_bus_iw_I\[1\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[1\].a sky130_fd_sc_hd__buf_6
XFILLER_0_12_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_344_ col\[4\].zbuf_top_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[167] sky130_fd_sc_hd__buf_2
X_275_ col\[2\].zbuf_top_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[98] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].zbuf_bot_iw_I\[8\].genblk1.cell0_I net477 col\[2\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[2\].zbuf_bot_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_10_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_2781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_bot_iw_I\[3\].genblk1.cell0_I net487 col\[4\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[4\].zbuf_bot_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_15_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[4\].zbuf_top_iw_I\[14\].genblk1.cell0_I net499 net425 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_060_ net4 _004_ net1 _005_ _007_ vssd1 vssd1 vccd1 vccd1 _008_ sky130_fd_sc_hd__a221oi_1
Xfanout482 col\[0\].zbuf_bot_iw_I\[6\].a vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__clkbuf_4
Xfanout493 col\[0\].zbuf_bot_iw_I\[17\].a vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__buf_6
Xfanout460 zbuf_bus_sel_I\[1\].z vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_2
Xfanout471 net474 vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__buf_4
XFILLER_0_9_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[4\].genblk1.tbuf_spine_ow_I\[5\].cell0_I col\[4\].genblk1.mux4_I\[5\].x net439
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[5\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_13_2875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_327_ col\[4\].zbuf_bot_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[150] sky130_fd_sc_hd__buf_2
Xcol\[0\].zbuf_top_iw_I\[7\].genblk1.cell0_I net479 net433 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_2597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_258_ col\[2\].zbuf_bot_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[81] sky130_fd_sc_hd__buf_2
XFILLER_0_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_189_ col\[0\].zbuf_bot_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[12] sky130_fd_sc_hd__buf_2
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.tbuf_spine_ow_I\[14\].cell0_I col\[2\].genblk1.mux4_I\[14\].x net441
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[14\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_14_2628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_2617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[2\].zbuf_top_iw_I\[2\].genblk1.cell0_I net489 net430 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_1605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[7\].zbuf_top_ena_I.genblk1.cell0_I net551 net420 vssd1 vssd1 vccd1 vccd1 col\[7\].zbuf_top_ena_I.z
+ sky130_fd_sc_hd__and2_1
XFILLER_0_1_1649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[6\].zbuf_top_iw_I\[13\].genblk1.cell0_I net502 net421 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[10\].genblk1.cell0_I net19 net515 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[10\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_0_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[7\].zbuf_bot_iw_I\[6\].genblk1.cell0_I net482 col\[7\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[7\].zbuf_bot_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_2136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput303 um_ow[341] vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput325 um_ow[361] vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput336 um_ow[371] vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput314 um_ow[351] vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput347 um_ow[381] vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput358 um_ow[45] vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__clkbuf_2
Xinput369 um_ow[55] vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_2025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_2069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_7 col\[0\].genblk1.tbuf_spine_ow_I\[0\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_2824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_2200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[5\].zbuf_top_iw_I\[5\].genblk1.cell0_I net484 net424 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput111 um_ow[169] vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_1
Xinput100 um_ow[159] vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_1
Xinput122 um_ow[179] vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__clkbuf_1
Xinput133 um_ow[189] vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_1
Xinput144 um_ow[199] vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_1
Xinput166 um_ow[218] vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_1
Xinput177 um_ow[228] vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_1
Xinput155 um_ow[208] vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__clkbuf_1
Xcol\[7\].zbuf_top_iw_I\[0\].genblk1.cell0_I net510 net420 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[0\].z sky130_fd_sc_hd__and2_1
Xinput188 um_ow[238] vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_1
Xcol\[0\].genblk1.mux4_I\[21\].cell0_I net168 net358 net384 net411 net461 net447 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[21\].x sky130_fd_sc_hd__mux4_2
Xinput199 um_ow[248] vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_8_1408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_2653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_216 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_205 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_227 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_238 col\[0\].genblk1.tbuf_spine_ow_I\[17\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_249 col\[0\].genblk1.tbuf_spine_ow_I\[18\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_2153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_360_ col\[5\].zbuf_bot_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[183] sky130_fd_sc_hd__buf_2
XFILLER_0_3_2017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_291_ col\[3\].zbuf_bot_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[114] sky130_fd_sc_hd__buf_2
XFILLER_0_9_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[0\].genblk1.tbuf_spine_ow_I\[4\].cell0_I col\[0\].genblk1.mux4_I\[4\].x net444
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_3_1861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtbuf_spine_ow_I\[1\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[1\].z net512 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[1\].z sky130_fd_sc_hd__ebufn_1
XFILLER_0_15_2372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[1\].zbuf_bot_iw_I\[17\].genblk1.cell0_I net493 col\[1\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[1\].zbuf_bot_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_2061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_412_ col\[6\].zbuf_top_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[235] sky130_fd_sc_hd__buf_2
XFILLER_0_9_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_343_ col\[4\].zbuf_top_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[166] sky130_fd_sc_hd__buf_2
X_274_ col\[2\].zbuf_top_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[97] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_2793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_2523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[6\].genblk1.tbuf_spine_ow_I\[22\].cell0_I col\[6\].genblk1.mux4_I\[22\].x net435
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[22\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtt_mux_530 vssd1 vssd1 vccd1 vccd1 tt_mux_530/HI um_k_zero[10] sky130_fd_sc_hd__conb_1
XFILLER_0_13_2309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtt_mux_552 vssd1 vssd1 vccd1 vccd1 k_one tt_mux_552/LO sky130_fd_sc_hd__conb_1
XFILLER_0_15_2191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout450 net453 vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__buf_2
Xfanout483 col\[0\].zbuf_bot_iw_I\[5\].a vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__buf_6
Xfanout472 net474 vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__clkbuf_2
Xfanout461 net463 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__buf_4
Xfanout494 col\[0\].zbuf_bot_iw_I\[17\].a vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_2911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_326_ col\[4\].zbuf_bot_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[149] sky130_fd_sc_hd__buf_2
Xcol\[4\].genblk1.tbuf_spine_ow_I\[9\].cell0_I col\[4\].genblk1.mux4_I\[9\].x net439
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[9\].z sky130_fd_sc_hd__ebufn_8
X_257_ col\[2\].zbuf_bot_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[80] sky130_fd_sc_hd__buf_2
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_188_ col\[0\].zbuf_bot_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[11] sky130_fd_sc_hd__buf_2
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[3\].zbuf_bot_iw_I\[16\].genblk1.cell0_I net495 col\[3\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[3\].zbuf_bot_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[2\].genblk1.tbuf_spine_ow_I\[18\].cell0_I col\[2\].genblk1.mux4_I\[18\].x net441
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[18\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_5_2421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[0\].zbuf_bot_iw_I\[0\].genblk1.cell0_I net509 col\[0\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[0\].zbuf_bot_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[1\].zbuf_top_iw_I\[13\].genblk1.cell0_I net501 net431 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_sel_I\[3\].genblk1.cell1_I zbuf_bus_sel_I\[3\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 zbuf_bus_sel_I\[3\].z sky130_fd_sc_hd__buf_6
XFILLER_0_13_1961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_309_ col\[3\].zbuf_top_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[132] sky130_fd_sc_hd__buf_2
XFILLER_0_13_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput326 um_ow[362] vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput304 um_ow[342] vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput315 um_ow[352] vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput348 um_ow[382] vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput359 um_ow[46] vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__clkbuf_2
Xinput337 um_ow[372] vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__dlymetal6s2s_1
Xcol\[5\].zbuf_bot_iw_I\[15\].genblk1.cell0_I net498 col\[5\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[5\].zbuf_bot_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_2903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_2846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_8 col\[0\].genblk1.tbuf_spine_ow_I\[0\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_2713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_2757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[3\].zbuf_top_iw_I\[12\].genblk1.cell0_I net503 net427 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_2335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_2070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[1\].zbuf_bot_iw_I\[8\].genblk1.cell0_I net477 col\[1\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[1\].zbuf_bot_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput101 um_ow[15] vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_2
Xinput112 um_ow[16] vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__clkbuf_2
Xinput123 um_ow[17] vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput134 um_ow[18] vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput145 um_ow[19] vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput167 um_ow[219] vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_1
Xinput178 um_ow[229] vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_1
Xinput156 um_ow[209] vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_1
Xinput189 um_ow[239] vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_1
Xcol\[3\].zbuf_bot_iw_I\[3\].genblk1.cell0_I net487 col\[3\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[3\].zbuf_bot_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_2532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_2210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[7\].zbuf_bot_iw_I\[14\].genblk1.cell0_I net500 col\[7\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[7\].zbuf_bot_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_11_1717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.tbuf_spine_ow_I\[11\].cell0_I col\[4\].genblk1.mux4_I\[11\].x net438
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[11\].z sky130_fd_sc_hd__ebufn_8
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_206 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_217 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_228 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_239 col\[0\].genblk1.tbuf_spine_ow_I\[17\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_2165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_290_ col\[3\].zbuf_bot_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[113] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[5\].zbuf_top_iw_I\[11\].genblk1.cell0_I net506 net423 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[11\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_iw_I\[2\].genblk1.cell0_I net489 net432 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_15_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_2574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[0\].genblk1.tbuf_spine_ow_I\[8\].cell0_I col\[0\].genblk1.mux4_I\[8\].x net445
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_3_1873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xzbuf_bus_iw_I\[9\].genblk1.cell1_I zbuf_bus_iw_I\[9\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[9\].a sky130_fd_sc_hd__buf_6
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xtbuf_spine_ow_I\[5\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[5\].z net512 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[5\].z sky130_fd_sc_hd__ebufn_2
XFILLER_0_11_1525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_411_ col\[6\].zbuf_top_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[234] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_342_ col\[4\].zbuf_top_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[165] sky130_fd_sc_hd__buf_2
X_273_ col\[2\].zbuf_top_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[96] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_2793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[6\].zbuf_bot_iw_I\[6\].genblk1.cell0_I net482 col\[6\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[6\].zbuf_bot_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_12_2535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtt_mux_531 vssd1 vssd1 vccd1 vccd1 tt_mux_531/HI um_k_zero[11] sky130_fd_sc_hd__conb_1
Xtt_mux_520 vssd1 vssd1 vccd1 vccd1 tt_mux_520/HI um_k_zero[0] sky130_fd_sc_hd__conb_1
XFILLER_0_4_2113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[7\].zbuf_top_iw_I\[10\].genblk1.cell0_I net508 net419 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout440 col\[4\].genblk1.tbuf_row_ena_I.tx vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__buf_6
Xfanout484 col\[0\].zbuf_bot_iw_I\[5\].a vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__clkbuf_4
Xfanout462 net463 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__buf_4
Xfanout473 net474 vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__clkbuf_4
Xcol\[4\].genblk1.mux4_I\[12\].cell0_I net151 net177 net204 net230 net468 net454 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[12\].x sky130_fd_sc_hd__mux4_1
Xfanout451 net453 vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__clkbuf_2
Xfanout495 col\[0\].zbuf_bot_iw_I\[16\].a vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_6
XFILLER_0_9_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_2899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_325_ col\[4\].zbuf_bot_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[148] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_256_ col\[2\].zbuf_bot_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[79] sky130_fd_sc_hd__buf_2
X_187_ col\[0\].zbuf_bot_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[10] sky130_fd_sc_hd__buf_2
XFILLER_0_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[4\].zbuf_top_iw_I\[5\].genblk1.cell0_I net483 net426 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_2488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].zbuf_top_iw_I\[0\].genblk1.cell0_I net510 net422 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_2129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.mux4_I\[22\].cell0_I net269 net295 net321 net348 net471 net457 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[22\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_13_1973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_2330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_308_ col\[3\].zbuf_top_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[131] sky130_fd_sc_hd__buf_2
X_239_ col\[1\].zbuf_top_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[62] sky130_fd_sc_hd__buf_2
XFILLER_0_13_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_2427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].zbuf_bot_iw_I\[15\].genblk1.cell0_I net497 col\[0\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[0\].zbuf_bot_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput327 um_ow[363] vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput305 um_ow[343] vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput316 um_ow[353] vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput338 um_ow[373] vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput349 um_ow[383] vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_9 col\[0\].genblk1.tbuf_spine_ow_I\[0\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_2561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xzbuf_bus_iw_I\[5\].genblk1.cell0_I net13 net514 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[5\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_13_2471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[7\].zbuf_top_iw_I\[8\].genblk1.cell0_I net478 net420 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput102 um_ow[160] vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_1
Xinput113 um_ow[170] vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__clkbuf_1
Xinput135 um_ow[190] vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__clkbuf_1
Xinput124 um_ow[180] vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__clkbuf_1
Xinput146 um_ow[1] vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__clkbuf_2
Xinput157 um_ow[20] vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_2
Xinput168 um_ow[21] vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput179 um_ow[22] vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_15_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_2701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[2\].zbuf_bot_iw_I\[14\].genblk1.cell0_I net499 col\[2\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[2\].zbuf_bot_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_1933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[4\].genblk1.tbuf_spine_ow_I\[15\].cell0_I col\[4\].genblk1.mux4_I\[15\].x net440
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[15\].z sky130_fd_sc_hd__ebufn_8
XANTENNA_207 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_218 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_229 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_2177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_2907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_2920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].zbuf_top_iw_I\[11\].genblk1.cell0_I net505 net433 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_2829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_2330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtbuf_spine_ow_I\[9\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[9\].z net513 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[9\].z sky130_fd_sc_hd__ebufn_1
XFILLER_0_13_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_2239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_410_ col\[6\].zbuf_bot_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[233] sky130_fd_sc_hd__buf_2
X_341_ col\[4\].zbuf_top_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[164] sky130_fd_sc_hd__buf_2
Xcol\[4\].zbuf_bot_iw_I\[13\].genblk1.cell0_I net501 col\[4\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[4\].zbuf_bot_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_2895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_272_ col\[2\].zbuf_top_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[95] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_2637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_2547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_2350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtt_mux_521 vssd1 vssd1 vccd1 vccd1 tt_mux_521/HI um_k_zero[1] sky130_fd_sc_hd__conb_1
Xtt_mux_532 vssd1 vssd1 vccd1 vccd1 tt_mux_532/HI um_k_zero[12] sky130_fd_sc_hd__conb_1
Xcol\[2\].zbuf_top_iw_I\[10\].genblk1.cell0_I net507 net429 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_2125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[0\].genblk1.tbuf_spine_ow_I\[22\].cell0_I col\[0\].genblk1.mux4_I\[22\].x net444
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[22\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_11_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtbuf_spine_ow_I\[20\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[20\].z net511 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[20\].z sky130_fd_sc_hd__ebufn_2
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout430 col\[2\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout441 net443 vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__buf_12
Xfanout463 net467 vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__clkbuf_4
Xfanout452 net453 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__buf_2
Xfanout474 zbuf_bus_sel_I\[0\].z vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__clkbuf_4
Xfanout485 col\[0\].zbuf_bot_iw_I\[4\].a vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_8
Xfanout496 col\[0\].zbuf_bot_iw_I\[16\].a vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_2047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[16\].cell0_I net155 net182 net208 net235 net469 net455 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[16\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_6_2935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_324_ col\[4\].zbuf_bot_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[147] sky130_fd_sc_hd__buf_2
X_255_ col\[2\].zbuf_bot_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[78] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_186_ col\[0\].zbuf_bot_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[9] sky130_fd_sc_hd__buf_2
Xcol\[6\].genblk1.tbuf_spine_ow_I\[1\].cell0_I col\[6\].genblk1.mux4_I\[1\].x net436
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[1\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_5_2401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_2333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.tbuf_row_ena_I.cell0_I col\[6\].genblk1.tbuf_row_ena_I.t vssd1 vssd1
+ vccd1 vccd1 col\[6\].genblk1.tbuf_row_ena_I.tx sky130_fd_sc_hd__clkinv_4
XFILLER_0_12_1621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].zbuf_bot_iw_I\[8\].genblk1.cell0_I net477 col\[0\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[0\].zbuf_bot_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[6\].zbuf_bot_iw_I\[12\].genblk1.cell0_I net504 col\[6\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[6\].zbuf_bot_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].zbuf_bot_iw_I\[3\].genblk1.cell0_I net487 col\[2\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[2\].zbuf_bot_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_2765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_2629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_307_ col\[3\].zbuf_top_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[130] sky130_fd_sc_hd__buf_2
XFILLER_0_13_2697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_238_ col\[1\].zbuf_top_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[61] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_169_ col\[4\].zbuf_bot_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[8] sky130_fd_sc_hd__buf_2
XFILLER_0_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput306 um_ow[344] vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput317 um_ow[354] vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput328 um_ow[364] vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput339 um_ow[374] vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__dlymetal6s2s_1
Xcol\[0\].zbuf_top_iw_I\[2\].genblk1.cell0_I net489 net434 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_10_2815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_2826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_2426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_2459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_2225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[3\].zbuf_top_ena_I.genblk1.cell0_I net543 net428 vssd1 vssd1 vccd1 vccd1 col\[3\].zbuf_top_ena_I.z
+ sky130_fd_sc_hd__and2_1
XFILLER_0_1_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput114 um_ow[171] vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkbuf_1
Xinput125 um_ow[181] vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_1
Xinput136 um_ow[191] vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_1
Xinput103 um_ow[161] vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_1
Xinput169 um_ow[220] vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_1
Xinput147 um_ow[200] vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_1
Xinput158 um_ow[210] vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__clkbuf_1
Xcol\[5\].zbuf_bot_iw_I\[6\].genblk1.cell0_I net482 col\[5\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[5\].zbuf_bot_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_2713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_2757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[7\].zbuf_bot_iw_I\[1\].genblk1.cell0_I net492 col\[7\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[7\].zbuf_bot_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_1901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_219 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_208 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_2009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[4\].genblk1.tbuf_spine_ow_I\[19\].cell0_I col\[4\].genblk1.mux4_I\[19\].x net438
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[19\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_7_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_top_ena_I.genblk1.cell0_I_537 vssd1 vssd1 vccd1 vccd1 net537 col\[0\].zbuf_top_ena_I.genblk1.cell0_I_537/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_9_2911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[3\].zbuf_top_iw_I\[5\].genblk1.cell0_I net483 net428 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.tbuf_spine_ow_I\[0\].cell0_I col\[2\].genblk1.mux4_I\[0\].x net442
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[0\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[5\].zbuf_top_iw_I\[0\].genblk1.cell0_I net510 net424 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_2318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_2097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].genblk1.mux4_I\[11\].cell0_I net57 net323 net373 net400 net462 net448 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[11\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_6_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_340_ col\[4\].zbuf_top_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[163] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_271_ col\[2\].zbuf_top_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[94] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_2261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtt_mux_522 vssd1 vssd1 vccd1 vccd1 tt_mux_522/HI um_k_zero[2] sky130_fd_sc_hd__conb_1
Xtt_mux_533 vssd1 vssd1 vccd1 vccd1 tt_mux_533/HI um_k_zero[13] sky130_fd_sc_hd__conb_1
XFILLER_0_4_2137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout420 col\[7\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout431 col\[1\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__clkbuf_2
Xcol\[2\].genblk1.mux4_I\[21\].cell0_I net54 net81 net107 net133 net464 net450 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[21\].x sky130_fd_sc_hd__mux4_1
Xfanout475 col\[0\].zbuf_bot_iw_I\[9\].a vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__buf_6
Xfanout453 zbuf_bus_sel_I\[1\].z vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_4
Xfanout442 net443 vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__buf_12
Xfanout464 net465 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__clkbuf_4
Xfanout486 col\[0\].zbuf_bot_iw_I\[4\].a vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__clkbuf_4
Xfanout497 col\[0\].zbuf_bot_iw_I\[15\].a vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__buf_6
XFILLER_0_9_2015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_2059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_323_ col\[4\].zbuf_bot_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[146] sky130_fd_sc_hd__buf_2
X_254_ col\[2\].zbuf_bot_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[77] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_2535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_185_ col\[0\].zbuf_bot_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[8] sky130_fd_sc_hd__buf_2
Xcol\[6\].genblk1.tbuf_spine_ow_I\[5\].cell0_I col\[6\].genblk1.mux4_I\[5\].x net436
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[5\].z sky130_fd_sc_hd__ebufn_8
Xcol\[6\].zbuf_top_iw_I\[8\].genblk1.cell0_I net478 net421 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[8\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_ena_I.genblk1.cell0_I_539 vssd1 vssd1 vccd1 vccd1 net539 col\[1\].zbuf_top_ena_I.genblk1.cell0_I_539/LO
+ sky130_fd_sc_hd__conb_1
Xcol\[1\].zbuf_bot_iw_I\[12\].genblk1.cell0_I net503 col\[1\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[1\].zbuf_bot_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_2424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[6\].genblk1.tbuf_spine_ow_I\[12\].cell0_I col\[6\].genblk1.mux4_I\[12\].x net435
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[12\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_9_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_306_ col\[3\].zbuf_top_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[129] sky130_fd_sc_hd__buf_2
XFILLER_0_2_1918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_237_ col\[1\].zbuf_top_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[60] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_168_ col\[3\].zbuf_top_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[7] sky130_fd_sc_hd__buf_2
X_099_ _013_ _011_ _028_ vssd1 vssd1 vccd1 vccd1 _031_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput307 um_ow[345] vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__clkbuf_2
Xinput318 um_ow[355] vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput329 um_ow[365] vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_6_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[3\].zbuf_bot_iw_I\[11\].genblk1.cell0_I net505 col\[3\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[3\].zbuf_bot_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_2541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_2237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput115 um_ow[172] vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__clkbuf_1
Xinput126 um_ow[182] vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_1
Xinput104 um_ow[162] vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_1
Xinput148 um_ow[201] vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__clkbuf_1
Xinput159 um_ow[211] vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__clkbuf_1
Xinput137 um_ow[192] vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_2725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_2883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_2769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_2603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[5\].zbuf_bot_iw_I\[10\].genblk1.cell0_I net508 col\[5\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[5\].zbuf_bot_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_2001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_209 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_2533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_2577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[2\].genblk1.tbuf_spine_ow_I\[4\].cell0_I col\[2\].genblk1.mux4_I\[4\].x net442
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_8_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[1\].zbuf_bot_iw_I\[3\].genblk1.cell0_I net487 col\[1\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[1\].zbuf_bot_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_1765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[0\].genblk1.mux4_I\[15\].cell0_I net101 net351 net378 net404 net461 net447 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[15\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_10_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_2717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xzbuf_bus_iw_I\[17\].genblk1.cell1_I zbuf_bus_iw_I\[17\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[17\].a sky130_fd_sc_hd__buf_6
X_270_ col\[2\].zbuf_top_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[93] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_2606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_2363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_399_ col\[6\].zbuf_bot_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[222] sky130_fd_sc_hd__buf_2
XFILLER_0_3_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtt_mux_523 vssd1 vssd1 vccd1 vccd1 tt_mux_523/HI um_k_zero[3] sky130_fd_sc_hd__conb_1
Xtt_mux_534 vssd1 vssd1 vccd1 vccd1 tt_mux_534/HI um_k_zero[14] sky130_fd_sc_hd__conb_1
XFILLER_0_15_2151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout421 col\[6\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__clkbuf_2
Xfanout432 col\[1\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout454 net455 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__buf_2
Xfanout443 col\[2\].genblk1.tbuf_row_ena_I.tx vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__buf_6
Xfanout465 net467 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__buf_2
Xfanout476 col\[0\].zbuf_bot_iw_I\[9\].a vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__clkbuf_4
Xfanout498 col\[0\].zbuf_bot_iw_I\[15\].a vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__clkbuf_4
Xfanout487 col\[0\].zbuf_bot_iw_I\[3\].a vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__buf_8
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_322_ col\[4\].zbuf_bot_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[145] sky130_fd_sc_hd__buf_2
XFILLER_0_4_2661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_253_ col\[2\].zbuf_bot_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[76] sky130_fd_sc_hd__buf_2
X_184_ col\[0\].zbuf_bot_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[7] sky130_fd_sc_hd__buf_2
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.mux4_I\[2\].cell0_I net246 net273 net299 net326 net474 net459 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[2\].x sky130_fd_sc_hd__mux4_1
Xcol\[6\].genblk1.tbuf_spine_ow_I\[9\].cell0_I col\[6\].genblk1.mux4_I\[9\].x net435
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[9\].z sky130_fd_sc_hd__ebufn_8
Xzbuf_bus_iw_I\[4\].genblk1.cell1_I zbuf_bus_iw_I\[4\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[4\].a sky130_fd_sc_hd__buf_6
XFILLER_0_5_2447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[4\].zbuf_bot_iw_I\[6\].genblk1.cell0_I net481 col\[4\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[4\].zbuf_bot_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[4\].zbuf_top_iw_I\[17\].genblk1.cell0_I net493 net425 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_12_2891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.mux4_I\[0\].cell0_I net414 net58 net84 net110 net466 net452 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[0\].x sky130_fd_sc_hd__mux4_1
Xcol\[6\].zbuf_bot_iw_I\[1\].genblk1.cell0_I net492 col\[6\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[6\].zbuf_bot_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.tbuf_spine_ow_I\[16\].cell0_I col\[6\].genblk1.mux4_I\[16\].x net436
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[16\].z sky130_fd_sc_hd__ebufn_8
X_305_ col\[3\].zbuf_top_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[128] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_236_ col\[1\].zbuf_top_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[59] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_167_ col\[3\].zbuf_bot_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[6] sky130_fd_sc_hd__buf_2
X_098_ _030_ vssd1 vssd1 vccd1 vccd1 col\[7\].zbuf_bot_ena_I.e sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput308 um_ow[346] vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_2
Xinput319 um_ow[356] vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__dlymetal6s2s_1
Xcol\[2\].zbuf_top_iw_I\[5\].genblk1.cell0_I net483 net430 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_2920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_2839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[4\].zbuf_top_iw_I\[0\].genblk1.cell0_I net509 net426 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_219_ col\[1\].zbuf_bot_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[42] sky130_fd_sc_hd__buf_2
XFILLER_0_0_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].zbuf_top_iw_I\[16\].genblk1.cell0_I net496 net421 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_2085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[13\].genblk1.cell0_I net22 net516 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[13\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_12_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.mux4_I\[12\].cell0_I net258 net284 net310 net337 net471 net457 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[12\].x sky130_fd_sc_hd__mux4_1
Xinput127 um_ow[183] vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_1
Xinput116 um_ow[173] vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_1
Xinput105 um_ow[163] vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_1
Xcol\[7\].zbuf_bot_iw_I\[9\].genblk1.cell0_I net476 col\[7\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[7\].zbuf_bot_iw_I\[9\].z sky130_fd_sc_hd__and2_1
Xinput138 um_ow[193] vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__clkbuf_1
Xinput149 um_ow[202] vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_2737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_2472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].genblk1.tbuf_spine_ow_I\[23\].cell0_I col\[2\].genblk1.mux4_I\[23\].x net441
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[23\].z sky130_fd_sc_hd__ebufn_8
XTAP_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_2659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_2236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[0\].zbuf_bot_iw_I\[10\].genblk1.cell0_I net507 col\[0\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[0\].zbuf_bot_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[4\].genblk1.mux4_I\[3\].cell0_I net140 net167 net194 net220 net469 net456 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[3\].x sky130_fd_sc_hd__mux4_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[5\].zbuf_top_iw_I\[8\].genblk1.cell0_I net478 net424 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xzbuf_bus_iw_I\[0\].genblk1.cell0_I net8 net514 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[0\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_2681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_top_iw_I\[3\].genblk1.cell0_I net488 net420 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[3\].z sky130_fd_sc_hd__and2_1
Xcol\[2\].genblk1.tbuf_spine_ow_I\[8\].cell0_I col\[2\].genblk1.mux4_I\[8\].x net442
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z sky130_fd_sc_hd__ebufn_8
Xcol\[0\].genblk1.mux4_I\[1\].cell0_I net146 net212 net362 net389 net463 net449 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[1\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_8_2434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[0\].genblk1.mux4_I\[19\].cell0_I net145 net356 net382 net409 net461 net447 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[19\].x sky130_fd_sc_hd__mux4_2
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_2743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_2618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_2375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_398_ col\[6\].zbuf_bot_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[221] sky130_fd_sc_hd__buf_2
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtt_mux_535 vssd1 vssd1 vccd1 vccd1 tt_mux_535/HI um_k_zero[15] sky130_fd_sc_hd__conb_1
Xtt_mux_524 vssd1 vssd1 vccd1 vccd1 tt_mux_524/HI um_k_zero[4] sky130_fd_sc_hd__conb_1
XFILLER_0_8_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout422 col\[6\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_10_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout433 net434 vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout466 net467 vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__buf_4
Xfanout444 net446 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__buf_12
Xfanout455 net456 vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__clkbuf_4
Xfanout488 col\[0\].zbuf_bot_iw_I\[3\].a vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__clkbuf_4
Xfanout477 col\[0\].zbuf_bot_iw_I\[8\].a vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__buf_6
Xfanout499 col\[0\].zbuf_bot_iw_I\[14\].a vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__buf_6
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_321_ col\[4\].zbuf_bot_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[144] sky130_fd_sc_hd__buf_2
XFILLER_0_4_2673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_252_ col\[2\].zbuf_bot_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[75] sky130_fd_sc_hd__buf_2
XFILLER_0_11_2550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_2572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_183_ col\[0\].zbuf_bot_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[6] sky130_fd_sc_hd__buf_2
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].genblk1.mux4_I\[6\].cell0_I net250 net277 net304 net330 net473 net459 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[6\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_9_1861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_2183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.mux4_I\[4\].cell0_I net36 net62 net88 net115 net466 net452 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[4\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_13_2601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_304_ col\[3\].zbuf_top_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[127] sky130_fd_sc_hd__buf_2
XFILLER_0_13_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_235_ col\[1\].zbuf_top_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[58] sky130_fd_sc_hd__buf_2
XFILLER_0_11_2380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_166_ col\[2\].zbuf_top_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[5] sky130_fd_sc_hd__buf_2
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_097_ _013_ net460 _028_ vssd1 vssd1 vccd1 vccd1 _030_ sky130_fd_sc_hd__and3b_1
Xcol\[0\].genblk1.tbuf_spine_ow_I\[12\].cell0_I col\[0\].genblk1.mux4_I\[12\].x net445
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[12\].z sky130_fd_sc_hd__ebufn_8
Xtbuf_spine_ow_I\[10\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[10\].z net512 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[10\].z sky130_fd_sc_hd__ebufn_1
XFILLER_0_1_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_2234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_190 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput309 um_ow[347] vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_10_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[1\].zbuf_top_iw_I\[16\].genblk1.cell0_I net495 net431 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[16\].z sky130_fd_sc_hd__and2_1
Xcol\[0\].zbuf_bot_iw_I\[3\].genblk1.cell0_I net487 col\[0\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[0\].zbuf_bot_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_2598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_218_ col\[1\].zbuf_bot_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[41] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_149_ tbuf_spine_ow_I\[12\].z vssd1 vssd1 vccd1 vccd1 spine_ow[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_2097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.tbuf_row_ena_I.cell0_I col\[2\].genblk1.tbuf_row_ena_I.t vssd1 vssd1
+ vccd1 vccd1 col\[2\].genblk1.tbuf_row_ena_I.tx sky130_fd_sc_hd__inv_2
XFILLER_0_8_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput117 um_ow[174] vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_1
Xinput106 um_ow[164] vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_1
Xinput128 um_ow[184] vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__clkbuf_1
Xinput139 um_ow[194] vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__clkbuf_1
Xcol\[6\].genblk1.mux4_I\[16\].cell0_I net262 net288 net315 net341 net471 net457 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[16\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_90 col\[0\].genblk1.tbuf_spine_ow_I\[5\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_2605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[7\].cell0_I net144 net172 net198 net225 net468 net455 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[7\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_7_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[3\].zbuf_top_iw_I\[15\].genblk1.cell0_I net497 net427 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[3\].zbuf_bot_iw_I\[6\].genblk1.cell0_I net481 col\[3\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[3\].zbuf_bot_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[0\].genblk1.mux4_I\[5\].cell0_I net374 net256 net367 net393 net462 net448 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[5\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_6_2181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[5\].zbuf_bot_iw_I\[1\].genblk1.cell0_I net492 col\[5\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[5\].zbuf_bot_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[7\].zbuf_bot_iw_I\[17\].genblk1.cell0_I net494 col\[7\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[7\].zbuf_bot_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_2822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_397_ col\[6\].zbuf_bot_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[220] sky130_fd_sc_hd__buf_2
XFILLER_0_3_2387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[5\].zbuf_top_iw_I\[14\].genblk1.cell0_I net500 net423 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[14\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_iw_I\[5\].genblk1.cell0_I net483 net432 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[5\].z sky130_fd_sc_hd__and2_1
Xtt_mux_525 vssd1 vssd1 vccd1 vccd1 tt_mux_525/HI um_k_zero[5] sky130_fd_sc_hd__conb_1
XFILLER_0_15_2164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_2017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout423 col\[5\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__clkbuf_2
Xcol\[3\].zbuf_top_iw_I\[0\].genblk1.cell0_I net509 net428 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[0\].z sky130_fd_sc_hd__and2_1
Xfanout434 col\[0\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__clkbuf_2
Xfanout456 zbuf_bus_sel_I\[1\].z vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout445 net446 vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__buf_12
Xfanout478 col\[0\].zbuf_bot_iw_I\[8\].a vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__clkbuf_4
Xfanout489 col\[0\].zbuf_bot_iw_I\[2\].a vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_8
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout467 zbuf_bus_sel_I\[0\].z vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_2029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_320_ col\[3\].zbuf_top_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[143] sky130_fd_sc_hd__buf_2
XFILLER_0_4_2641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_251_ col\[2\].zbuf_bot_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[74] sky130_fd_sc_hd__buf_2
X_182_ col\[0\].zbuf_bot_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[5] sky130_fd_sc_hd__buf_2
XFILLER_0_11_1861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xzbuf_bus_sel_I\[2\].genblk1.cell0_I net28 net516 vssd1 vssd1 vccd1 vccd1 zbuf_bus_sel_I\[2\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_9_2563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_449_ col\[7\].zbuf_top_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[272] sky130_fd_sc_hd__buf_2
XFILLER_0_15_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[4\].genblk1.tbuf_spine_ow_I\[20\].cell0_I col\[4\].genblk1.mux4_I\[20\].x net438
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[20\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_10_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[6\].zbuf_bot_iw_I\[9\].genblk1.cell0_I net476 col\[6\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[6\].zbuf_bot_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_top_iw_I\[13\].genblk1.cell0_I net502 net419 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_2657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_2460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_303_ col\[3\].zbuf_top_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[126] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].genblk1.mux4_I\[8\].cell0_I net40 net66 net93 net119 net466 net452 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[8\].x sky130_fd_sc_hd__mux4_1
X_234_ col\[1\].zbuf_top_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[57] sky130_fd_sc_hd__buf_2
X_165_ col\[2\].zbuf_bot_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[4] sky130_fd_sc_hd__buf_2
X_096_ _029_ vssd1 vssd1 vccd1 vccd1 col\[6\].zbuf_top_ena_I.e sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[0\].genblk1.tbuf_spine_ow_I\[16\].cell0_I col\[0\].genblk1.mux4_I\[16\].x net445
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[16\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_14_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtbuf_spine_ow_I\[14\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[14\].z net511 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[14\].z sky130_fd_sc_hd__ebufn_1
XFILLER_0_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_191 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_180 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcol\[2\].genblk1.mux4_I\[11\].cell0_I net43 net70 net96 net122 net465 net451 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[11\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_2891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[4\].zbuf_top_iw_I\[8\].genblk1.cell0_I net477 net425 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].zbuf_top_iw_I\[3\].genblk1.cell0_I net488 net422 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_2408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_217_ col\[1\].zbuf_bot_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[40] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_148_ tbuf_spine_ow_I\[11\].z vssd1 vssd1 vccd1 vccd1 spine_ow[12] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_079_ _013_ _011_ _018_ vssd1 vssd1 vccd1 vccd1 _020_ sky130_fd_sc_hd__and3b_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[21\].cell0_I net161 net187 net214 net240 net469 net455 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[21\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_3_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput118 um_ow[175] vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_1
Xinput107 um_ow[165] vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_1
Xinput129 um_ow[185] vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_2785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_2605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_91 col\[0\].genblk1.tbuf_spine_ow_I\[5\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_80 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_2617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_2385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_bot_ena_I.genblk1.cell0_I net544 col\[4\].zbuf_bot_ena_I.e vssd1 vssd1
+ vccd1 vccd1 col\[4\].zbuf_bot_ena_I.z sky130_fd_sc_hd__and2_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xzbuf_bus_iw_I\[8\].genblk1.cell0_I net17 net514 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[8\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_2903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[4\].genblk1.tbuf_spine_ow_I\[0\].cell0_I col\[4\].genblk1.mux4_I\[0\].x net439
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[0\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_6_2193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[0\].genblk1.mux4_I\[9\].cell0_I net418 net301 net371 net398 net462 net448 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[9\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_14_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].zbuf_bot_iw_I\[17\].genblk1.cell0_I net493 col\[2\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[2\].zbuf_bot_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_2701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_396_ col\[6\].zbuf_bot_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[219] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_top_iw_I\[14\].genblk1.cell0_I net499 net433 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_10_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput290 um_ow[32] vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_8_2211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtt_mux_526 vssd1 vssd1 vccd1 vccd1 tt_mux_526/HI um_k_zero[6] sky130_fd_sc_hd__conb_1
XFILLER_0_8_1521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_2143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout424 col\[5\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout457 net460 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__clkbuf_4
Xfanout435 net436 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__buf_12
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout446 col\[0\].genblk1.tbuf_row_ena_I.tx vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__buf_6
Xfanout479 col\[0\].zbuf_bot_iw_I\[7\].a vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__buf_6
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout468 net469 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__buf_4
XFILLER_0_9_1307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_2839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_2653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_250_ col\[2\].zbuf_bot_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[73] sky130_fd_sc_hd__buf_2
XFILLER_0_4_2697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_181_ col\[0\].zbuf_bot_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[4] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[4\].zbuf_bot_iw_I\[16\].genblk1.cell0_I net495 col\[4\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[4\].zbuf_bot_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_2575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_2305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_448_ col\[7\].zbuf_top_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[271] sky130_fd_sc_hd__buf_2
X_379_ col\[5\].zbuf_top_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[202] sky130_fd_sc_hd__buf_2
Xzbuf_bus_iw_I\[12\].genblk1.cell1_I zbuf_bus_iw_I\[12\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[12\].a sky130_fd_sc_hd__buf_6
XFILLER_0_8_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_2826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[2\].zbuf_top_iw_I\[13\].genblk1.cell0_I net501 net429 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_302_ col\[3\].zbuf_bot_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[125] sky130_fd_sc_hd__buf_2
XFILLER_0_13_1979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_233_ col\[1\].zbuf_top_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[56] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_164_ col\[1\].zbuf_top_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[3] sky130_fd_sc_hd__buf_2
XFILLER_0_11_1681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_095_ _011_ _028_ net473 vssd1 vssd1 vccd1 vccd1 _029_ sky130_fd_sc_hd__and3b_1
XFILLER_0_9_1660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_170 net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_2113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_181 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_192 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtbuf_spine_ow_I\[18\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[18\].z net511 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[18\].z sky130_fd_sc_hd__ebufn_1
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].genblk1.mux4_I\[15\].cell0_I net48 net74 net100 net127 net464 net450 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[15\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_2809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_2645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[6\].zbuf_bot_iw_I\[15\].genblk1.cell0_I net498 col\[6\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[6\].zbuf_bot_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].zbuf_bot_iw_I\[6\].genblk1.cell0_I net481 col\[2\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[2\].zbuf_bot_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_1833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_216_ col\[1\].zbuf_bot_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[39] sky130_fd_sc_hd__buf_2
X_147_ tbuf_spine_ow_I\[10\].z vssd1 vssd1 vccd1 vccd1 spine_ow[11] sky130_fd_sc_hd__clkbuf_4
X_078_ _019_ vssd1 vssd1 vccd1 vccd1 col\[2\].zbuf_top_ena_I.e sky130_fd_sc_hd__clkbuf_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[4\].zbuf_bot_iw_I\[1\].genblk1.cell0_I net491 col\[4\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[4\].zbuf_bot_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_2309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[4\].zbuf_top_iw_I\[12\].genblk1.cell0_I net503 net425 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtbuf_row_ena_I.cell0_I net516 vssd1 vssd1 vccd1 vccd1 tbuf_row_ena_I.tx sky130_fd_sc_hd__clkinv_2
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput108 um_ow[166] vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_1
Xinput119 um_ow[176] vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_2810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_81 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_70 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_92 col\[0\].genblk1.tbuf_spine_ow_I\[5\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcol\[0\].zbuf_top_iw_I\[5\].genblk1.cell0_I net483 net434 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_2364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_2241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[2\].zbuf_top_iw_I\[0\].genblk1.cell0_I net509 net430 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput90 um_ow[14] vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_bot_ena_I.genblk1.cell0_I_550 vssd1 vssd1 vccd1 vccd1 net550 col\[7\].zbuf_bot_ena_I.genblk1.cell0_I_550/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_14_2572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[6\].zbuf_top_iw_I\[11\].genblk1.cell0_I net506 net421 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_10_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[5\].zbuf_bot_iw_I\[9\].genblk1.cell0_I net476 col\[5\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[5\].zbuf_bot_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[4\].genblk1.tbuf_spine_ow_I\[4\].cell0_I col\[4\].genblk1.mux4_I\[4\].x net440
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_2_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[7\].zbuf_bot_iw_I\[4\].genblk1.cell0_I net486 col\[7\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[7\].zbuf_bot_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[2\].genblk1.tbuf_spine_ow_I\[13\].cell0_I col\[2\].genblk1.mux4_I\[13\].x net441
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[13\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_7_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_2701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_464_ col\[7\].zbuf_top_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[287] sky130_fd_sc_hd__buf_2
XFILLER_0_10_2211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_395_ col\[6\].zbuf_bot_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[218] sky130_fd_sc_hd__buf_2
XFILLER_0_1_2080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[3\].zbuf_top_iw_I\[8\].genblk1.cell0_I net477 net427 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput280 um_ow[320] vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_1
Xinput291 um_ow[330] vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_1
Xtt_mux_527 vssd1 vssd1 vccd1 vccd1 tt_mux_527/HI um_k_zero[7] sky130_fd_sc_hd__conb_1
XFILLER_0_8_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_2267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[5\].zbuf_top_iw_I\[3\].genblk1.cell0_I net488 net424 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout436 col\[6\].genblk1.tbuf_row_ena_I.tx vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_12
Xfanout447 net449 vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__clkbuf_4
Xfanout425 col\[4\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__clkbuf_2
Xfanout458 net460 vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__clkbuf_2
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout469 net470 vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__buf_4
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_180_ col\[0\].zbuf_bot_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[3] sky130_fd_sc_hd__buf_2
XFILLER_0_11_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_2521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_2317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_447_ col\[7\].zbuf_top_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[270] sky130_fd_sc_hd__buf_2
XFILLER_0_15_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_378_ col\[5\].zbuf_top_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[201] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_301_ col\[3\].zbuf_bot_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[124] sky130_fd_sc_hd__buf_2
X_232_ col\[1\].zbuf_top_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[55] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_2350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_163_ col\[1\].zbuf_bot_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[2] sky130_fd_sc_hd__buf_2
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_094_ zbuf_bus_ena_I.z col\[6\].genblk1.tbuf_row_ena_I.t vssd1 vssd1 vccd1 vccd1
+ _028_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[0\].genblk1.mux4_I\[20\].cell0_I net157 net357 net383 net410 net461 net447 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[20\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_9_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_160 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_182 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_171 net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_193 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_2125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.mux4_I\[19\].cell0_I net52 net78 net105 net131 net464 net450 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[19\].x sky130_fd_sc_hd__mux4_1
Xcol\[1\].zbuf_bot_iw_I\[15\].genblk1.cell0_I net497 col\[1\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[1\].zbuf_bot_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_2760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_215_ col\[1\].zbuf_bot_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[38] sky130_fd_sc_hd__buf_2
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_146_ tbuf_spine_ow_I\[9\].z vssd1 vssd1 vccd1 vccd1 spine_ow[10] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_077_ _011_ _018_ _013_ vssd1 vssd1 vccd1 vccd1 _019_ sky130_fd_sc_hd__and3b_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].genblk1.tbuf_spine_ow_I\[3\].cell0_I col\[0\].genblk1.mux4_I\[3\].x net444
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[3\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput109 um_ow[167] vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_2743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_2629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtbuf_spine_ow_I\[0\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[0\].z net512 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[0\].z sky130_fd_sc_hd__ebufn_1
XANTENNA_60 col\[0\].genblk1.tbuf_spine_ow_I\[22\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_82 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_71 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_93 col\[0\].genblk1.tbuf_spine_ow_I\[5\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_2507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[3\].zbuf_bot_iw_I\[14\].genblk1.cell0_I net499 col\[3\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[3\].zbuf_bot_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_2253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput80 um_ow[140] vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput91 um_ow[150] vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[6\].genblk1.tbuf_spine_ow_I\[21\].cell0_I col\[6\].genblk1.mux4_I\[21\].x net435
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[21\].z sky130_fd_sc_hd__ebufn_8
Xcol\[1\].zbuf_top_iw_I\[11\].genblk1.cell0_I net505 net431 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_2584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xzbuf_bus_sel_I\[1\].genblk1.cell1_I zbuf_bus_sel_I\[1\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 zbuf_bus_sel_I\[1\].z sky130_fd_sc_hd__buf_6
XFILLER_0_15_2337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.tbuf_spine_ow_I\[8\].cell0_I col\[4\].genblk1.mux4_I\[8\].x net439
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_1_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].genblk1.tbuf_spine_ow_I\[17\].cell0_I col\[2\].genblk1.mux4_I\[17\].x net443
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[17\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[5\].zbuf_bot_iw_I\[13\].genblk1.cell0_I net502 col\[5\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[5\].zbuf_bot_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_2725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_463_ col\[7\].zbuf_top_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[286] sky130_fd_sc_hd__buf_2
XFILLER_0_3_2324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_394_ col\[6\].zbuf_bot_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[217] sky130_fd_sc_hd__buf_2
XFILLER_0_10_2267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput281 um_ow[321] vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__clkbuf_1
Xinput270 um_ow[311] vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_2213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput292 um_ow[331] vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_1
Xtt_mux_528 vssd1 vssd1 vccd1 vccd1 tt_mux_528/HI um_k_zero[8] sky130_fd_sc_hd__conb_1
Xtt_mux_517 vssd1 vssd1 vccd1 vccd1 tt_mux_517/HI k_zero sky130_fd_sc_hd__conb_1
XFILLER_0_15_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[3\].zbuf_top_iw_I\[10\].genblk1.cell0_I net507 net427 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout426 col\[4\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout448 net449 vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_2
Xfanout437 col\[6\].genblk1.tbuf_row_ena_I.tx vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__clkbuf_8
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout459 net460 vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_2
Xcol\[1\].zbuf_bot_iw_I\[6\].genblk1.cell0_I net481 col\[1\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[1\].zbuf_bot_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_2819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_2808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_2521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[3\].zbuf_bot_iw_I\[1\].genblk1.cell0_I net491 col\[3\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[3\].zbuf_bot_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_320 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_2121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_2165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_446_ col\[7\].zbuf_bot_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[269] sky130_fd_sc_hd__buf_2
X_377_ col\[5\].zbuf_top_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[200] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_bot_iw_I\[12\].genblk1.cell0_I net504 col\[7\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[7\].zbuf_bot_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_2863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_300_ col\[3\].zbuf_bot_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[123] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_231_ col\[1\].zbuf_top_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[54] sky130_fd_sc_hd__buf_2
XFILLER_0_13_1959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_162_ col\[0\].zbuf_top_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[1] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_2384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_093_ _027_ vssd1 vssd1 vccd1 vccd1 col\[6\].zbuf_bot_ena_I.e sky130_fd_sc_hd__buf_2
Xcol\[1\].zbuf_top_iw_I\[0\].genblk1.cell0_I net509 net432 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XANTENNA_150 col\[0\].zbuf_bot_iw_I\[6\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_2238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_161 net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_183 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_194 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_172 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_2137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_429_ col\[7\].zbuf_bot_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[252] sky130_fd_sc_hd__buf_2
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[7\].genblk1.cell1_I zbuf_bus_iw_I\[7\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[7\].a sky130_fd_sc_hd__buf_6
XFILLER_0_12_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput1 addr[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_90 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[4\].zbuf_bot_iw_I\[9\].genblk1.cell0_I net475 col\[4\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[4\].zbuf_bot_iw_I\[9\].z sky130_fd_sc_hd__and2_1
Xcol\[4\].genblk1.tbuf_spine_ow_I\[10\].cell0_I col\[4\].genblk1.mux4_I\[10\].x net439
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[10\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_6_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_2547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_214_ col\[1\].zbuf_bot_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[37] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_145_ tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 spine_ow[9] sky130_fd_sc_hd__clkbuf_4
X_076_ zbuf_bus_ena_I.z col\[2\].genblk1.tbuf_row_ena_I.t vssd1 vssd1 vccd1 vccd1
+ _018_ sky130_fd_sc_hd__and2_1
Xcol\[6\].zbuf_bot_iw_I\[4\].genblk1.cell0_I net486 col\[6\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[6\].zbuf_bot_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_2901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].genblk1.tbuf_spine_ow_I\[7\].cell0_I col\[0\].genblk1.mux4_I\[7\].x net446
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[7\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_2799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_50 col\[0\].genblk1.tbuf_spine_ow_I\[21\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_61 col\[0\].genblk1.tbuf_spine_ow_I\[22\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_72 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_83 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtbuf_spine_ow_I\[4\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[4\].z net512 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[4\].z sky130_fd_sc_hd__ebufn_2
XANTENNA_94 col\[0\].genblk1.tbuf_spine_ow_I\[5\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcol\[2\].zbuf_top_iw_I\[8\].genblk1.cell0_I net477 net429 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_15_2519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_2265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[4\].zbuf_top_iw_I\[3\].genblk1.cell0_I net487 net426 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_059_ net5 net7 vssd1 vssd1 vccd1 vccd1 _007_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_2029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput70 um_ow[131] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput81 um_ow[141] vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput92 um_ow[151] vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_2907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xzbuf_bus_iw_I\[16\].genblk1.cell0_I net25 net515 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[16\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_7_2631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_2596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_2241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[4\].genblk1.mux4_I\[11\].cell0_I net150 net176 net203 net229 net468 net454 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[11\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_15_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[0\].zbuf_bot_iw_I\[13\].genblk1.cell0_I net501 col\[0\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[0\].zbuf_bot_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_2737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_462_ col\[7\].zbuf_top_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[285] sky130_fd_sc_hd__buf_2
XFILLER_0_7_2494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_393_ col\[6\].zbuf_bot_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[216] sky130_fd_sc_hd__buf_2
XFILLER_0_14_2393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xzbuf_bus_iw_I\[3\].genblk1.cell0_I net11 net514 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[3\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput271 um_ow[312] vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_1
Xinput260 um_ow[302] vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_1
Xinput282 um_ow[322] vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__clkbuf_1
Xinput293 um_ow[332] vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_1
Xtt_mux_529 vssd1 vssd1 vccd1 vccd1 tt_mux_529/HI um_k_zero[9] sky130_fd_sc_hd__conb_1
Xtt_mux_518 vssd1 vssd1 vccd1 vccd1 tt_mux_518/HI spine_ow[0] sky130_fd_sc_hd__conb_1
XFILLER_0_8_2225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_2269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_2135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_top_iw_I\[6\].genblk1.cell0_I net482 net420 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.mux4_I\[21\].cell0_I net267 net294 net320 net347 net471 net457 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[21\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_2_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[0\].zbuf_bot_ena_I.genblk1.cell0_I net536 col\[0\].zbuf_bot_ena_I.e vssd1 vssd1
+ vccd1 vccd1 col\[0\].zbuf_bot_ena_I.z sky130_fd_sc_hd__and2_1
Xfanout427 col\[3\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__clkbuf_2
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout438 net440 vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_12
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout449 net453 vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__clkbuf_2
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_2588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_2409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_310 col\[0\].genblk1.tbuf_spine_ow_I\[1\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_321 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_2589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_445_ col\[7\].zbuf_bot_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[268] sky130_fd_sc_hd__buf_2
X_376_ col\[5\].zbuf_top_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[199] sky130_fd_sc_hd__buf_2
XFILLER_0_3_2177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[2\].zbuf_bot_iw_I\[12\].genblk1.cell0_I net503 col\[2\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[2\].zbuf_bot_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_10_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_230_ col\[1\].zbuf_bot_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[53] sky130_fd_sc_hd__buf_2
XFILLER_0_4_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_161_ col\[0\].zbuf_bot_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[0] sky130_fd_sc_hd__buf_2
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_092_ net473 net459 col\[6\].genblk1.tbuf_row_ena_I.t zbuf_bus_ena_I.z vssd1 vssd1
+ vccd1 vccd1 _027_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_0_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_151 col\[0\].zbuf_bot_iw_I\[7\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_140 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_184 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_173 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_162 net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_428_ col\[6\].zbuf_top_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[251] sky130_fd_sc_hd__buf_2
XANTENNA_195 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_2149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_2851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_359_ col\[5\].zbuf_bot_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[182] sky130_fd_sc_hd__buf_2
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput2 addr[1] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XTAP_91 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_2661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[4\].zbuf_bot_iw_I\[11\].genblk1.cell0_I net505 col\[4\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[4\].zbuf_bot_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[4\].genblk1.tbuf_spine_ow_I\[14\].cell0_I col\[4\].genblk1.mux4_I\[14\].x net438
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[14\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_4_2261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_213_ col\[1\].zbuf_bot_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[36] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_144_ tbuf_spine_ow_I\[7\].z vssd1 vssd1 vccd1 vccd1 spine_ow[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_075_ _017_ vssd1 vssd1 vccd1 vccd1 col\[2\].zbuf_bot_ena_I.e sky130_fd_sc_hd__clkbuf_4
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_2058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_2701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_2868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_40 col\[0\].genblk1.tbuf_spine_ow_I\[1\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_51 col\[0\].genblk1.tbuf_spine_ow_I\[21\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_62 col\[0\].genblk1.tbuf_spine_ow_I\[22\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_73 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_84 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_95 col\[0\].genblk1.tbuf_spine_ow_I\[5\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xtbuf_spine_ow_I\[8\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[8\].z net513 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[8\].z sky130_fd_sc_hd__ebufn_1
XFILLER_0_6_2323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_2378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_058_ net4 _004_ net1 _005_ vssd1 vssd1 vccd1 vccd1 _006_ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[0\].zbuf_bot_iw_I\[6\].genblk1.cell0_I net481 col\[0\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[0\].zbuf_bot_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_2109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_top_ena_I.genblk1.cell0_I net545 net426 vssd1 vssd1 vccd1 vccd1 col\[4\].zbuf_top_ena_I.z
+ sky130_fd_sc_hd__and2_1
Xcol\[6\].zbuf_bot_iw_I\[10\].genblk1.cell0_I net508 col\[6\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[6\].zbuf_bot_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_2798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput71 um_ow[132] vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput82 um_ow[142] vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput60 um_ow[122] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_2
Xinput93 um_ow[152] vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[2\].zbuf_bot_iw_I\[1\].genblk1.cell0_I net491 col\[2\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[2\].zbuf_bot_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_2507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_2687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_2406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].genblk1.tbuf_spine_ow_I\[21\].cell0_I col\[0\].genblk1.mux4_I\[21\].x net444
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[21\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_8_1717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_2030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[15\].cell0_I net154 net181 net207 net233 net468 net454 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[15\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_6_1485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].genblk1.tbuf_spine_ow_I\[0\].cell0_I col\[6\].genblk1.mux4_I\[0\].x net437
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[0\].z sky130_fd_sc_hd__ebufn_8
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_2873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[0\].zbuf_top_iw_I\[0\].genblk1.cell0_I net509 net434 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[0\].z sky130_fd_sc_hd__and2_1
X_461_ col\[7\].zbuf_top_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[284] sky130_fd_sc_hd__buf_2
XFILLER_0_7_2462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_392_ col\[5\].zbuf_top_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[215] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput272 um_ow[313] vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_1
Xinput250 um_ow[294] vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_1
Xinput261 um_ow[303] vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_1
Xinput283 um_ow[323] vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_1
Xinput294 um_ow[333] vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_1
Xtt_mux_519 vssd1 vssd1 vccd1 vccd1 tt_mux_519/HI spine_ow[25] sky130_fd_sc_hd__conb_1
XFILLER_0_8_2237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[3\].zbuf_bot_iw_I\[9\].genblk1.cell0_I net475 col\[3\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[3\].zbuf_bot_iw_I\[9\].z sky130_fd_sc_hd__and2_1
Xfanout428 col\[3\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout439 net440 vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__buf_12
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[5\].zbuf_bot_iw_I\[4\].genblk1.cell0_I net486 col\[5\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[5\].zbuf_bot_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_300 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_322 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_311 col\[0\].genblk1.tbuf_spine_ow_I\[1\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_444_ col\[7\].zbuf_bot_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[267] sky130_fd_sc_hd__buf_2
X_375_ col\[5\].zbuf_top_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[198] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_2808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[5\].zbuf_top_iw_I\[17\].genblk1.cell0_I net494 net423 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[17\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_iw_I\[8\].genblk1.cell0_I net477 net431 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_2410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_160_ tbuf_spine_ow_I\[23\].z vssd1 vssd1 vccd1 vccd1 spine_ow[24] sky130_fd_sc_hd__buf_4
XFILLER_0_11_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[3\].zbuf_top_iw_I\[3\].genblk1.cell0_I net487 net428 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[3\].z sky130_fd_sc_hd__and2_1
X_091_ _026_ vssd1 vssd1 vccd1 vccd1 col\[5\].zbuf_top_ena_I.e sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_2376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_152 col\[0\].zbuf_bot_iw_I\[7\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_2229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_141 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_130 col\[0\].genblk1.tbuf_spine_ow_I\[7\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_185 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_163 net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_174 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_427_ col\[6\].zbuf_top_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[250] sky130_fd_sc_hd__buf_2
XANTENNA_196 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_358_ col\[5\].zbuf_bot_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[181] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_289_ col\[3\].zbuf_bot_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[112] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput3 addr[2] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XTAP_92 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_70 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_2673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_2505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_212_ col\[0\].zbuf_top_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[35] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_2126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[4\].genblk1.tbuf_spine_ow_I\[18\].cell0_I col\[4\].genblk1.mux4_I\[18\].x net438
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[18\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_11_2183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_143_ tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 spine_ow[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_1493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_074_ net464 net450 col\[2\].genblk1.tbuf_row_ena_I.t zbuf_bus_ena_I.z vssd1 vssd1
+ vccd1 vccd1 _017_ sky130_fd_sc_hd__and4bb_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[7\].zbuf_top_iw_I\[16\].genblk1.cell0_I net496 net419 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_2015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_2757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_30 col\[0\].genblk1.tbuf_spine_ow_I\[19\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_41 col\[0\].genblk1.tbuf_spine_ow_I\[1\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_52 col\[0\].genblk1.tbuf_spine_ow_I\[21\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_63 col\[0\].genblk1.tbuf_spine_ow_I\[22\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_74 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_85 col\[0\].genblk1.tbuf_spine_ow_I\[5\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_96 col\[0\].genblk1.tbuf_spine_ow_I\[5\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[0\].genblk1.mux4_I\[10\].cell0_I net46 net312 net372 net399 net462 net448 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[10\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_15_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_2289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_2081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[6\].zbuf_top_iw_I\[6\].genblk1.cell0_I net482 net422 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[1\].zbuf_bot_iw_I\[10\].genblk1.cell0_I net507 col\[1\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[1\].zbuf_bot_iw_I\[10\].z sky130_fd_sc_hd__and2_1
X_057_ net31 vssd1 vssd1 vccd1 vccd1 _005_ sky130_fd_sc_hd__inv_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_2700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput61 um_ow[123] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_13_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput72 um_ow[133] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput50 um_ow[113] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput83 um_ow[143] vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput94 um_ow[153] vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_2633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput410 um_ow[92] vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_1
Xtbuf_spine_ow_I\[23\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[23\].z net511 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[23\].z sky130_fd_sc_hd__ebufn_1
Xcol\[2\].genblk1.mux4_I\[20\].cell0_I net53 net80 net106 net132 net464 net450 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[20\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_6_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[4\].genblk1.mux4_I\[19\].cell0_I net159 net185 net211 net238 net469 net455 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[19\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_10_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[6\].genblk1.tbuf_spine_ow_I\[4\].cell0_I col\[6\].genblk1.mux4_I\[4\].x net436
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_8_2931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_460_ col\[7\].zbuf_top_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[283] sky130_fd_sc_hd__buf_2
XFILLER_0_7_2485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_391_ col\[5\].zbuf_top_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[214] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput240 um_ow[285] vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_2
Xinput251 um_ow[295] vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_1
Xinput262 um_ow[304] vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_1
Xinput284 um_ow[324] vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_1
Xinput295 um_ow[334] vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_1
Xinput273 um_ow[314] vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_2205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_2249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.tbuf_spine_ow_I\[11\].cell0_I col\[6\].genblk1.mux4_I\[11\].x net435
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[11\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_6_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout429 col\[2\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__clkbuf_2
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_2603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_301 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_312 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_323 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_443_ col\[7\].zbuf_bot_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[266] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_374_ col\[5\].zbuf_bot_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[197] sky130_fd_sc_hd__buf_2
XFILLER_0_10_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_2056 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_2057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_top_iw_I\[17\].genblk1.cell0_I net493 net433 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_2934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_2422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_2376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_090_ _013_ _011_ _023_ vssd1 vssd1 vccd1 vccd1 _026_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_120 col\[0\].genblk1.tbuf_spine_ow_I\[7\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_131 col\[0\].genblk1.tbuf_spine_ow_I\[7\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_142 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_153 col\[0\].zbuf_bot_iw_I\[8\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_175 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_164 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_426_ col\[6\].zbuf_top_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[249] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_186 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_197 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_357_ col\[5\].zbuf_bot_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[180] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_288_ col\[3\].zbuf_bot_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[111] sky130_fd_sc_hd__buf_2
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[1\].zbuf_bot_iw_I\[1\].genblk1.cell0_I net491 col\[1\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[1\].zbuf_bot_iw_I\[1\].z sky130_fd_sc_hd__and2_1
Xinput4 addr[3] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_2906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_60 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_2720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_93 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_2641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xzbuf_bus_iw_I\[15\].genblk1.cell1_I zbuf_bus_iw_I\[15\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[15\].a sky130_fd_sc_hd__buf_6
XFILLER_0_6_2517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_211_ col\[0\].zbuf_top_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[34] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_142_ tbuf_spine_ow_I\[5\].z vssd1 vssd1 vccd1 vccd1 spine_ow[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].zbuf_top_iw_I\[16\].genblk1.cell0_I net495 net429 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[16\].z sky130_fd_sc_hd__and2_1
X_073_ _016_ vssd1 vssd1 vccd1 vccd1 col\[1\].zbuf_top_ena_I.e sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_409_ col\[6\].zbuf_bot_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[232] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.tbuf_spine_ow_I\[3\].cell0_I col\[2\].genblk1.mux4_I\[3\].x net443
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[3\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_7_2826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_2447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_31 col\[0\].genblk1.tbuf_spine_ow_I\[19\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_20 col\[0\].genblk1.tbuf_spine_ow_I\[11\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_64 col\[0\].genblk1.tbuf_spine_ow_I\[23\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 col\[0\].genblk1.tbuf_spine_ow_I\[21\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_75 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_42 col\[0\].genblk1.tbuf_spine_ow_I\[1\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_97 col\[0\].genblk1.tbuf_spine_ow_I\[5\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_86 col\[0\].genblk1.tbuf_spine_ow_I\[5\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[0\].genblk1.mux4_I\[14\].cell0_I net90 net350 net377 net403 net461 net447 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[14\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_6_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_2093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xzbuf_bus_iw_I\[2\].genblk1.cell1_I zbuf_bus_iw_I\[2\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[2\].a sky130_fd_sc_hd__buf_6
X_056_ net6 vssd1 vssd1 vccd1 vccd1 _004_ sky130_fd_sc_hd__inv_2
Xcol\[2\].zbuf_bot_iw_I\[9\].genblk1.cell0_I net475 col\[2\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[2\].zbuf_bot_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_2712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput40 um_ow[104] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput62 um_ow[124] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput73 um_ow[134] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput51 um_ow[114] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__dlymetal6s2s_1
Xcol\[4\].zbuf_bot_iw_I\[4\].genblk1.cell0_I net485 col\[4\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[4\].zbuf_bot_iw_I\[4\].z sky130_fd_sc_hd__and2_1
Xinput84 um_ow[144] vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__clkbuf_1
Xinput95 um_ow[154] vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_top_iw_I\[15\].genblk1.cell0_I net497 net425 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_2689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput400 um_ow[83] vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__clkbuf_1
Xinput411 um_ow[93] vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_2019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].zbuf_top_iw_I\[8\].genblk1.cell0_I net477 net433 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[6\].genblk1.mux4_I\[1\].cell0_I net244 net272 net298 net325 net473 net459 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[1\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_15_2820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.tbuf_spine_ow_I\[8\].cell0_I col\[6\].genblk1.mux4_I\[8\].x net437
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_2864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].zbuf_top_iw_I\[3\].genblk1.cell0_I net487 net430 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_2431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_390_ col\[5\].zbuf_top_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[213] sky130_fd_sc_hd__buf_2
XFILLER_0_3_2328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput241 um_ow[286] vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_2
Xinput230 um_ow[276] vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput252 um_ow[296] vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_1
Xinput263 um_ow[305] vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__clkbuf_1
Xinput274 um_ow[315] vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_1
Xinput285 um_ow[325] vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_1
Xinput296 um_ow[335] vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_1
Xcol\[6\].zbuf_top_iw_I\[14\].genblk1.cell0_I net500 net421 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.tbuf_spine_ow_I\[15\].cell0_I col\[6\].genblk1.mux4_I\[15\].x net436
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[15\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout419 col\[7\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__clkbuf_2
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xzbuf_bus_iw_I\[11\].genblk1.cell0_I net20 net515 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[11\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_2773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_2659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_bot_iw_I\[7\].genblk1.cell0_I net480 col\[7\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[7\].zbuf_bot_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_302 col\[0\].genblk1.tbuf_spine_ow_I\[1\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_324 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_313 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_442_ col\[7\].zbuf_bot_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[265] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_373_ col\[5\].zbuf_bot_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[196] sky130_fd_sc_hd__buf_2
XFILLER_0_7_1593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_2434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[5\].zbuf_top_iw_I\[6\].genblk1.cell0_I net482 net424 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_2309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].genblk1.mux4_I\[11\].cell0_I net255 net283 net309 net336 net471 net458 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[11\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_5_2209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_132 col\[0\].genblk1.tbuf_spine_ow_I\[7\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_121 col\[0\].genblk1.tbuf_spine_ow_I\[7\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_143 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_110 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_154 col\[0\].zbuf_bot_iw_I\[8\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcol\[7\].zbuf_top_iw_I\[1\].genblk1.cell0_I net492 net420 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XANTENNA_165 net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_176 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_425_ col\[6\].zbuf_top_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[248] sky130_fd_sc_hd__buf_2
XANTENNA_187 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_198 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_356_ col\[4\].zbuf_top_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[179] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_287_ col\[3\].zbuf_bot_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[110] sky130_fd_sc_hd__buf_2
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.tbuf_spine_ow_I\[22\].cell0_I col\[2\].genblk1.mux4_I\[22\].x net441
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[22\].z sky130_fd_sc_hd__ebufn_8
Xinput5 addr[4] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XTAP_50 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_94 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_2743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_2529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[2\].cell0_I net139 net166 net193 net219 net470 net456 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[2\].x sky130_fd_sc_hd__mux4_1
X_210_ col\[0\].zbuf_top_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[33] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_2141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_141_ tbuf_spine_ow_I\[4\].z vssd1 vssd1 vccd1 vccd1 spine_ow[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_072_ _013_ _011_ _012_ vssd1 vssd1 vccd1 vccd1 _016_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_2153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_408_ col\[6\].zbuf_bot_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[231] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_339_ col\[4\].zbuf_top_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[162] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.tbuf_spine_ow_I\[7\].cell0_I col\[2\].genblk1.mux4_I\[7\].x net442
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[7\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_12_2461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].genblk1.mux4_I\[0\].cell0_I net35 net201 net361 net388 net463 net449 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[0\].x sky130_fd_sc_hd__mux4_2
XANTENNA_32 col\[0\].genblk1.tbuf_spine_ow_I\[19\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 col\[0\].genblk1.tbuf_spine_ow_I\[0\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 col\[0\].genblk1.tbuf_spine_ow_I\[11\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_54 col\[0\].genblk1.tbuf_spine_ow_I\[22\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_65 col\[0\].genblk1.tbuf_spine_ow_I\[23\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_43 col\[0\].genblk1.tbuf_spine_ow_I\[1\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_98 col\[0\].genblk1.tbuf_spine_ow_I\[5\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_87 col\[0\].genblk1.tbuf_spine_ow_I\[5\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_76 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcol\[0\].genblk1.mux4_I\[18\].cell0_I net134 net355 net381 net408 net461 net447 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[18\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_6_2348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_055_ _001_ _002_ vssd1 vssd1 vccd1 vccd1 _003_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput30 spine_iw[5] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput63 um_ow[125] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_0_1780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput41 um_ow[105] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput52 um_ow[115] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput74 um_ow[135] vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_13_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput85 um_ow[145] vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_1
Xinput96 um_ow[155] vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput401 um_ow[84] vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__clkbuf_1
Xinput412 um_ow[94] vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_2101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[3\].zbuf_bot_iw_I\[17\].genblk1.cell0_I net493 col\[3\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[3\].zbuf_bot_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[6\].genblk1.mux4_I\[5\].cell0_I net249 net276 net303 net329 net473 net459 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[5\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_15_2854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[0\].zbuf_bot_iw_I\[1\].genblk1.cell0_I net491 col\[0\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[0\].zbuf_bot_iw_I\[1\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_iw_I\[14\].genblk1.cell0_I net499 net431 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[14\].z sky130_fd_sc_hd__and2_1
Xinput220 um_ow[267] vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput242 um_ow[287] vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_2
Xinput231 um_ow[277] vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput253 um_ow[297] vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_1
Xinput275 um_ow[316] vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_1
Xinput286 um_ow[326] vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_1
Xinput297 um_ow[336] vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput264 um_ow[306] vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[2\].genblk1.mux4_I\[3\].cell0_I net417 net61 net87 net114 net466 net452 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[3\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_sel_I\[4\].genblk1.cell1_I zbuf_bus_sel_I\[4\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 zbuf_bus_sel_I\[4\].z sky130_fd_sc_hd__buf_6
XFILLER_0_14_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[6\].genblk1.tbuf_spine_ow_I\[19\].cell0_I col\[6\].genblk1.mux4_I\[19\].x net435
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[19\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_10_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[0\].genblk1.tbuf_spine_ow_I\[11\].cell0_I col\[0\].genblk1.mux4_I\[11\].x net445
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[11\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_8_2741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_top_ena_I.genblk1.cell0_I net537 net434 vssd1 vssd1 vccd1 vccd1 col\[0\].zbuf_top_ena_I.z
+ sky130_fd_sc_hd__and2_1
XFILLER_0_8_2785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_303 col\[0\].genblk1.tbuf_spine_ow_I\[1\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_314 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_325 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_441_ col\[7\].zbuf_bot_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[264] sky130_fd_sc_hd__buf_2
X_372_ col\[5\].zbuf_bot_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[195] sky130_fd_sc_hd__buf_2
XFILLER_0_7_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_2295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[5\].zbuf_bot_iw_I\[16\].genblk1.cell0_I net496 col\[5\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[5\].zbuf_bot_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[3\].zbuf_top_iw_I\[13\].genblk1.cell0_I net501 net427 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[1\].zbuf_bot_iw_I\[9\].genblk1.cell0_I net475 col\[1\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[1\].zbuf_bot_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XANTENNA_100 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[6\].genblk1.mux4_I\[15\].cell0_I net261 net287 net314 net340 net472 net458 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[15\].x sky130_fd_sc_hd__mux4_1
XANTENNA_133 col\[0\].genblk1.tbuf_spine_ow_I\[7\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_122 col\[0\].genblk1.tbuf_spine_ow_I\[7\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_111 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_424_ col\[6\].zbuf_top_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[247] sky130_fd_sc_hd__buf_2
XANTENNA_155 col\[0\].zbuf_bot_iw_I\[9\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_166 net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_144 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_177 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_199 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_188 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_355_ col\[4\].zbuf_top_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[178] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_2855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_286_ col\[3\].zbuf_bot_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[109] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[3\].zbuf_bot_iw_I\[4\].genblk1.cell0_I net485 col\[3\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[3\].zbuf_bot_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput6 spine_iw[10] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XTAP_40 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_51 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_84 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_95 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[7\].zbuf_bot_iw_I\[15\].genblk1.cell0_I net498 col\[7\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[7\].zbuf_bot_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_2210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_2129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_2107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[4\].genblk1.mux4_I\[6\].cell0_I net143 net171 net197 net224 net470 net456 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[6\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_140_ tbuf_spine_ow_I\[3\].z vssd1 vssd1 vccd1 vccd1 spine_ow[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_2197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_071_ _015_ vssd1 vssd1 vccd1 vccd1 col\[1\].zbuf_bot_ena_I.e sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_2121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_2165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_2917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_407_ col\[6\].zbuf_bot_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[230] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_338_ col\[4\].zbuf_bot_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[161] sky130_fd_sc_hd__buf_2
Xcol\[5\].zbuf_top_iw_I\[12\].genblk1.cell0_I net504 net423 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[12\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_iw_I\[3\].genblk1.cell0_I net487 net432 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_269_ col\[2\].zbuf_top_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[92] sky130_fd_sc_hd__buf_2
XFILLER_0_4_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_2574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_2473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_11 col\[0\].genblk1.tbuf_spine_ow_I\[0\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 col\[0\].genblk1.tbuf_spine_ow_I\[11\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_55 col\[0\].genblk1.tbuf_spine_ow_I\[22\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_44 col\[0\].genblk1.tbuf_spine_ow_I\[21\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_66 col\[0\].genblk1.tbuf_spine_ow_I\[23\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcol\[0\].genblk1.mux4_I\[4\].cell0_I net363 net245 net366 net392 net463 net449 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[4\].x sky130_fd_sc_hd__mux4_2
XANTENNA_33 col\[0\].genblk1.tbuf_spine_ow_I\[19\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_88 col\[0\].genblk1.tbuf_spine_ow_I\[5\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_99 col\[0\].genblk1.tbuf_spine_ow_I\[5\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_77 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xzbuf_bus_sel_I\[0\].genblk1.cell0_I net32 net516 vssd1 vssd1 vccd1 vccd1 zbuf_bus_sel_I\[0\].genblk1.l
+ sky130_fd_sc_hd__and2_1
X_054_ net3 net34 vssd1 vssd1 vccd1 vccd1 _002_ sky130_fd_sc_hd__xor2_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xzbuf_bus_ena_I.genblk1.cell1_I zbuf_bus_ena_I.genblk1.l vssd1 vssd1 vccd1 vccd1 zbuf_bus_ena_I.z
+ sky130_fd_sc_hd__buf_8
XFILLER_0_6_2850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[6\].zbuf_bot_iw_I\[7\].genblk1.cell0_I net480 col\[6\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[6\].zbuf_bot_iw_I\[7\].z sky130_fd_sc_hd__and2_1
Xinput31 spine_iw[6] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput20 spine_iw[23] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput64 um_ow[126] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput42 um_ow[106] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput53 um_ow[116] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_4_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput75 um_ow[136] vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput86 um_ow[146] vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_1
Xinput97 um_ow[156] vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_2669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_2224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput402 um_ow[85] vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__clkbuf_1
Xcol\[7\].zbuf_top_iw_I\[11\].genblk1.cell0_I net506 net419 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[11\].z sky130_fd_sc_hd__and2_1
Xinput413 um_ow[95] vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_2113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[5\].zbuf_bot_ena_I.genblk1.cell0_I net546 col\[5\].zbuf_bot_ena_I.e vssd1 vssd1
+ vccd1 vccd1 col\[5\].zbuf_bot_ena_I.z sky130_fd_sc_hd__and2_1
XFILLER_0_11_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[4\].zbuf_top_iw_I\[6\].genblk1.cell0_I net481 net426 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_2544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.mux4_I\[9\].cell0_I net253 net281 net307 net333 net472 net458 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[9\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_2_2599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[6\].zbuf_top_iw_I\[1\].genblk1.cell0_I net492 net422 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_1620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput210 um_ow[258] vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput232 um_ow[278] vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput221 um_ow[268] vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput254 um_ow[298] vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_1
Xinput243 um_ow[288] vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_1
Xinput276 um_ow[317] vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_1
Xinput287 um_ow[327] vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_1
Xinput265 um_ow[307] vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_1
Xinput298 um_ow[337] vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_15_2129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_2853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_2741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.mux4_I\[7\].cell0_I net39 net65 net92 net118 net466 net452 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[7\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_10_2785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].genblk1.tbuf_spine_ow_I\[15\].cell0_I col\[0\].genblk1.mux4_I\[15\].x net446
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[15\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_4_2617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtbuf_spine_ow_I\[13\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[13\].z net511 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[13\].z sky130_fd_sc_hd__ebufn_1
XFILLER_0_5_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[2\].genblk1.mux4_I\[10\].cell0_I net42 net69 net95 net121 net464 net450 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[10\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_13_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].zbuf_bot_iw_I\[16\].genblk1.cell0_I net495 col\[0\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[0\].zbuf_bot_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_304 col\[0\].genblk1.tbuf_spine_ow_I\[1\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_2241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_315 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_440_ col\[7\].zbuf_bot_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[263] sky130_fd_sc_hd__buf_2
XANTENNA_326 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_2151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_371_ col\[5\].zbuf_bot_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[194] sky130_fd_sc_hd__buf_2
XFILLER_0_3_2127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_2037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_2847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xzbuf_bus_iw_I\[6\].genblk1.cell0_I net14 net514 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[6\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_10_2593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[7\].zbuf_top_iw_I\[9\].genblk1.cell0_I net476 net419 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[20\].cell0_I net160 net186 net213 net239 net469 net455 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[20\].x sky130_fd_sc_hd__mux4_1
XANTENNA_101 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_123 col\[0\].genblk1.tbuf_spine_ow_I\[7\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_134 col\[0\].genblk1.tbuf_spine_ow_I\[7\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_112 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_156 col\[0\].zbuf_bot_iw_I\[9\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_423_ col\[6\].zbuf_top_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[246] sky130_fd_sc_hd__buf_2
XANTENNA_145 col\[0\].zbuf_bot_iw_I\[10\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_2071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_167 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_189 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_178 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_354_ col\[4\].zbuf_top_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[177] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].genblk1.mux4_I\[19\].cell0_I net265 net292 net318 net344 net471 net457 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[19\].x sky130_fd_sc_hd__mux4_1
X_285_ col\[3\].zbuf_bot_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[108] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput7 spine_iw[11] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XTAP_41 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_2701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_85 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[2\].zbuf_bot_iw_I\[15\].genblk1.cell0_I net497 col\[2\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[2\].zbuf_bot_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XTAP_63 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_52 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_2609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_96 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_070_ _013_ _011_ _012_ vssd1 vssd1 vccd1 vccd1 _015_ sky130_fd_sc_hd__and3b_1
XFILLER_0_14_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].zbuf_top_iw_I\[12\].genblk1.cell0_I net503 net433 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_1421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_2920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_406_ col\[6\].zbuf_bot_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[229] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_337_ col\[4\].zbuf_bot_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[160] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_268_ col\[2\].zbuf_top_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[91] sky130_fd_sc_hd__buf_2
X_199_ col\[0\].zbuf_top_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[22] sky130_fd_sc_hd__buf_2
XFILLER_0_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_2597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_2485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_12 col\[0\].genblk1.tbuf_spine_ow_I\[0\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 col\[0\].genblk1.tbuf_spine_ow_I\[11\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_45 col\[0\].genblk1.tbuf_spine_ow_I\[21\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_56 col\[0\].genblk1.tbuf_spine_ow_I\[22\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 col\[0\].genblk1.tbuf_spine_ow_I\[19\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_89 col\[0\].genblk1.tbuf_spine_ow_I\[5\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_67 col\[0\].genblk1.tbuf_spine_ow_I\[23\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_78 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[0\].genblk1.mux4_I\[8\].cell0_I net407 net290 net370 net397 net462 net448 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[8\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_3_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_053_ net2 net33 vssd1 vssd1 vccd1 vccd1 _001_ sky130_fd_sc_hd__xor2_1
Xcol\[4\].zbuf_bot_iw_I\[14\].genblk1.cell0_I net499 col\[4\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[4\].zbuf_bot_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_2873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput21 spine_iw[24] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
Xinput10 spine_iw[14] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput32 spine_iw[7] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput54 um_ow[117] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_0_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput43 um_ow[107] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput65 um_ow[127] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput76 um_ow[137] vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput87 um_ow[147] vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_1
Xinput98 um_ow[157] vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[10\].genblk1.cell1_I zbuf_bus_iw_I\[10\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[10\].a sky130_fd_sc_hd__buf_6
XFILLER_0_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].zbuf_top_iw_I\[11\].genblk1.cell0_I net505 net429 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_2236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput403 um_ow[86] vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__clkbuf_1
Xinput414 um_ow[96] vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_6_2125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_bot_iw_I\[9\].genblk1.cell0_I net475 col\[0\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[0\].zbuf_bot_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[6\].zbuf_bot_iw_I\[13\].genblk1.cell0_I net502 col\[6\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[6\].zbuf_bot_iw_I\[13\].z sky130_fd_sc_hd__and2_1
Xcol\[4\].genblk1.tbuf_spine_ow_I\[23\].cell0_I col\[4\].genblk1.mux4_I\[23\].x net438
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[23\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_14_2322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_2066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[2\].zbuf_bot_iw_I\[4\].genblk1.cell0_I net485 col\[2\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[2\].zbuf_bot_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput200 um_ow[249] vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput211 um_ow[259] vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput222 um_ow[269] vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput233 um_ow[279] vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput244 um_ow[289] vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_1
Xinput277 um_ow[318] vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_1
Xinput288 um_ow[328] vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_1
Xinput255 um_ow[299] vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_1
Xinput266 um_ow[308] vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_1
Xinput299 um_ow[338] vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_15_2108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_2753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[4\].zbuf_top_iw_I\[10\].genblk1.cell0_I net507 net425 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_10_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_2765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_2620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_2386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[0\].genblk1.tbuf_spine_ow_I\[19\].cell0_I col\[0\].genblk1.mux4_I\[19\].x net446
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[19\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_11_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtbuf_spine_ow_I\[17\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[17\].z net511 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[17\].z sky130_fd_sc_hd__ebufn_1
XFILLER_0_1_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[2\].genblk1.mux4_I\[14\].cell0_I net47 net73 net99 net126 net464 net451 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[14\].x sky130_fd_sc_hd__mux4_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_305 col\[0\].genblk1.tbuf_spine_ow_I\[1\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_316 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_327 zbuf_bus_ena_I.z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_2253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_370_ col\[5\].zbuf_bot_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[193] sky130_fd_sc_hd__buf_2
XFILLER_0_7_2297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_top_iw_I\[3\].genblk1.cell0_I net487 net434 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_2927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_102 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_124 col\[0\].genblk1.tbuf_spine_ow_I\[7\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_113 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_146 col\[0\].zbuf_bot_iw_I\[2\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_422_ col\[6\].zbuf_top_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[245] sky130_fd_sc_hd__buf_2
XANTENNA_135 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_157 zbuf_bus_ena_I.z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_168 net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_179 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_353_ col\[4\].zbuf_top_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[176] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[5\].zbuf_bot_iw_I\[7\].genblk1.cell0_I net480 col\[5\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[5\].zbuf_bot_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_284_ col\[2\].zbuf_top_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[107] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 spine_iw[12] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XTAP_42 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_2713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_2601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_75 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_53 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_2724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[7\].zbuf_bot_iw_I\[2\].genblk1.cell0_I net490 col\[7\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[7\].zbuf_bot_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XTAP_97 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_2177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_2009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[3\].zbuf_top_iw_I\[6\].genblk1.cell0_I net481 net428 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_2910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_405_ col\[6\].zbuf_bot_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[228] sky130_fd_sc_hd__buf_2
X_336_ col\[4\].zbuf_bot_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[159] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_267_ col\[2\].zbuf_top_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[90] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_198_ col\[0\].zbuf_top_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[21] sky130_fd_sc_hd__buf_2
Xcol\[5\].zbuf_top_iw_I\[1\].genblk1.cell0_I net492 net424 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_2521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_13 col\[0\].genblk1.tbuf_spine_ow_I\[11\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_46 col\[0\].genblk1.tbuf_spine_ow_I\[21\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 col\[0\].genblk1.tbuf_spine_ow_I\[19\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_57 col\[0\].genblk1.tbuf_spine_ow_I\[22\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_24 col\[0\].genblk1.tbuf_spine_ow_I\[11\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_68 col\[0\].genblk1.tbuf_spine_ow_I\[23\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_79 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.tbuf_spine_ow_I\[3\].cell0_I col\[4\].genblk1.mux4_I\[3\].x net440
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[3\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.tbuf_spine_ow_I\[12\].cell0_I col\[2\].genblk1.mux4_I\[12\].x net443
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[12\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_13_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_052_ _000_ vssd1 vssd1 vccd1 vccd1 col\[6\].genblk1.tbuf_row_ena_I.t sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_2863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_319_ col\[3\].zbuf_top_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[142] sky130_fd_sc_hd__buf_2
Xinput22 spine_iw[25] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
Xinput11 spine_iw[15] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
Xinput44 um_ow[108] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_0_1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput55 um_ow[118] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput33 spine_iw[8] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
Xinput66 um_ow[128] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput77 um_ow[138] vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput88 um_ow[148] vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput99 um_ow[158] vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_2261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput404 um_ow[87] vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__clkbuf_1
Xinput415 um_ow[97] vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_6_2137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_2924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[2\].zbuf_bot_ena_I.genblk1.cell0_I_540 vssd1 vssd1 vccd1 vccd1 net540 col\[2\].zbuf_bot_ena_I.genblk1.cell0_I_540/LO
+ sky130_fd_sc_hd__conb_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[6\].zbuf_top_iw_I\[9\].genblk1.cell0_I net476 net421 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_15_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[1\].zbuf_bot_iw_I\[13\].genblk1.cell0_I net501 col\[1\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[1\].zbuf_bot_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_1845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_2435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_2089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput201 um_ow[24] vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_2
Xinput212 um_ow[25] vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__clkbuf_2
Xinput245 um_ow[28] vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_2
Xinput234 um_ow[27] vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_2
Xinput223 um_ow[26] vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_2
Xinput278 um_ow[319] vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_1
Xinput256 um_ow[29] vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_2
Xinput267 um_ow[309] vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_1
Xinput289 um_ow[329] vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_1509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[2\].genblk1.mux4_I\[18\].cell0_I net51 net77 net104 net130 net464 net450 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[18\].x sky130_fd_sc_hd__mux4_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_306 col\[0\].genblk1.tbuf_spine_ow_I\[1\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_317 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_2265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_328 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_2142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[3\].zbuf_bot_iw_I\[12\].genblk1.cell0_I net503 col\[3\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[3\].zbuf_bot_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_2805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[3\].zbuf_bot_ena_I.genblk1.cell0_I_542 vssd1 vssd1 vccd1 vccd1 net542 col\[3\].zbuf_bot_ena_I.genblk1.cell0_I_542/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_10_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_2405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].genblk1.tbuf_spine_ow_I\[2\].cell0_I col\[0\].genblk1.mux4_I\[2\].x net444
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[2\].z sky130_fd_sc_hd__ebufn_8
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_103 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_125 col\[0\].genblk1.tbuf_spine_ow_I\[7\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_114 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_147 col\[0\].zbuf_bot_iw_I\[5\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_421_ col\[6\].zbuf_top_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[244] sky130_fd_sc_hd__buf_2
XANTENNA_136 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_2073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_158 zbuf_bus_ena_I.z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_352_ col\[4\].zbuf_top_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[175] sky130_fd_sc_hd__buf_2
XANTENNA_169 net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_283_ col\[2\].zbuf_top_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[106] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput9 spine_iw[13] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XTAP_32 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_76 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_43 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_54 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_98 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_2769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[5\].zbuf_bot_iw_I\[11\].genblk1.cell0_I net506 col\[5\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[5\].zbuf_bot_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.tbuf_spine_ow_I\[20\].cell0_I col\[6\].genblk1.mux4_I\[20\].x net435
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[20\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_9_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_404_ col\[6\].zbuf_bot_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[227] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_335_ col\[4\].zbuf_bot_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[158] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_266_ col\[2\].zbuf_bot_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[89] sky130_fd_sc_hd__buf_2
X_197_ col\[0\].zbuf_top_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[20] sky130_fd_sc_hd__buf_2
XFILLER_0_5_2533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_2577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_14 col\[0\].genblk1.tbuf_spine_ow_I\[11\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_47 col\[0\].genblk1.tbuf_spine_ow_I\[21\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_36 col\[0\].genblk1.tbuf_spine_ow_I\[19\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 col\[0\].genblk1.tbuf_spine_ow_I\[11\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[1\].zbuf_bot_iw_I\[4\].genblk1.cell0_I net485 col\[1\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[1\].zbuf_bot_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XANTENNA_58 col\[0\].genblk1.tbuf_spine_ow_I\[22\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_69 col\[0\].genblk1.tbuf_spine_ow_I\[4\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.tbuf_spine_ow_I\[7\].cell0_I col\[4\].genblk1.mux4_I\[7\].x net439
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[7\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_11_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_bot_ena_I.genblk1.cell0_I_544 vssd1 vssd1 vccd1 vccd1 net544 col\[4\].zbuf_bot_ena_I.genblk1.cell0_I_544/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_2043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[2\].genblk1.tbuf_spine_ow_I\[16\].cell0_I col\[2\].genblk1.mux4_I\[16\].x net441
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[16\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_4_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_051_ zbuf_bus_sel_I\[4\].z zbuf_bus_sel_I\[2\].z zbuf_bus_sel_I\[3\].z vssd1 vssd1
+ vccd1 vccd1 _000_ sky130_fd_sc_hd__and3b_1
XFILLER_0_2_2717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_318_ col\[3\].zbuf_top_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[141] sky130_fd_sc_hd__buf_2
Xcol\[7\].zbuf_bot_iw_I\[10\].genblk1.cell0_I net508 col\[7\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[7\].zbuf_bot_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_2463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 spine_iw[16] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_249_ col\[2\].zbuf_bot_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[72] sky130_fd_sc_hd__buf_2
Xinput45 um_ow[109] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput23 spine_iw[26] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 spine_iw[9] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
Xinput78 um_ow[139] vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput67 um_ow[129] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput89 um_ow[149] vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_1
Xinput56 um_ow[119] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput405 um_ow[88] vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__clkbuf_1
Xinput416 um_ow[98] vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_6_2149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_2836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[5\].genblk1.cell1_I zbuf_bus_iw_I\[5\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[5\].a sky130_fd_sc_hd__buf_6
XFILLER_0_0_2260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_2302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_bot_iw_I\[7\].genblk1.cell0_I net479 col\[4\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[4\].zbuf_bot_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_2057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput202 um_ow[250] vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__clkbuf_2
Xinput224 um_ow[270] vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput235 um_ow[280] vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_2
Xinput213 um_ow[260] vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__dlymetal6s2s_1
Xcol\[5\].zbuf_bot_ena_I.genblk1.cell0_I_546 vssd1 vssd1 vccd1 vccd1 net546 col\[5\].zbuf_bot_ena_I.genblk1.cell0_I_546/LO
+ sky130_fd_sc_hd__conb_1
Xinput268 um_ow[30] vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_2
Xinput279 um_ow[31] vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_2
Xinput246 um_ow[290] vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_1
Xinput257 um_ow[2] vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[6\].zbuf_bot_iw_I\[2\].genblk1.cell0_I net490 col\[6\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[6\].zbuf_bot_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_2344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].genblk1.mux4_I\[23\].cell0_I net190 net360 net387 net413 net461 net447 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[23\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_307 col\[0\].genblk1.tbuf_spine_ow_I\[1\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_2233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_318 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_329 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcol\[2\].zbuf_top_iw_I\[6\].genblk1.cell0_I net481 net430 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_2277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_top_iw_I\[1\].genblk1.cell0_I net491 net426 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_2631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[1\].zbuf_bot_ena_I.genblk1.cell0_I net538 col\[1\].zbuf_bot_ena_I.e vssd1 vssd1
+ vccd1 vccd1 col\[1\].zbuf_bot_ena_I.z sky130_fd_sc_hd__and2_1
XFILLER_0_1_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].zbuf_top_iw_I\[17\].genblk1.cell0_I net494 net421 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_2463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[14\].genblk1.cell0_I net23 net516 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[14\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].genblk1.tbuf_spine_ow_I\[6\].cell0_I col\[0\].genblk1.mux4_I\[6\].x net446
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z sky130_fd_sc_hd__ebufn_8
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_115 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_420_ col\[6\].zbuf_top_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[243] sky130_fd_sc_hd__buf_2
XANTENNA_148 col\[0\].zbuf_bot_iw_I\[5\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_137 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_126 col\[0\].genblk1.tbuf_spine_ow_I\[7\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_351_ col\[4\].zbuf_top_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[174] sky130_fd_sc_hd__buf_2
XFILLER_0_7_2085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_159 zbuf_bus_ena_I.z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_282_ col\[2\].zbuf_top_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[105] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtbuf_spine_ow_I\[3\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[3\].z net512 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[3\].z sky130_fd_sc_hd__ebufn_1
Xcol\[6\].zbuf_bot_ena_I.genblk1.cell0_I_548 vssd1 vssd1 vccd1 vccd1 net548 col\[6\].zbuf_bot_ena_I.genblk1.cell0_I_548/LO
+ sky130_fd_sc_hd__conb_1
XTAP_33 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_44 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_99 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_bot_iw_I\[11\].genblk1.cell0_I net505 col\[0\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[0\].zbuf_bot_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_2350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_2236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[5\].zbuf_top_iw_I\[9\].genblk1.cell0_I net476 net423 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_403_ col\[6\].zbuf_bot_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[226] sky130_fd_sc_hd__buf_2
XFILLER_0_13_2934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xzbuf_bus_iw_I\[1\].genblk1.cell0_I net9 net514 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[1\].genblk1.l
+ sky130_fd_sc_hd__and2_1
X_334_ col\[4\].zbuf_bot_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[157] sky130_fd_sc_hd__buf_2
X_265_ col\[2\].zbuf_bot_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[88] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_196_ col\[0\].zbuf_top_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[19] sky130_fd_sc_hd__buf_2
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_top_iw_I\[4\].genblk1.cell0_I net486 net420 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_2545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_48 col\[0\].genblk1.tbuf_spine_ow_I\[21\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 col\[0\].genblk1.tbuf_spine_ow_I\[19\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 col\[0\].genblk1.tbuf_spine_ow_I\[11\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_15 col\[0\].genblk1.tbuf_spine_ow_I\[11\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcol\[4\].genblk1.mux4_I\[10\].cell0_I net149 net175 net202 net228 net468 net454 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[10\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_12_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_59 col\[0\].genblk1.tbuf_spine_ow_I\[22\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_050_ zbuf_bus_sel_I\[4\].z zbuf_bus_sel_I\[2\].z zbuf_bus_sel_I\[3\].z vssd1 vssd1
+ vccd1 vccd1 col\[4\].genblk1.tbuf_row_ena_I.t sky130_fd_sc_hd__nor3b_2
XFILLER_0_15_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].zbuf_bot_iw_I\[10\].genblk1.cell0_I net507 col\[2\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[2\].zbuf_bot_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_2720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_2898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_317_ col\[3\].zbuf_top_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[140] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput13 spine_iw[17] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
X_248_ col\[1\].zbuf_top_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[71] sky130_fd_sc_hd__buf_2
Xinput35 um_ow[0] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_2
Xinput46 um_ow[10] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput24 spine_iw[27] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
Xinput68 um_ow[12] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_2
Xinput57 um_ow[11] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_2
Xinput79 um_ow[13] vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_2
X_179_ col\[0\].zbuf_bot_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[2] sky130_fd_sc_hd__buf_2
XFILLER_0_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[6\].genblk1.mux4_I\[20\].cell0_I net266 net293 net319 net346 net471 net457 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[20\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_11_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput406 um_ow[89] vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__clkbuf_1
Xinput417 um_ow[99] vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_6_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_2740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[5\].zbuf_top_ena_I.genblk1.cell0_I net547 net423 vssd1 vssd1 vccd1 vccd1 col\[5\].zbuf_top_ena_I.z
+ sky130_fd_sc_hd__and2_1
XFILLER_0_15_2826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_2325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_2358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput225 um_ow[271] vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput236 um_ow[281] vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__clkbuf_2
Xinput203 um_ow[251] vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__clkbuf_2
Xinput214 um_ow[261] vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput247 um_ow[291] vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_1
Xinput258 um_ow[300] vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_1
Xinput269 um_ow[310] vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_2857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_2645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_308 col\[0\].genblk1.tbuf_spine_ow_I\[1\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_319 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_2109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[0\].zbuf_bot_iw_I\[4\].genblk1.cell0_I net485 col\[0\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[0\].zbuf_bot_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_1953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[1\].zbuf_top_iw_I\[17\].genblk1.cell0_I net493 net431 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[4\].genblk1.tbuf_spine_ow_I\[13\].cell0_I col\[4\].genblk1.mux4_I\[13\].x net439
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[13\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_3_1997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_116 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_149 col\[0\].zbuf_bot_iw_I\[6\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_138 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_127 col\[0\].genblk1.tbuf_spine_ow_I\[7\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_2097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_350_ col\[4\].zbuf_top_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[173] sky130_fd_sc_hd__buf_2
X_281_ col\[2\].zbuf_top_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[104] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtbuf_spine_ow_I\[7\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[7\].z net513 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[7\].z sky130_fd_sc_hd__ebufn_1
XTAP_67 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_34 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_45 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_2716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_89 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_2495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[7\].zbuf_top_ena_I.genblk1.cell0_I_551 vssd1 vssd1 vccd1 vccd1 net551 col\[7\].zbuf_top_ena_I.genblk1.cell0_I_551/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[3\].zbuf_top_iw_I\[16\].genblk1.cell0_I net495 net427 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_402_ col\[6\].zbuf_bot_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[225] sky130_fd_sc_hd__buf_2
XFILLER_0_9_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_333_ col\[4\].zbuf_bot_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[156] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_264_ col\[2\].zbuf_bot_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[87] sky130_fd_sc_hd__buf_2
XFILLER_0_11_2681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_195_ col\[0\].zbuf_top_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[18] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].genblk1.tbuf_spine_ow_I\[20\].cell0_I col\[0\].genblk1.mux4_I\[20\].x net444
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[20\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[3\].zbuf_bot_iw_I\[7\].genblk1.cell0_I net479 col\[3\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[3\].zbuf_bot_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_38 col\[0\].genblk1.tbuf_spine_ow_I\[19\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_2292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_27 col\[0\].genblk1.tbuf_spine_ow_I\[11\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_16 col\[0\].genblk1.tbuf_spine_ow_I\[11\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_49 col\[0\].genblk1.tbuf_spine_ow_I\[21\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[14\].cell0_I net153 net180 net206 net232 net468 net454 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[14\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[5\].zbuf_bot_iw_I\[2\].genblk1.cell0_I net490 col\[5\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[5\].zbuf_bot_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_2001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_316_ col\[3\].zbuf_top_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[139] sky130_fd_sc_hd__buf_2
XFILLER_0_13_2776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_247_ col\[1\].zbuf_top_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[70] sky130_fd_sc_hd__buf_2
Xinput36 um_ow[100] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput25 spine_iw[28] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
Xinput14 spine_iw[18] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
Xinput58 um_ow[120] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput69 um_ow[130] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput47 um_ow[110] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dlymetal6s2s_1
X_178_ col\[0\].zbuf_bot_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[1] sky130_fd_sc_hd__buf_2
XFILLER_0_0_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[1\].zbuf_top_iw_I\[6\].genblk1.cell0_I net481 net432 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_1929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[5\].zbuf_top_iw_I\[15\].genblk1.cell0_I net498 net423 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_2365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput407 um_ow[8] vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__clkbuf_2
Xinput418 um_ow[9] vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_2
Xcol\[3\].zbuf_top_iw_I\[1\].genblk1.cell0_I net491 net428 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_2785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_2685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_sel_I\[3\].genblk1.cell0_I net29 net516 vssd1 vssd1 vccd1 vccd1 zbuf_bus_sel_I\[3\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_13_2562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput226 um_ow[272] vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput204 um_ow[252] vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__clkbuf_2
Xinput215 um_ow[262] vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput237 um_ow[282] vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_2
Xinput248 um_ow[292] vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_1
Xinput259 um_ow[301] vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_2893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_top_iw_I\[14\].genblk1.cell0_I net500 net419 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_2602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_2471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[4\].zbuf_top_iw_I\[9\].genblk1.cell0_I net475 net425 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_309 col\[0\].genblk1.tbuf_spine_ow_I\[1\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].zbuf_top_iw_I\[4\].genblk1.cell0_I net486 net422 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_2633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.tbuf_spine_ow_I\[17\].cell0_I col\[4\].genblk1.mux4_I\[17\].x net440
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[17\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_139 col\[0\].genblk1.tbuf_spine_ow_I\[8\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_117 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_128 col\[0\].genblk1.tbuf_spine_ow_I\[7\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_280_ col\[2\].zbuf_top_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[103] sky130_fd_sc_hd__buf_2
XFILLER_0_11_2863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_35 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_46 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_57 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_2605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_79 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_2739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_2374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xzbuf_bus_iw_I\[9\].genblk1.cell0_I net18 net514 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[9\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout510 col\[0\].zbuf_bot_iw_I\[0\].a vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__clkbuf_4
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_401_ col\[6\].zbuf_bot_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[224] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_332_ col\[4\].zbuf_bot_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[155] sky130_fd_sc_hd__buf_2
XFILLER_0_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_263_ col\[2\].zbuf_bot_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[86] sky130_fd_sc_hd__buf_2
X_194_ col\[0\].zbuf_bot_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[17] sky130_fd_sc_hd__clkbuf_4
Xtbuf_spine_ow_I\[22\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[22\].z net513 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[22\].z sky130_fd_sc_hd__ebufn_1
XFILLER_0_12_2435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_39 col\[0\].genblk1.tbuf_spine_ow_I\[1\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 col\[0\].genblk1.tbuf_spine_ow_I\[12\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_17 col\[0\].genblk1.tbuf_spine_ow_I\[11\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_2181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[4\].genblk1.mux4_I\[18\].cell0_I net158 net184 net210 net237 net469 net455 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[18\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.tbuf_spine_ow_I\[3\].cell0_I col\[6\].genblk1.mux4_I\[3\].x net436
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[3\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_2092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_2057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_2788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_315_ col\[3\].zbuf_top_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[138] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_2455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_2444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_246_ col\[1\].zbuf_top_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[69] sky130_fd_sc_hd__buf_2
Xinput37 um_ow[101] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_0_2499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput26 spine_iw[29] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
Xinput15 spine_iw[19] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
Xinput59 um_ow[121] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_2
X_177_ col\[0\].zbuf_bot_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[0] sky130_fd_sc_hd__buf_2
Xinput48 um_ow[111] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[0\].zbuf_top_iw_I\[15\].genblk1.cell0_I net497 net433 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.tbuf_spine_ow_I\[10\].cell0_I col\[6\].genblk1.mux4_I\[10\].x net436
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[10\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_12_1597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput408 um_ow[90] vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_100_ _031_ vssd1 vssd1 vccd1 vccd1 col\[7\].zbuf_top_ena_I.e sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[4\].zbuf_bot_iw_I\[17\].genblk1.cell0_I net493 col\[4\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[4\].zbuf_bot_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_2697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_229_ col\[1\].zbuf_bot_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[52] sky130_fd_sc_hd__buf_2
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_2406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[13\].genblk1.cell1_I zbuf_bus_iw_I\[13\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[13\].a sky130_fd_sc_hd__buf_6
XFILLER_0_1_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput227 um_ow[273] vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput216 um_ow[263] vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput205 um_ow[253] vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput238 um_ow[283] vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_2
Xinput249 um_ow[293] vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_1
Xcol\[2\].zbuf_top_iw_I\[14\].genblk1.cell0_I net499 net429 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_2572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_2715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_2358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_2093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].zbuf_bot_iw_I\[16\].genblk1.cell0_I net496 col\[6\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[6\].zbuf_bot_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xzbuf_bus_iw_I\[0\].genblk1.cell1_I zbuf_bus_iw_I\[0\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[0\].a sky130_fd_sc_hd__buf_6
XFILLER_0_3_2601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[2\].zbuf_bot_iw_I\[7\].genblk1.cell0_I net479 col\[2\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[2\].zbuf_bot_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_2781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[4\].zbuf_bot_iw_I\[2\].genblk1.cell0_I net489 col\[4\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[4\].zbuf_bot_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_1833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[4\].zbuf_top_iw_I\[13\].genblk1.cell0_I net501 net425 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_2188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_107 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_129 col\[0\].genblk1.tbuf_spine_ow_I\[7\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_118 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcol\[2\].genblk1.tbuf_spine_ow_I\[2\].cell0_I col\[2\].genblk1.mux4_I\[2\].x net442
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[2\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_4_2932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_2897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[0\].genblk1.mux4_I\[13\].cell0_I net79 net345 net376 net402 net462 net448 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[13\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_9_2854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[0\].zbuf_top_iw_I\[6\].genblk1.cell0_I net481 net434 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XTAP_36 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_47 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_58 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_69 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_2617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[2\].zbuf_top_iw_I\[1\].genblk1.cell0_I net491 net430 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_15_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_2206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout500 col\[0\].zbuf_bot_iw_I\[14\].a vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__clkbuf_4
Xfanout511 net513 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_400_ col\[6\].zbuf_bot_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[223] sky130_fd_sc_hd__buf_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_331_ col\[4\].zbuf_bot_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[154] sky130_fd_sc_hd__buf_2
XFILLER_0_7_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_262_ col\[2\].zbuf_bot_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[85] sky130_fd_sc_hd__buf_2
X_193_ col\[0\].zbuf_bot_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[16] sky130_fd_sc_hd__clkbuf_4
Xcol\[6\].zbuf_top_iw_I\[12\].genblk1.cell0_I net504 net421 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_29 col\[0\].genblk1.tbuf_spine_ow_I\[19\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_18 col\[0\].genblk1.tbuf_spine_ow_I\[11\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcol\[2\].genblk1.mux4_I\[23\].cell0_I net56 net83 net109 net136 net465 net450 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[23\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_2193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_bot_iw_I\[5\].genblk1.cell0_I net484 col\[7\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[7\].zbuf_bot_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_2025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.mux4_I\[0\].cell0_I net243 net271 net297 net324 net473 net459 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[0\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_15_2071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].genblk1.tbuf_spine_ow_I\[7\].cell0_I col\[6\].genblk1.mux4_I\[7\].x net437
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[7\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_11_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_314_ col\[3\].zbuf_top_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[137] sky130_fd_sc_hd__buf_2
X_245_ col\[1\].zbuf_top_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[68] sky130_fd_sc_hd__buf_2
Xinput27 spine_iw[2] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput16 spine_iw[1] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_0_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput49 um_ow[112] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput38 um_ow[102] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__dlymetal6s2s_1
X_176_ col\[7\].zbuf_top_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[15] sky130_fd_sc_hd__buf_2
Xcol\[3\].zbuf_top_iw_I\[9\].genblk1.cell0_I net475 net427 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_2345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_2389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_290 col\[0\].genblk1.tbuf_spine_ow_I\[9\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.tbuf_spine_ow_I\[14\].cell0_I col\[6\].genblk1.mux4_I\[14\].x net436
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[14\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_12_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput409 um_ow[91] vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__clkbuf_1
Xcol\[5\].zbuf_top_iw_I\[4\].genblk1.cell0_I net486 net424 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[4\].genblk1.tbuf_row_ena_I.cell0_I col\[4\].genblk1.tbuf_row_ena_I.t vssd1 vssd1
+ vccd1 vccd1 col\[4\].genblk1.tbuf_row_ena_I.tx sky130_fd_sc_hd__inv_2
XFILLER_0_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_228_ col\[1\].zbuf_bot_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[51] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_159_ tbuf_spine_ow_I\[22\].z vssd1 vssd1 vccd1 vccd1 spine_ow[23] sky130_fd_sc_hd__buf_4
XFILLER_0_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_2153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_2197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput217 um_ow[264] vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput206 um_ow[254] vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_11_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput239 um_ow[284] vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput228 um_ow[274] vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[6\].genblk1.mux4_I\[10\].cell0_I net254 net282 net308 net335 net471 net457 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[10\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_2_2304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[2\].genblk1.tbuf_spine_ow_I\[21\].cell0_I col\[2\].genblk1.mux4_I\[21\].x net441
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[21\].z sky130_fd_sc_hd__ebufn_8
Xcol\[1\].zbuf_bot_iw_I\[16\].genblk1.cell0_I net495 col\[1\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[1\].zbuf_bot_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_1525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_2793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[1\].cell0_I net138 net165 net192 net218 net470 net456 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[1\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_10_2534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[1\].zbuf_top_ena_I.genblk1.cell0_I net539 net432 vssd1 vssd1 vccd1 vccd1 col\[1\].zbuf_top_ena_I.z
+ sky130_fd_sc_hd__and2_1
XFILLER_0_8_1801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_2281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_119 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_108 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[2\].genblk1.tbuf_spine_ow_I\[6\].cell0_I col\[2\].genblk1.mux4_I\[6\].x net442
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_10_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_37 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_48 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_59 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_2629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].genblk1.mux4_I\[17\].cell0_I net123 net354 net380 net406 net461 net447 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[17\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_3_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[3\].zbuf_bot_iw_I\[15\].genblk1.cell0_I net497 col\[3\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[3\].zbuf_bot_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout501 col\[0\].zbuf_bot_iw_I\[13\].a vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__buf_6
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout512 net513 vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_330_ col\[4\].zbuf_bot_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[153] sky130_fd_sc_hd__buf_2
Xcol\[1\].zbuf_top_iw_I\[12\].genblk1.cell0_I net503 net431 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_261_ col\[2\].zbuf_bot_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[84] sky130_fd_sc_hd__buf_2
X_192_ col\[0\].zbuf_bot_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_1961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xzbuf_bus_sel_I\[2\].genblk1.cell1_I zbuf_bus_sel_I\[2\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 zbuf_bus_sel_I\[2\].z sky130_fd_sc_hd__buf_6
XFILLER_0_9_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_19 col\[0\].genblk1.tbuf_spine_ow_I\[11\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_459_ col\[7\].zbuf_top_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[282] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_2037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_2083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[6\].genblk1.mux4_I\[4\].cell0_I net248 net275 net302 net328 net473 net459 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[4\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_15_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[5\].zbuf_bot_iw_I\[14\].genblk1.cell0_I net500 col\[5\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[5\].zbuf_bot_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_313_ col\[3\].zbuf_top_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[136] sky130_fd_sc_hd__buf_2
X_244_ col\[1\].zbuf_top_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[67] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput17 spine_iw[20] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
Xinput28 spine_iw[3] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput39 um_ow[103] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__dlymetal6s2s_1
X_175_ col\[7\].zbuf_bot_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[14] sky130_fd_sc_hd__buf_2
XFILLER_0_0_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_280 col\[0\].genblk1.tbuf_spine_ow_I\[3\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_291 col\[0\].genblk1.tbuf_spine_ow_I\[9\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_2267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[2\].genblk1.mux4_I\[2\].cell0_I net416 net60 net86 net113 net466 net452 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[2\].x sky130_fd_sc_hd__mux4_1
Xcol\[3\].zbuf_top_iw_I\[11\].genblk1.cell0_I net505 net427 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].genblk1.tbuf_spine_ow_I\[18\].cell0_I col\[6\].genblk1.mux4_I\[18\].x net435
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[18\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[1\].zbuf_bot_iw_I\[7\].genblk1.cell0_I net479 col\[1\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[1\].zbuf_bot_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].genblk1.tbuf_spine_ow_I\[10\].cell0_I col\[0\].genblk1.mux4_I\[10\].x net445
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[10\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_8_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[3\].zbuf_bot_iw_I\[2\].genblk1.cell0_I net489 col\[3\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[3\].zbuf_bot_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_227_ col\[1\].zbuf_bot_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[50] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_158_ tbuf_spine_ow_I\[21\].z vssd1 vssd1 vccd1 vccd1 spine_ow[22] sky130_fd_sc_hd__buf_4
XFILLER_0_0_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_089_ _025_ vssd1 vssd1 vccd1 vccd1 col\[5\].zbuf_bot_ena_I.e sky130_fd_sc_hd__clkbuf_4
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[7\].zbuf_bot_iw_I\[13\].genblk1.cell0_I net502 col\[7\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[7\].zbuf_bot_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_2121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput218 um_ow[265] vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput207 um_ow[255] vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput229 um_ow[275] vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_7_2920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[6\].zbuf_bot_ena_I.genblk1.cell0_I net548 col\[6\].zbuf_bot_ena_I.e vssd1 vssd1
+ vccd1 vccd1 col\[6\].zbuf_bot_ena_I.z sky130_fd_sc_hd__and2_1
XFILLER_0_14_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[5\].zbuf_top_iw_I\[10\].genblk1.cell0_I net508 net423 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[10\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_iw_I\[1\].genblk1.cell0_I net491 net432 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_2351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.mux4_I\[14\].cell0_I net260 net286 net313 net339 net472 net457 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[14\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_13_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_2084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xzbuf_bus_iw_I\[8\].genblk1.cell1_I zbuf_bus_iw_I\[8\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[8\].a sky130_fd_sc_hd__buf_6
XFILLER_0_14_2126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[5\].cell0_I net142 net170 net196 net222 net470 net454 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[5\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_10_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].zbuf_bot_iw_I\[5\].genblk1.cell0_I net484 col\[6\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[6\].zbuf_bot_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_2293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_2181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_2157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_109 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].genblk1.mux4_I\[3\].cell0_I net352 net234 net365 net391 net463 net449 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[3\].x sky130_fd_sc_hd__mux4_2
Xcol\[2\].zbuf_top_iw_I\[9\].genblk1.cell0_I net475 net429 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_38 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_49 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[4\].zbuf_top_iw_I\[4\].genblk1.cell0_I net485 net426 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[4\].z sky130_fd_sc_hd__and2_1
Xinput390 um_ow[74] vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_2322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout502 col\[0\].zbuf_bot_iw_I\[13\].a vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__clkbuf_4
Xfanout513 tbuf_row_ena_I.tx vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__buf_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_2617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[17\].genblk1.cell0_I net26 net514 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[17\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_7_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_260_ col\[2\].zbuf_bot_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[83] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_191_ col\[0\].zbuf_bot_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_458_ col\[7\].zbuf_top_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[281] sky130_fd_sc_hd__buf_2
X_389_ col\[5\].zbuf_top_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[212] sky130_fd_sc_hd__buf_2
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_bot_iw_I\[14\].genblk1.cell0_I net499 col\[0\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[0\].zbuf_bot_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_11_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.mux4_I\[8\].cell0_I net252 net280 net306 net332 net473 net459 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[8\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_312_ col\[3\].zbuf_top_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[135] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_2561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_243_ col\[1\].zbuf_top_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[66] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 spine_iw[21] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
Xinput29 spine_iw[4] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__dlymetal6s2s_1
X_174_ col\[6\].zbuf_top_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[13] sky130_fd_sc_hd__buf_2
XFILLER_0_11_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xzbuf_bus_iw_I\[4\].genblk1.cell0_I net12 net515 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[4\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XANTENNA_270 col\[0\].genblk1.tbuf_spine_ow_I\[2\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_281 col\[0\].genblk1.tbuf_spine_ow_I\[3\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_292 col\[0\].genblk1.tbuf_spine_ow_I\[9\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_2071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[7\].zbuf_top_iw_I\[7\].genblk1.cell0_I net480 net420 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.mux4_I\[6\].cell0_I net38 net64 net91 net117 net466 net452 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[6\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_1_2723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_2701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[0\].genblk1.tbuf_spine_ow_I\[14\].cell0_I col\[0\].genblk1.mux4_I\[14\].x net445
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[14\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_1_2789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtbuf_spine_ow_I\[12\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[12\].z net512 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[12\].z sky130_fd_sc_hd__ebufn_1
XFILLER_0_6_2623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_2500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_2288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_226_ col\[1\].zbuf_bot_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[49] sky130_fd_sc_hd__buf_2
X_157_ tbuf_spine_ow_I\[20\].z vssd1 vssd1 vccd1 vccd1 spine_ow[21] sky130_fd_sc_hd__buf_4
Xcol\[2\].zbuf_bot_iw_I\[13\].genblk1.cell0_I net501 col\[2\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[2\].zbuf_bot_iw_I\[13\].z sky130_fd_sc_hd__and2_1
X_088_ _013_ net460 _023_ vssd1 vssd1 vccd1 vccd1 _025_ sky130_fd_sc_hd__and3b_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_2177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput208 um_ow[256] vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput219 um_ow[266] vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_14_2820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_2807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_2829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].zbuf_top_iw_I\[10\].genblk1.cell0_I net507 net433 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_2063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_209_ col\[0\].zbuf_top_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[32] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[6\].genblk1.mux4_I\[18\].cell0_I net264 net291 net317 net343 net472 net458 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[18\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_1_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_2862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[4\].zbuf_bot_iw_I\[12\].genblk1.cell0_I net503 col\[4\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[4\].zbuf_bot_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[4\].genblk1.mux4_I\[9\].cell0_I net148 net174 net200 net227 net468 net454 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[9\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_15_2414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].genblk1.mux4_I\[7\].cell0_I net396 net279 net369 net395 net462 net448 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[7\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_9_2813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_39 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_2480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput380 um_ow[65] vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__clkbuf_1
Xinput391 um_ow[75] vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_2211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[0\].zbuf_bot_iw_I\[7\].genblk1.cell0_I net479 col\[0\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[0\].zbuf_bot_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_2288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].zbuf_bot_iw_I\[11\].genblk1.cell0_I net506 col\[6\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[6\].zbuf_bot_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout503 col\[0\].zbuf_bot_iw_I\[12\].a vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__buf_6
Xfanout514 net515 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].zbuf_bot_iw_I\[2\].genblk1.cell0_I net489 col\[2\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[2\].zbuf_bot_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_2629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_2798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_190_ col\[0\].zbuf_bot_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[13] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_2687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_457_ col\[7\].zbuf_top_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[280] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_388_ col\[5\].zbuf_top_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[211] sky130_fd_sc_hd__buf_2
XFILLER_0_3_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_top_iw_I\[1\].genblk1.cell0_I net491 net434 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[4\].genblk1.tbuf_spine_ow_I\[22\].cell0_I col\[4\].genblk1.mux4_I\[22\].x net438
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[22\].z sky130_fd_sc_hd__ebufn_8
X_311_ col\[3\].zbuf_top_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[134] sky130_fd_sc_hd__buf_2
XFILLER_0_4_2573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_242_ col\[1\].zbuf_top_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[65] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_173_ col\[6\].zbuf_bot_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[12] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput19 spine_iw[22] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_1793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_260 col\[0\].genblk1.tbuf_spine_ow_I\[2\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_271 col\[0\].genblk1.tbuf_spine_ow_I\[2\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_293 col\[0\].genblk1.tbuf_spine_ow_I\[9\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_282 col\[0\].genblk1.tbuf_spine_ow_I\[3\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_2225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[0\].genblk1.tbuf_spine_ow_I\[18\].cell0_I col\[0\].genblk1.mux4_I\[18\].x net445
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[18\].z sky130_fd_sc_hd__ebufn_8
Xtbuf_spine_ow_I\[16\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[16\].z net511 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[16\].z sky130_fd_sc_hd__ebufn_1
Xcol\[5\].zbuf_bot_iw_I\[5\].genblk1.cell0_I net484 col\[5\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[5\].zbuf_bot_iw_I\[5\].z sky130_fd_sc_hd__and2_1
Xcol\[2\].genblk1.mux4_I\[13\].cell0_I net45 net72 net98 net125 net465 net451 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[13\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_6_2602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_2381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_225_ col\[1\].zbuf_bot_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[48] sky130_fd_sc_hd__buf_2
X_156_ tbuf_spine_ow_I\[19\].z vssd1 vssd1 vccd1 vccd1 spine_ow[20] sky130_fd_sc_hd__buf_4
XFILLER_0_0_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_087_ _024_ vssd1 vssd1 vccd1 vccd1 col\[4\].zbuf_top_ena_I.e sky130_fd_sc_hd__clkbuf_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[7\].zbuf_bot_iw_I\[0\].genblk1.cell0_I net510 col\[7\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[7\].zbuf_bot_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput209 um_ow[257] vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__dlymetal6s2s_1
Xcol\[1\].zbuf_top_iw_I\[9\].genblk1.cell0_I net475 net431 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_2900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[3\].zbuf_top_iw_I\[4\].genblk1.cell0_I net485 net428 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_2432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[23\].cell0_I net163 net189 net216 net242 net469 net455 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[23\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_5_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_208_ col\[0\].zbuf_top_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[31] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_139_ tbuf_spine_ow_I\[2\].z vssd1 vssd1 vccd1 vccd1 spine_ow[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_2117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_2673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].genblk1.tbuf_row_ena_I.cell0_I col\[0\].genblk1.tbuf_row_ena_I.t vssd1 vssd1
+ vccd1 vccd1 col\[0\].genblk1.tbuf_row_ena_I.tx sky130_fd_sc_hd__inv_2
XFILLER_0_8_2549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[7\].zbuf_top_iw_I\[17\].genblk1.cell0_I net494 net419 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_15_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_2835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_2879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[4\].genblk1.tbuf_spine_ow_I\[2\].cell0_I col\[4\].genblk1.mux4_I\[2\].x net439
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[2\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_9_2825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_2424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[2\].genblk1.tbuf_spine_ow_I\[11\].cell0_I col\[2\].genblk1.mux4_I\[11\].x net443
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[11\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_10_2378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].zbuf_top_iw_I\[7\].genblk1.cell0_I net480 net422 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[7\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_bot_iw_I\[11\].genblk1.cell0_I net505 col\[1\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[1\].zbuf_bot_iw_I\[11\].z sky130_fd_sc_hd__and2_1
Xinput381 um_ow[66] vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__clkbuf_1
Xinput370 um_ow[56] vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__clkbuf_1
Xinput392 um_ow[76] vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_2234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_2081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout504 col\[0\].zbuf_bot_iw_I\[12\].a vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout515 tbuf_row_ena_I.t vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__clkbuf_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_2733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_456_ col\[7\].zbuf_top_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[279] sky130_fd_sc_hd__buf_2
X_387_ col\[5\].zbuf_top_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[210] sky130_fd_sc_hd__buf_2
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_310_ col\[3\].zbuf_top_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[133] sky130_fd_sc_hd__buf_2
Xcol\[3\].zbuf_bot_iw_I\[10\].genblk1.cell0_I net507 col\[3\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[3\].zbuf_bot_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_2585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_241_ col\[1\].zbuf_top_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[64] sky130_fd_sc_hd__buf_2
X_172_ col\[5\].zbuf_top_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[11] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_250 col\[0\].genblk1.tbuf_spine_ow_I\[18\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_261 col\[0\].genblk1.tbuf_spine_ow_I\[2\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_272 col\[0\].genblk1.tbuf_spine_ow_I\[3\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_294 col\[0\].genblk1.tbuf_spine_ow_I\[9\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_283 col\[0\].genblk1.tbuf_spine_ow_I\[3\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_2237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_439_ col\[7\].zbuf_bot_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[262] sky130_fd_sc_hd__buf_2
XFILLER_0_3_2073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_2872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.mux4_I\[17\].cell0_I net50 net76 net103 net129 net465 net451 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[17\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_6_1913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_2393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_224_ col\[1\].zbuf_bot_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[47] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_155_ tbuf_spine_ow_I\[18\].z vssd1 vssd1 vccd1 vccd1 spine_ow[19] sky130_fd_sc_hd__buf_4
X_086_ _011_ _023_ net470 vssd1 vssd1 vccd1 vccd1 _024_ sky130_fd_sc_hd__and3b_1
XFILLER_0_0_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_2001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].genblk1.tbuf_spine_ow_I\[1\].cell0_I col\[0\].genblk1.mux4_I\[1\].x net444
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[1\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_8_2709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_2411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_207_ col\[0\].zbuf_top_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[30] sky130_fd_sc_hd__buf_2
X_138_ tbuf_spine_ow_I\[1\].z vssd1 vssd1 vccd1 vccd1 spine_ow[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_069_ _014_ vssd1 vssd1 vccd1 vccd1 col\[0\].zbuf_top_ena_I.e sky130_fd_sc_hd__clkbuf_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[1\].zbuf_bot_iw_I\[2\].genblk1.cell0_I net489 col\[1\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[1\].zbuf_bot_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[16\].genblk1.cell1_I zbuf_bus_iw_I\[16\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[16\].a sky130_fd_sc_hd__buf_6
XFILLER_0_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].zbuf_top_iw_I\[17\].genblk1.cell0_I net493 net429 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.tbuf_spine_ow_I\[6\].cell0_I col\[4\].genblk1.mux4_I\[6\].x net439
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_14_2471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[2\].zbuf_bot_ena_I.genblk1.cell0_I net540 col\[2\].zbuf_bot_ena_I.e vssd1 vssd1
+ vccd1 vccd1 col\[2\].zbuf_bot_ena_I.z sky130_fd_sc_hd__and2_1
XFILLER_0_3_2436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.tbuf_spine_ow_I\[15\].cell0_I col\[2\].genblk1.mux4_I\[15\].x net441
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[15\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_11_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[3\].genblk1.cell1_I zbuf_bus_iw_I\[3\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[3\].a sky130_fd_sc_hd__buf_6
Xinput360 um_ow[47] vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__clkbuf_2
Xinput371 um_ow[57] vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_1
Xinput393 um_ow[77] vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__clkbuf_1
Xinput382 um_ow[67] vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_2891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout505 col\[0\].zbuf_bot_iw_I\[11\].a vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__buf_6
XFILLER_0_1_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[4\].zbuf_bot_iw_I\[5\].genblk1.cell0_I net483 col\[4\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[4\].zbuf_bot_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout516 tbuf_row_ena_I.t vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__buf_2
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[4\].zbuf_top_iw_I\[16\].genblk1.cell0_I net495 net425 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_2745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].zbuf_bot_iw_I\[0\].genblk1.cell0_I net510 col\[6\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[6\].zbuf_bot_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_455_ col\[7\].zbuf_top_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[278] sky130_fd_sc_hd__buf_2
XFILLER_0_14_2290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_386_ col\[5\].zbuf_top_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[209] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_top_iw_I\[9\].genblk1.cell0_I net475 net434 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[9\].z sky130_fd_sc_hd__and2_1
Xinput190 um_ow[23] vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_8_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_2920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[2\].zbuf_top_iw_I\[4\].genblk1.cell0_I net485 net430 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_2829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_240_ col\[1\].zbuf_top_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[63] sky130_fd_sc_hd__buf_2
XFILLER_0_4_2597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_171_ col\[5\].zbuf_bot_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[10] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_2496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_240 col\[0\].genblk1.tbuf_spine_ow_I\[17\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_251 col\[0\].genblk1.tbuf_spine_ow_I\[18\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_262 col\[0\].genblk1.tbuf_spine_ow_I\[2\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_2041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_284 col\[0\].genblk1.tbuf_spine_ow_I\[3\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_295 col\[0\].genblk1.tbuf_spine_ow_I\[9\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_273 col\[0\].genblk1.tbuf_spine_ow_I\[3\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_2249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_438_ col\[7\].zbuf_bot_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[261] sky130_fd_sc_hd__buf_2
XFILLER_0_3_2085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_369_ col\[5\].zbuf_bot_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[192] sky130_fd_sc_hd__buf_2
Xcol\[6\].zbuf_top_iw_I\[15\].genblk1.cell0_I net498 net421 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_10_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xzbuf_bus_iw_I\[12\].genblk1.cell0_I net21 net516 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[12\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_1_2715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[7\].zbuf_bot_iw_I\[8\].genblk1.cell0_I net478 col\[7\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[7\].zbuf_bot_iw_I\[8\].z sky130_fd_sc_hd__and2_1
Xcol\[0\].genblk1.mux4_I\[22\].cell0_I net179 net359 net386 net412 net461 net447 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[22\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_9_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_2637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_223_ col\[1\].zbuf_bot_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[46] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_154_ tbuf_spine_ow_I\[17\].z vssd1 vssd1 vccd1 vccd1 spine_ow[18] sky130_fd_sc_hd__buf_4
XFILLER_0_11_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_085_ zbuf_bus_ena_I.z col\[4\].genblk1.tbuf_row_ena_I.t vssd1 vssd1 vccd1 vccd1
+ _023_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_2709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[5\].zbuf_top_iw_I\[7\].genblk1.cell0_I net480 net424 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[7\].z sky130_fd_sc_hd__and2_1
Xcol\[6\].zbuf_top_ena_I.genblk1.cell0_I net549 net422 vssd1 vssd1 vccd1 vccd1 col\[6\].zbuf_top_ena_I.z
+ sky130_fd_sc_hd__and2_1
Xcol\[0\].genblk1.tbuf_spine_ow_I\[5\].cell0_I col\[0\].genblk1.mux4_I\[5\].x net444
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[5\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_2609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_top_iw_I\[2\].genblk1.cell0_I net490 net420 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_2099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_206_ col\[0\].zbuf_top_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[29] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_137_ tbuf_spine_ow_I\[0\].z vssd1 vssd1 vccd1 vccd1 spine_ow[1] sky130_fd_sc_hd__clkbuf_4
Xcol\[0\].zbuf_bot_ena_I.genblk1.cell0_I_536 vssd1 vssd1 vccd1 vccd1 net536 col\[0\].zbuf_bot_ena_I.genblk1.cell0_I_536/LO
+ sky130_fd_sc_hd__conb_1
X_068_ _011_ _012_ _013_ vssd1 vssd1 vccd1 vccd1 _014_ sky130_fd_sc_hd__and3b_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtbuf_spine_ow_I\[2\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[2\].z net512 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[2\].z sky130_fd_sc_hd__ebufn_1
XFILLER_0_14_2108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_2743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[6\].genblk1.tbuf_spine_ow_I\[23\].cell0_I col\[6\].genblk1.mux4_I\[23\].x net435
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[23\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_0_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_2404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.tbuf_spine_ow_I\[19\].cell0_I col\[2\].genblk1.mux4_I\[19\].x net441
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[19\].z sky130_fd_sc_hd__ebufn_8
Xinput350 um_ow[38] vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__clkbuf_2
Xinput372 um_ow[58] vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__clkbuf_1
Xinput361 um_ow[48] vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__clkbuf_1
Xinput394 um_ow[78] vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__clkbuf_1
Xinput383 um_ow[68] vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[1\].zbuf_bot_ena_I.genblk1.cell0_I_538 vssd1 vssd1 vccd1 vccd1 net538 col\[1\].zbuf_bot_ena_I.genblk1.cell0_I_538/LO
+ sky130_fd_sc_hd__conb_1
Xfanout506 col\[0\].zbuf_bot_iw_I\[11\].a vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__clkbuf_4
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_2613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_454_ col\[7\].zbuf_top_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[277] sky130_fd_sc_hd__buf_2
XFILLER_0_3_2245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_2267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_385_ col\[5\].zbuf_top_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[208] sky130_fd_sc_hd__buf_2
XFILLER_0_10_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput180 um_ow[230] vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_2101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput191 um_ow[240] vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_8_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_2808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_170_ col\[4\].zbuf_top_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[9] sky130_fd_sc_hd__buf_2
XFILLER_0_4_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].zbuf_bot_iw_I\[2\].genblk1.cell0_I net489 col\[0\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[0\].zbuf_bot_iw_I\[2\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_iw_I\[15\].genblk1.cell0_I net497 net431 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_230 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_241 col\[0\].genblk1.tbuf_spine_ow_I\[17\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_252 col\[0\].genblk1.tbuf_spine_ow_I\[18\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_263 col\[0\].genblk1.tbuf_spine_ow_I\[2\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_285 col\[0\].genblk1.tbuf_spine_ow_I\[3\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_274 col\[0\].genblk1.tbuf_spine_ow_I\[3\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_437_ col\[7\].zbuf_bot_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[260] sky130_fd_sc_hd__buf_2
XFILLER_0_3_2053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_296 col\[0\].genblk1.tbuf_spine_ow_I\[9\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_368_ col\[5\].zbuf_bot_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[191] sky130_fd_sc_hd__buf_2
XFILLER_0_3_2097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_299_ col\[3\].zbuf_bot_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[122] sky130_fd_sc_hd__buf_2
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_222_ col\[1\].zbuf_bot_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[45] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_153_ tbuf_spine_ow_I\[16\].z vssd1 vssd1 vccd1 vccd1 spine_ow[17] sky130_fd_sc_hd__buf_4
Xcol\[5\].zbuf_bot_iw_I\[17\].genblk1.cell0_I net494 col\[5\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[5\].zbuf_bot_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_084_ _022_ vssd1 vssd1 vccd1 vccd1 col\[4\].zbuf_bot_ena_I.e sky130_fd_sc_hd__buf_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_2025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_2069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.tbuf_spine_ow_I\[12\].cell0_I col\[4\].genblk1.mux4_I\[12\].x net438
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[12\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[3\].zbuf_top_iw_I\[14\].genblk1.cell0_I net499 net427 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_2546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].genblk1.tbuf_spine_ow_I\[9\].cell0_I col\[0\].genblk1.mux4_I\[9\].x net445
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[9\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_13_2345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_205_ col\[0\].zbuf_top_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[28] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_067_ net467 vssd1 vssd1 vccd1 vccd1 _013_ sky130_fd_sc_hd__buf_6
XFILLER_0_0_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[3\].zbuf_bot_iw_I\[5\].genblk1.cell0_I net483 col\[3\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[3\].zbuf_bot_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtbuf_spine_ow_I\[6\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[6\].z net512 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[6\].z sky130_fd_sc_hd__ebufn_2
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[5\].zbuf_bot_iw_I\[0\].genblk1.cell0_I net510 col\[5\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[5\].zbuf_bot_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[7\].zbuf_bot_iw_I\[16\].genblk1.cell0_I net496 col\[7\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[7\].zbuf_bot_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_2799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_2129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[5\].zbuf_top_iw_I\[13\].genblk1.cell0_I net502 net423 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[13\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_iw_I\[4\].genblk1.cell0_I net485 net432 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[4\].genblk1.mux4_I\[13\].cell0_I net152 net178 net205 net231 net468 net454 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[13\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_7_2585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xzbuf_bus_sel_I\[1\].genblk1.cell0_I net27 net516 vssd1 vssd1 vccd1 vccd1 zbuf_bus_sel_I\[1\].genblk1.l
+ sky130_fd_sc_hd__and2_1
Xinput351 um_ow[39] vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_2
Xinput340 um_ow[375] vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput362 um_ow[49] vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_1
Xinput395 um_ow[79] vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__clkbuf_1
Xinput384 um_ow[69] vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__clkbuf_1
Xinput373 um_ow[59] vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_2226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].zbuf_bot_iw_I\[8\].genblk1.cell0_I net478 col\[6\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[6\].zbuf_bot_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout507 col\[0\].zbuf_bot_iw_I\[10\].a vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__buf_6
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_2725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_2769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_2624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_2471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[7\].zbuf_top_iw_I\[12\].genblk1.cell0_I net504 net419 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[2\].zbuf_top_ena_I.genblk1.cell0_I_541 vssd1 vssd1 vccd1 vccd1 net541 col\[2\].zbuf_top_ena_I.genblk1.cell0_I_541/LO
+ sky130_fd_sc_hd__conb_1
Xcol\[6\].genblk1.mux4_I\[23\].cell0_I net270 net296 net322 net349 net471 net457 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[23\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_9_2669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_453_ col\[7\].zbuf_top_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[276] sky130_fd_sc_hd__buf_2
XFILLER_0_14_2281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_384_ col\[5\].zbuf_top_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[207] sky130_fd_sc_hd__buf_2
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput170 um_ow[221] vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_1
Xinput181 um_ow[231] vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_2113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput192 um_ow[241] vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_15_2001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[4\].zbuf_top_iw_I\[7\].genblk1.cell0_I net479 net426 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_2708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_2465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].zbuf_top_iw_I\[2\].genblk1.cell0_I net490 net422 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_220 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_231 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_242 col\[0\].genblk1.tbuf_spine_ow_I\[17\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_264 col\[0\].genblk1.tbuf_spine_ow_I\[2\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_253 col\[0\].genblk1.tbuf_spine_ow_I\[18\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_286 col\[0\].genblk1.tbuf_spine_ow_I\[3\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_275 col\[0\].genblk1.tbuf_spine_ow_I\[3\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_2207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_297 col\[0\].zbuf_bot_iw_I\[0\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_2920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_436_ col\[7\].zbuf_bot_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[259] sky130_fd_sc_hd__buf_2
XFILLER_0_3_2065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_367_ col\[5\].zbuf_bot_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[190] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_298_ col\[3\].zbuf_bot_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[121] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_2741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].zbuf_bot_iw_I\[17\].genblk1.cell0_I net493 col\[0\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[0\].zbuf_bot_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_2527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_221_ col\[1\].zbuf_bot_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[44] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_152_ tbuf_spine_ow_I\[15\].z vssd1 vssd1 vccd1 vccd1 spine_ow[16] sky130_fd_sc_hd__buf_4
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_083_ net470 net456 col\[4\].genblk1.tbuf_row_ena_I.t zbuf_bus_ena_I.z vssd1 vssd1
+ vccd1 vccd1 _022_ sky130_fd_sc_hd__and4bb_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[3\].zbuf_top_ena_I.genblk1.cell0_I_543 vssd1 vssd1 vccd1 vccd1 net543 col\[3\].zbuf_top_ena_I.genblk1.cell0_I_543/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_9_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_2127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_419_ col\[6\].zbuf_top_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[242] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[7\].genblk1.cell0_I net15 net514 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[7\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_12_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.tbuf_spine_ow_I\[16\].cell0_I col\[4\].genblk1.mux4_I\[16\].x net438
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[16\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_8_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_2193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_2057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_204_ col\[0\].zbuf_top_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[27] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_066_ zbuf_bus_ena_I.z col\[0\].genblk1.tbuf_row_ena_I.t vssd1 vssd1 vccd1 vccd1
+ _012_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_2878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].zbuf_bot_iw_I\[16\].genblk1.cell0_I net495 col\[2\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[2\].zbuf_bot_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_12_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_2509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].zbuf_top_iw_I\[13\].genblk1.cell0_I net501 net433 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_049_ zbuf_bus_sel_I\[4\].z zbuf_bus_sel_I\[3\].z zbuf_bus_sel_I\[2\].z vssd1 vssd1
+ vccd1 vccd1 col\[2\].genblk1.tbuf_row_ena_I.t sky130_fd_sc_hd__nor3b_4
XFILLER_0_0_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[4\].zbuf_top_ena_I.genblk1.cell0_I_545 vssd1 vssd1 vccd1 vccd1 net545 col\[4\].zbuf_top_ena_I.genblk1.cell0_I_545/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_15_2920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].genblk1.tbuf_spine_ow_I\[23\].cell0_I col\[0\].genblk1.mux4_I\[23\].x net444
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[23\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_2_1930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtbuf_spine_ow_I\[21\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[21\].z net511 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[21\].z sky130_fd_sc_hd__ebufn_1
XFILLER_0_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[4\].genblk1.mux4_I\[17\].cell0_I net156 net183 net209 net236 net469 net455 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[17\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_3_2417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_2575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[6\].genblk1.tbuf_spine_ow_I\[2\].cell0_I col\[6\].genblk1.mux4_I\[2\].x net436
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[2\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_8_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[4\].zbuf_bot_iw_I\[15\].genblk1.cell0_I net497 col\[4\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[4\].zbuf_bot_iw_I\[15\].z sky130_fd_sc_hd__and2_1
Xinput330 um_ow[366] vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput341 um_ow[376] vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput352 um_ow[3] vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__clkbuf_2
Xinput363 um_ow[4] vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__clkbuf_2
Xinput396 um_ow[7] vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__clkbuf_2
Xinput385 um_ow[6] vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput374 um_ow[5] vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_15_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout508 col\[0\].zbuf_bot_iw_I\[10\].a vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_4
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xzbuf_bus_iw_I\[11\].genblk1.cell1_I zbuf_bus_iw_I\[11\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[11\].a sky130_fd_sc_hd__buf_6
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_2840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_2715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].zbuf_top_iw_I\[12\].genblk1.cell0_I net503 net429 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_2361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_452_ col\[7\].zbuf_top_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[275] sky130_fd_sc_hd__buf_2
X_383_ col\[5\].zbuf_top_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[206] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_2113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput171 um_ow[222] vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_1
Xinput160 um_ow[212] vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_1
Xinput182 um_ow[232] vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_1
Xinput193 um_ow[242] vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_8_2125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_2169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_2792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[6\].zbuf_bot_iw_I\[14\].genblk1.cell0_I net500 col\[6\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[6\].zbuf_bot_iw_I\[14\].z sky130_fd_sc_hd__and2_1
Xcol\[5\].zbuf_top_ena_I.genblk1.cell0_I_547 vssd1 vssd1 vccd1 vccd1 net547 col\[5\].zbuf_top_ena_I.genblk1.cell0_I_547/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_4_2523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[2\].zbuf_bot_iw_I\[5\].genblk1.cell0_I net483 col\[2\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[2\].zbuf_bot_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_1711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_221 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_210 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_243 col\[0\].genblk1.tbuf_spine_ow_I\[17\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_232 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_265 col\[0\].genblk1.tbuf_spine_ow_I\[2\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_254 col\[0\].genblk1.tbuf_spine_ow_I\[18\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_276 col\[0\].genblk1.tbuf_spine_ow_I\[3\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_435_ col\[7\].zbuf_bot_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[258] sky130_fd_sc_hd__buf_2
XANTENNA_287 col\[0\].genblk1.tbuf_spine_ow_I\[9\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_298 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_366_ col\[5\].zbuf_bot_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[189] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_297_ col\[3\].zbuf_bot_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[120] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_bot_iw_I\[0\].genblk1.cell0_I net509 col\[4\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[4\].zbuf_bot_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XFILLER_0_11_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_top_iw_I\[11\].genblk1.cell0_I net505 net425 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_2753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_220_ col\[1\].zbuf_bot_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[43] sky130_fd_sc_hd__buf_2
XFILLER_0_11_2241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_151_ tbuf_spine_ow_I\[14\].z vssd1 vssd1 vccd1 vccd1 spine_ow[15] sky130_fd_sc_hd__buf_4
XFILLER_0_9_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_082_ _021_ vssd1 vssd1 vccd1 vccd1 col\[3\].zbuf_top_ena_I.e sky130_fd_sc_hd__clkbuf_1
Xcol\[0\].zbuf_top_iw_I\[4\].genblk1.cell0_I net485 net434 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_418_ col\[6\].zbuf_top_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[241] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_349_ col\[4\].zbuf_top_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[172] sky130_fd_sc_hd__buf_2
XFILLER_0_4_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].zbuf_top_ena_I.genblk1.cell0_I_549 vssd1 vssd1 vccd1 vccd1 net549 col\[6\].zbuf_top_ena_I.genblk1.cell0_I_549/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_6_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[6\].zbuf_top_iw_I\[10\].genblk1.cell0_I net508 net421 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[10\].z sky130_fd_sc_hd__and2_1
X_203_ col\[0\].zbuf_top_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[26] sky130_fd_sc_hd__buf_2
XFILLER_0_13_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[2\].genblk1.tbuf_spine_ow_I\[1\].cell0_I col\[2\].genblk1.mux4_I\[1\].x net442
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[1\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_11_2071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[5\].zbuf_bot_iw_I\[8\].genblk1.cell0_I net478 col\[5\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[5\].zbuf_bot_iw_I\[8\].z sky130_fd_sc_hd__and2_1
X_065_ net453 vssd1 vssd1 vccd1 vccd1 _011_ sky130_fd_sc_hd__buf_6
XFILLER_0_0_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].genblk1.mux4_I\[12\].cell0_I net68 net334 net375 net401 net462 net448 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[12\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_12_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_bot_iw_I\[3\].genblk1.cell0_I net488 col\[7\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[7\].zbuf_bot_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_2267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[3\].zbuf_top_iw_I\[7\].genblk1.cell0_I net479 net428 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_048_ zbuf_bus_sel_I\[4\].z zbuf_bus_sel_I\[2\].z zbuf_bus_sel_I\[3\].z vssd1 vssd1
+ vccd1 vccd1 col\[0\].genblk1.tbuf_row_ena_I.t sky130_fd_sc_hd__nor3_4
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_2790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[5\].zbuf_top_iw_I\[2\].genblk1.cell0_I net490 net424 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_2665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[2\].genblk1.mux4_I\[22\].cell0_I net55 net82 net108 net135 net464 net450 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[22\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_7_2521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].genblk1.tbuf_spine_ow_I\[6\].cell0_I col\[6\].genblk1.mux4_I\[6\].x net437
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[6\].z sky130_fd_sc_hd__ebufn_8
Xcol\[2\].zbuf_top_ena_I.genblk1.cell0_I net541 net430 vssd1 vssd1 vccd1 vccd1 col\[2\].zbuf_top_ena_I.z
+ sky130_fd_sc_hd__and2_1
Xinput320 um_ow[357] vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput342 um_ow[377] vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput353 um_ow[40] vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__clkbuf_2
Xinput331 um_ow[367] vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput397 um_ow[80] vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__clkbuf_1
Xinput386 um_ow[70] vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_1
Xinput375 um_ow[60] vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__clkbuf_1
Xinput364 um_ow[50] vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_1628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_2 _014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout509 col\[0\].zbuf_bot_iw_I\[0\].a vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__buf_8
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_2795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_2451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[6\].genblk1.tbuf_spine_ow_I\[13\].cell0_I col\[6\].genblk1.mux4_I\[13\].x net437
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[13\].z sky130_fd_sc_hd__ebufn_8
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_451_ col\[7\].zbuf_top_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[274] sky130_fd_sc_hd__buf_2
X_382_ col\[5\].zbuf_top_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[205] sky130_fd_sc_hd__buf_2
XFILLER_0_14_2261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput172 um_ow[223] vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_1
Xinput150 um_ow[203] vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_1
Xinput161 um_ow[213] vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__clkbuf_1
Xinput183 um_ow[233] vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_1
Xinput194 um_ow[243] vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_8_2137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[1\].zbuf_bot_iw_I\[14\].genblk1.cell0_I net499 col\[1\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[1\].zbuf_bot_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_2413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_200 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_233 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_222 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_211 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_434_ col\[7\].zbuf_bot_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[257] sky130_fd_sc_hd__buf_2
XANTENNA_255 col\[0\].genblk1.tbuf_spine_ow_I\[18\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_244 col\[0\].genblk1.tbuf_spine_ow_I\[17\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_266 col\[0\].genblk1.tbuf_spine_ow_I\[2\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_277 col\[0\].genblk1.tbuf_spine_ow_I\[3\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_2911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_299 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_288 col\[0\].genblk1.tbuf_spine_ow_I\[9\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_365_ col\[5\].zbuf_bot_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[188] sky130_fd_sc_hd__buf_2
X_296_ col\[3\].zbuf_bot_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[119] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_2619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].genblk1.tbuf_spine_ow_I\[20\].cell0_I col\[2\].genblk1.mux4_I\[20\].x net441
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[20\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_4_1620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_150_ tbuf_spine_ow_I\[13\].z vssd1 vssd1 vccd1 vccd1 spine_ow[14] sky130_fd_sc_hd__buf_4
XFILLER_0_11_2297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_081_ _013_ _011_ _018_ vssd1 vssd1 vccd1 vccd1 _021_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_1596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[3\].zbuf_bot_iw_I\[13\].genblk1.cell0_I net501 col\[3\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[3\].zbuf_bot_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_417_ col\[6\].zbuf_top_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[240] sky130_fd_sc_hd__buf_2
X_348_ col\[4\].zbuf_top_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[171] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_279_ col\[2\].zbuf_top_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[102] sky130_fd_sc_hd__buf_2
XFILLER_0_3_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[4\].genblk1.mux4_I\[0\].cell0_I net137 net164 net191 net217 net470 net456 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[0\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_11_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_2562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[1\].zbuf_top_iw_I\[10\].genblk1.cell0_I net507 net431 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_10_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_202_ col\[0\].zbuf_top_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[25] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xzbuf_bus_sel_I\[0\].genblk1.cell1_I zbuf_bus_sel_I\[0\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 zbuf_bus_sel_I\[0\].z sky130_fd_sc_hd__buf_6
Xcol\[2\].genblk1.tbuf_spine_ow_I\[5\].cell0_I col\[2\].genblk1.mux4_I\[5\].x net442
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[5\].z sky130_fd_sc_hd__ebufn_8
X_064_ _010_ vssd1 vssd1 vccd1 vccd1 col\[0\].zbuf_bot_ena_I.e sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[0\].genblk1.mux4_I\[16\].cell0_I net112 net353 net379 net405 net461 net447 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[16\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_bot_ena_I.genblk1.cell0_I net550 col\[7\].zbuf_bot_ena_I.e vssd1 vssd1
+ vccd1 vccd1 col\[7\].zbuf_bot_ena_I.z sky130_fd_sc_hd__and2_1
XFILLER_0_7_2725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[5\].zbuf_bot_iw_I\[12\].genblk1.cell0_I net504 col\[5\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[5\].zbuf_bot_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_2381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_2900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[1\].zbuf_bot_iw_I\[5\].genblk1.cell0_I net483 col\[1\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[1\].zbuf_bot_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[3\].zbuf_bot_iw_I\[0\].genblk1.cell0_I net509 col\[3\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[3\].zbuf_bot_iw_I\[0\].z sky130_fd_sc_hd__and2_1
Xcol\[6\].genblk1.mux4_I\[3\].cell0_I net247 net274 net300 net327 net473 net459 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[3\].x sky130_fd_sc_hd__mux4_1
Xinput310 um_ow[348] vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__clkbuf_2
Xinput321 um_ow[358] vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput354 um_ow[41] vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_2
Xinput332 um_ow[368] vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput343 um_ow[378] vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput387 um_ow[71] vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__clkbuf_1
Xinput376 um_ow[61] vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__clkbuf_1
Xinput365 um_ow[51] vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_1
Xinput398 um_ow[81] vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_2043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_3 col\[0\].genblk1.tbuf_spine_ow_I\[0\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_bot_iw_I\[11\].genblk1.cell0_I net506 col\[7\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[7\].zbuf_bot_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_10_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_2853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_2875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_2741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_2717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[2\].genblk1.mux4_I\[1\].cell0_I net415 net59 net85 net111 net466 net452 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[1\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[6\].genblk1.tbuf_spine_ow_I\[17\].cell0_I col\[6\].genblk1.mux4_I\[17\].x net435
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[17\].z sky130_fd_sc_hd__ebufn_8
XFILLER_0_9_1905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_450_ col\[7\].zbuf_top_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[273] sky130_fd_sc_hd__buf_2
X_381_ col\[5\].zbuf_top_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[204] sky130_fd_sc_hd__buf_2
XFILLER_0_7_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_2396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput140 um_ow[195] vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_1
Xinput151 um_ow[204] vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__clkbuf_1
Xinput162 um_ow[214] vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_1
Xinput173 um_ow[224] vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_1
Xinput184 um_ow[234] vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_1
Xinput195 um_ow[244] vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_8_2149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[6\].genblk1.cell1_I zbuf_bus_iw_I\[6\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[6\].a sky130_fd_sc_hd__buf_6
XFILLER_0_14_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_2661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_2547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[4\].zbuf_bot_iw_I\[8\].genblk1.cell0_I net477 col\[4\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[4\].zbuf_bot_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_2403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_234 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_212 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_223 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_201 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_433_ col\[7\].zbuf_bot_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[256] sky130_fd_sc_hd__buf_2
XANTENNA_256 col\[0\].genblk1.tbuf_spine_ow_I\[18\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_245 col\[0\].genblk1.tbuf_spine_ow_I\[17\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_267 col\[0\].genblk1.tbuf_spine_ow_I\[2\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_278 col\[0\].genblk1.tbuf_spine_ow_I\[3\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_289 col\[0\].genblk1.tbuf_spine_ow_I\[9\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_364_ col\[5\].zbuf_bot_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[187] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_295_ col\[3\].zbuf_bot_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[118] sky130_fd_sc_hd__buf_2
Xcol\[6\].zbuf_bot_iw_I\[3\].genblk1.cell0_I net488 col\[6\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[6\].zbuf_bot_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_2490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].genblk1.mux4_I\[13\].cell0_I net259 net285 net311 net338 net471 net457 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[13\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_2_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_2322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].zbuf_top_iw_I\[7\].genblk1.cell0_I net479 net430 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[7\].z sky130_fd_sc_hd__and2_1
X_080_ _020_ vssd1 vssd1 vccd1 vccd1 col\[3\].zbuf_bot_ena_I.e sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_2277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_416_ col\[6\].zbuf_top_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[239] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_top_iw_I\[2\].genblk1.cell0_I net489 net426 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[2\].z sky130_fd_sc_hd__and2_1
X_347_ col\[4\].zbuf_top_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[170] sky130_fd_sc_hd__buf_2
X_278_ col\[2\].zbuf_top_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[101] sky130_fd_sc_hd__buf_2
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[4\].genblk1.mux4_I\[4\].cell0_I net141 net169 net195 net221 net468 net454 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[4\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_7_2929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_2528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xzbuf_bus_iw_I\[15\].genblk1.cell0_I net24 net515 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[15\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_201_ col\[0\].zbuf_top_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[24] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_063_ net467 net453 col\[0\].genblk1.tbuf_row_ena_I.t zbuf_bus_ena_I.z vssd1 vssd1
+ vccd1 vccd1 _010_ sky130_fd_sc_hd__and4bb_2
Xcol\[2\].genblk1.tbuf_spine_ow_I\[9\].cell0_I col\[2\].genblk1.mux4_I\[9\].x net442
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[9\].z sky130_fd_sc_hd__ebufn_8
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[0\].genblk1.mux4_I\[2\].cell0_I net257 net223 net364 net390 net463 net449 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[2\].x sky130_fd_sc_hd__mux4_2
Xfanout490 col\[0\].zbuf_bot_iw_I\[2\].a vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_2041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_2085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[0\].zbuf_bot_iw_I\[12\].genblk1.cell0_I net503 col\[0\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[0\].zbuf_bot_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_2737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_2658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_2269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xzbuf_bus_iw_I\[2\].genblk1.cell0_I net10 net514 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[2\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_0_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_2934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[7\].zbuf_top_iw_I\[5\].genblk1.cell0_I net484 net419 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_2770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_2809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_2656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[6\].genblk1.mux4_I\[7\].cell0_I net251 net278 net305 net331 net473 net459 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[7\].x sky130_fd_sc_hd__mux4_1
Xinput300 um_ow[339] vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput311 um_ow[349] vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput333 um_ow[369] vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput344 um_ow[379] vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput322 um_ow[359] vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput388 um_ow[72] vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__clkbuf_1
Xinput355 um_ow[42] vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__clkbuf_2
Xinput377 um_ow[62] vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__clkbuf_1
Xinput366 um_ow[52] vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_1
Xinput399 um_ow[82] vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].zbuf_bot_iw_I\[11\].genblk1.cell0_I net505 col\[2\].zbuf_bot_ena_I.e vssd1
+ vssd1 vccd1 vccd1 col\[2\].zbuf_bot_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_2099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 col\[0\].genblk1.tbuf_spine_ow_I\[0\].z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_2420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[2\].genblk1.mux4_I\[5\].cell0_I net37 net63 net89 net116 net466 net452 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[5\].x sky130_fd_sc_hd__mux4_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_380_ col\[5\].zbuf_top_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[203] sky130_fd_sc_hd__buf_2
XFILLER_0_3_2228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[0\].genblk1.tbuf_spine_ow_I\[13\].cell0_I col\[0\].genblk1.mux4_I\[13\].x net445
+ vssd1 vssd1 vccd1 vccd1 col\[0\].genblk1.tbuf_spine_ow_I\[13\].z sky130_fd_sc_hd__ebufn_8
Xtbuf_spine_ow_I\[11\].cell0_I col\[0\].genblk1.tbuf_spine_ow_I\[11\].z net512 vssd1
+ vssd1 vccd1 vccd1 tbuf_spine_ow_I\[11\].z sky130_fd_sc_hd__ebufn_1
Xinput130 um_ow[186] vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__clkbuf_1
Xinput141 um_ow[196] vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__clkbuf_1
Xinput152 um_ow[205] vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__clkbuf_1
Xinput163 um_ow[215] vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_1
Xinput174 um_ow[225] vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_1
Xinput185 um_ow[235] vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_1
Xinput196 um_ow[245] vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

