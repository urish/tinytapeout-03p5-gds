magic
tech sky130A
magscale 1 2
timestamp 1685641958
<< obsli1 >>
rect 1104 1071 271492 9809
<< obsm1 >>
rect 842 8 272214 10872
<< obsm2 >>
rect 846 2 272210 10878
<< metal3 >>
rect 270554 9558 272504 9618
rect 272210 9422 272504 9482
rect 268070 9286 272504 9346
rect 268806 9150 272504 9210
rect 268714 9014 272504 9074
rect 272026 8878 272504 8938
rect 271830 8742 272504 8802
rect 272304 8606 272504 8666
rect 268346 8470 272504 8530
rect 268070 8334 272504 8394
rect 272014 8198 272504 8258
rect 272210 8062 272504 8122
rect 272210 7926 272504 7986
rect 264942 7790 272504 7850
rect 271842 7654 272504 7714
rect 271830 7518 272504 7578
rect 272026 7382 272504 7442
rect 262366 7246 272504 7306
rect 263286 7110 272504 7170
rect 267978 6974 272504 7034
rect 267978 6838 272504 6898
rect 271014 6702 272504 6762
rect 272118 6566 272504 6626
rect 271934 6430 272504 6490
rect 271382 6294 272504 6354
rect 270542 6158 272504 6218
rect 271750 6022 272504 6082
rect 271198 5886 272504 5946
rect 270910 5750 272504 5810
rect 270726 5614 272504 5674
rect 271842 5478 272504 5538
rect 271842 5342 272504 5402
rect 269082 5206 272504 5266
rect 268530 5070 272504 5130
rect 272026 4934 272504 4994
rect 268990 4798 272504 4858
rect 268346 4662 272504 4722
rect 272304 4526 272504 4586
rect 271830 4390 272504 4450
rect 271842 4254 272504 4314
rect 271830 4118 272504 4178
rect 272014 3982 272504 4042
rect 272210 3846 272504 3906
rect 268070 3710 272504 3770
rect 272210 3574 272504 3634
rect 272014 3438 272504 3498
rect 271830 3302 272504 3362
rect 271842 3166 272504 3226
rect 267978 3030 272504 3090
rect 258766 2894 272504 2954
rect 271290 2758 272504 2818
rect 267978 2622 272504 2682
rect 268438 2486 272504 2546
rect 248474 2350 272504 2410
rect 271830 2214 272504 2274
rect 272026 2078 272504 2138
rect 272118 1942 272504 2002
rect 268898 1806 272504 1866
rect 269622 1670 272504 1730
rect 272210 1534 272504 1594
rect 258778 1398 272504 1458
rect 272026 1262 272504 1322
rect 271830 1126 272504 1186
rect 272198 990 272504 1050
<< obsm3 >>
rect 750 9698 272258 10573
rect 750 9478 270474 9698
rect 750 9426 272130 9478
rect 750 9206 267990 9426
rect 750 9154 268726 9206
rect 750 8934 268634 9154
rect 750 8882 271946 8934
rect 750 8662 271750 8882
rect 750 8610 272224 8662
rect 750 8474 268266 8610
rect 750 8254 267990 8474
rect 750 8118 271934 8254
rect 750 7930 272130 8118
rect 750 7710 264862 7930
rect 750 7658 271762 7710
rect 750 7438 271750 7658
rect 750 7386 271946 7438
rect 750 7166 262286 7386
rect 750 7030 263206 7166
rect 750 6758 267898 7030
rect 750 6622 270934 6758
rect 750 6570 272038 6622
rect 750 6434 271854 6570
rect 750 6298 271302 6434
rect 750 6078 270462 6298
rect 750 6026 271670 6078
rect 750 5890 271118 6026
rect 750 5754 270830 5890
rect 750 5534 270646 5754
rect 750 5346 271762 5534
rect 750 5210 269002 5346
rect 750 4990 268450 5210
rect 750 4938 271946 4990
rect 750 4802 268910 4938
rect 750 4582 268266 4802
rect 750 4530 272224 4582
rect 750 4310 271750 4530
rect 750 4258 271762 4310
rect 750 4038 271750 4258
rect 750 3902 271934 4038
rect 750 3850 272130 3902
rect 750 3630 267990 3850
rect 750 3578 272130 3630
rect 750 3442 271934 3578
rect 750 3222 271750 3442
rect 750 3170 271762 3222
rect 750 3034 267898 3170
rect 750 2814 258686 3034
rect 750 2762 271210 2814
rect 750 2542 267898 2762
rect 750 2490 268358 2542
rect 750 2270 248394 2490
rect 750 2134 271750 2270
rect 750 1998 271946 2134
rect 750 1946 272038 1998
rect 750 1726 268818 1946
rect 750 1590 269542 1726
rect 750 1538 272130 1590
rect 750 1318 258698 1538
rect 750 1266 271946 1318
rect 750 1046 271750 1266
rect 750 910 272118 1046
rect 750 35 272258 910
<< metal4 >>
rect 798 9212 858 10880
rect 1534 10164 1594 10880
rect 2270 10164 2330 10880
rect 3006 9892 3066 10880
rect 3742 10164 3802 10880
rect 4478 10164 4538 10880
rect 5214 10164 5274 10880
rect 5950 10164 6010 10880
rect 6686 10164 6746 10880
rect 7422 10164 7482 10880
rect 8158 9892 8218 10880
rect 8894 10164 8954 10880
rect 9630 10164 9690 10880
rect 10366 10164 10426 10880
rect 11102 10164 11162 10880
rect 11838 10164 11898 10880
rect 12574 10164 12634 10880
rect 13310 9892 13370 10880
rect 14046 10164 14106 10880
rect 14782 10164 14842 10880
rect 15518 10164 15578 10880
rect 16254 10164 16314 10880
rect 16990 10164 17050 10880
rect 17726 10164 17786 10880
rect 18462 10164 18522 10880
rect 19198 6900 19258 10880
rect 19934 9892 19994 10880
rect 20670 8396 20730 10880
rect 21406 8668 21466 10880
rect 22142 8940 22202 10880
rect 22878 8396 22938 10880
rect 23614 8396 23674 10880
rect 24350 9212 24410 10880
rect 25086 8396 25146 10880
rect 25822 9756 25882 10880
rect 26558 9756 26618 10880
rect 27294 8668 27354 10880
rect 28030 8668 28090 10880
rect 28766 8668 28826 10880
rect 29502 9756 29562 10880
rect 30238 9756 30298 10880
rect 30974 8668 31034 10880
rect 31710 10300 31770 10880
rect 32446 9212 32506 10880
rect 34930 10300 34990 10880
rect 35666 10300 35726 10880
rect 36402 10300 36462 10880
rect 37138 10300 37198 10880
rect 37874 10300 37934 10880
rect 38610 10300 38670 10880
rect 39346 10300 39406 10880
rect 40082 10300 40142 10880
rect 40818 10300 40878 10880
rect 41554 10300 41614 10880
rect 42290 10300 42350 10880
rect 43026 10300 43086 10880
rect 43762 10300 43822 10880
rect 44498 10300 44558 10880
rect 45234 10300 45294 10880
rect 45970 10300 46030 10880
rect 46706 10300 46766 10880
rect 47442 10300 47502 10880
rect 48178 10300 48238 10880
rect 48914 10300 48974 10880
rect 49650 10300 49710 10880
rect 50386 10300 50446 10880
rect 51122 10300 51182 10880
rect 51858 10300 51918 10880
rect 52594 10572 52654 10880
rect 53330 10300 53390 10880
rect 54066 10300 54126 10880
rect 54802 10300 54862 10880
rect 55538 10300 55598 10880
rect 56274 10300 56334 10880
rect 57010 10300 57070 10880
rect 57746 10300 57806 10880
rect 58482 10300 58542 10880
rect 59218 10300 59278 10880
rect 59954 10300 60014 10880
rect 60690 10300 60750 10880
rect 61426 10300 61486 10880
rect 62162 10300 62222 10880
rect 62898 10300 62958 10880
rect 63634 10300 63694 10880
rect 64370 10300 64430 10880
rect 65106 10300 65166 10880
rect 65842 10300 65902 10880
rect 66578 10300 66638 10880
rect 798 0 858 2756
rect 1534 0 1594 988
rect 2270 0 2330 580
rect 3006 0 3066 716
rect 3742 0 3802 988
rect 4478 0 4538 1260
rect 5214 0 5274 988
rect 5950 0 6010 716
rect 6686 0 6746 1260
rect 7422 0 7482 988
rect 8158 0 8218 444
rect 8894 0 8954 308
rect 9630 0 9690 988
rect 10366 0 10426 716
rect 11102 0 11162 716
rect 11838 0 11898 988
rect 12574 0 12634 988
rect 13310 0 13370 580
rect 14046 0 14106 988
rect 14782 0 14842 1260
rect 15518 0 15578 988
rect 16254 0 16314 716
rect 16990 0 17050 716
rect 17726 0 17786 988
rect 18462 0 18522 308
rect 19198 0 19258 2756
rect 19934 0 19994 1532
rect 20670 0 20730 1396
rect 21406 0 21466 580
rect 22142 0 22202 1668
rect 22878 0 22938 2756
rect 23614 0 23674 1260
rect 24350 0 24410 1260
rect 25086 0 25146 2756
rect 25822 0 25882 1260
rect 26558 0 26618 1260
rect 27294 0 27354 2756
rect 28030 0 28090 580
rect 28766 0 28826 308
rect 29502 0 29562 1124
rect 30238 0 30298 580
rect 30974 0 31034 580
rect 31710 0 31770 580
rect 32446 0 32506 1532
rect 34742 1040 35062 9840
rect 68540 1040 68860 9840
rect 69062 9620 69122 10880
rect 69798 9892 69858 10880
rect 70534 9620 70594 10880
rect 71270 10164 71330 10880
rect 72006 10436 72066 10880
rect 72742 9620 72802 10880
rect 73478 9076 73538 10880
rect 74214 9620 74274 10880
rect 74950 9076 75010 10880
rect 75686 9620 75746 10880
rect 76422 9620 76482 10880
rect 77158 9892 77218 10880
rect 77894 9620 77954 10880
rect 78630 9892 78690 10880
rect 79366 10164 79426 10880
rect 80102 9620 80162 10880
rect 80838 9892 80898 10880
rect 81574 10572 81634 10880
rect 82310 10572 82370 10880
rect 83046 10164 83106 10880
rect 83782 10164 83842 10880
rect 84518 10164 84578 10880
rect 85254 10164 85314 10880
rect 85990 9892 86050 10880
rect 86726 10572 86786 10880
rect 87462 8668 87522 10880
rect 88198 9212 88258 10880
rect 88934 8124 88994 10880
rect 89670 10300 89730 10880
rect 90406 8668 90466 10880
rect 91142 10028 91202 10880
rect 91878 9212 91938 10880
rect 92614 9756 92674 10880
rect 93350 9756 93410 10880
rect 94086 8668 94146 10880
rect 94822 8668 94882 10880
rect 95558 9756 95618 10880
rect 96294 9756 96354 10880
rect 97030 8668 97090 10880
rect 97766 8668 97826 10880
rect 98502 9756 98562 10880
rect 99238 8668 99298 10880
rect 99974 9756 100034 10880
rect 100710 9212 100770 10880
rect 103194 10300 103254 10880
rect 103930 10300 103990 10880
rect 104666 10300 104726 10880
rect 105402 10300 105462 10880
rect 106138 10300 106198 10880
rect 106874 10300 106934 10880
rect 107610 10300 107670 10880
rect 108346 10300 108406 10880
rect 109082 10300 109142 10880
rect 109818 10300 109878 10880
rect 110554 10300 110614 10880
rect 111290 10300 111350 10880
rect 112026 10300 112086 10880
rect 112762 10300 112822 10880
rect 113498 10300 113558 10880
rect 114234 10300 114294 10880
rect 114970 10300 115030 10880
rect 115706 10300 115766 10880
rect 116442 10300 116502 10880
rect 117178 10300 117238 10880
rect 117914 10300 117974 10880
rect 118650 10300 118710 10880
rect 119386 10300 119446 10880
rect 120122 10300 120182 10880
rect 120858 10300 120918 10880
rect 121594 10300 121654 10880
rect 122330 10300 122390 10880
rect 123066 10300 123126 10880
rect 123802 10300 123862 10880
rect 124538 10300 124598 10880
rect 125274 10436 125334 10880
rect 126010 10300 126070 10880
rect 126746 10300 126806 10880
rect 127482 10300 127542 10880
rect 128218 10300 128278 10880
rect 128954 10300 129014 10880
rect 129690 10300 129750 10880
rect 130426 10300 130486 10880
rect 131162 10300 131222 10880
rect 131898 10300 131958 10880
rect 132634 10300 132694 10880
rect 133370 10300 133430 10880
rect 134106 10300 134166 10880
rect 134842 10300 134902 10880
rect 34930 0 34990 580
rect 35666 0 35726 580
rect 36402 0 36462 580
rect 37138 0 37198 580
rect 37874 0 37934 580
rect 38610 0 38670 580
rect 39346 0 39406 308
rect 40082 0 40142 580
rect 40818 0 40878 580
rect 41554 0 41614 580
rect 42290 0 42350 580
rect 43026 0 43086 580
rect 43762 0 43822 580
rect 44498 0 44558 580
rect 45234 0 45294 580
rect 45970 0 46030 580
rect 46706 0 46766 580
rect 47442 0 47502 580
rect 48178 0 48238 580
rect 48914 0 48974 580
rect 49650 0 49710 580
rect 50386 0 50446 580
rect 51122 0 51182 580
rect 51858 0 51918 580
rect 52594 0 52654 308
rect 53330 0 53390 580
rect 54066 0 54126 580
rect 54802 0 54862 370
rect 55538 0 55598 444
rect 56274 0 56334 444
rect 57010 0 57070 444
rect 57746 0 57806 370
rect 58482 0 58542 444
rect 59218 0 59278 370
rect 59954 0 60014 444
rect 60690 0 60750 444
rect 61426 0 61486 444
rect 62162 0 62222 444
rect 62898 0 62958 444
rect 63634 0 63694 308
rect 64370 0 64430 308
rect 65106 0 65166 308
rect 65842 0 65902 444
rect 66578 0 66638 444
rect 69062 0 69122 852
rect 69798 0 69858 852
rect 70534 0 70594 852
rect 71270 0 71330 988
rect 72006 0 72066 988
rect 72742 0 72802 852
rect 73478 0 73538 988
rect 74214 0 74274 852
rect 74950 0 75010 852
rect 75686 0 75746 988
rect 76422 0 76482 1260
rect 77158 0 77218 988
rect 77894 0 77954 852
rect 78630 0 78690 1260
rect 79366 0 79426 988
rect 80102 0 80162 852
rect 80838 0 80898 988
rect 81574 0 81634 1260
rect 82310 0 82370 988
rect 83046 0 83106 852
rect 83782 0 83842 1260
rect 84518 0 84578 988
rect 85254 0 85314 308
rect 85990 0 86050 988
rect 86726 0 86786 852
rect 87462 0 87522 444
rect 88198 0 88258 1396
rect 88934 0 88994 1260
rect 89670 0 89730 370
rect 90406 0 90466 1260
rect 91142 0 91202 1532
rect 91878 0 91938 1260
rect 92614 0 92674 580
rect 93350 0 93410 1260
rect 94086 0 94146 3028
rect 94822 0 94882 580
rect 95558 0 95618 2756
rect 96294 0 96354 1532
rect 97030 0 97090 2756
rect 97766 0 97826 3708
rect 98502 0 98562 1532
rect 99238 0 99298 852
rect 99974 0 100034 580
rect 100710 0 100770 3164
rect 102339 1040 102659 9840
rect 136137 1040 136457 9840
rect 137326 9620 137386 10880
rect 138062 10300 138122 10880
rect 138798 10164 138858 10880
rect 139534 9892 139594 10880
rect 140270 10164 140330 10880
rect 141006 10164 141066 10880
rect 141742 10164 141802 10880
rect 142478 10300 142538 10880
rect 143214 10164 143274 10880
rect 143950 10164 144010 10880
rect 144686 9892 144746 10880
rect 145422 10164 145482 10880
rect 146158 10164 146218 10880
rect 146894 10164 146954 10880
rect 147630 10572 147690 10880
rect 148366 10300 148426 10880
rect 149102 10164 149162 10880
rect 149838 9892 149898 10880
rect 150574 10164 150634 10880
rect 151310 10164 151370 10880
rect 152046 10164 152106 10880
rect 152782 10164 152842 10880
rect 153518 10164 153578 10880
rect 154254 10436 154314 10880
rect 154990 9892 155050 10880
rect 155726 8668 155786 10880
rect 156462 9484 156522 10880
rect 157198 8396 157258 10880
rect 157934 8124 157994 10880
rect 158670 8396 158730 10880
rect 159406 8124 159466 10880
rect 160142 8396 160202 10880
rect 160878 8124 160938 10880
rect 161614 8396 161674 10880
rect 162350 7852 162410 10880
rect 163086 8396 163146 10880
rect 163822 8124 163882 10880
rect 164558 8396 164618 10880
rect 165294 8124 165354 10880
rect 166030 8396 166090 10880
rect 166766 8396 166826 10880
rect 167502 9756 167562 10880
rect 168238 9212 168298 10880
rect 168974 9756 169034 10880
rect 171458 10300 171518 10880
rect 172194 10572 172254 10880
rect 172930 10436 172990 10880
rect 173666 10300 173726 10880
rect 174402 10300 174462 10880
rect 175138 10300 175198 10880
rect 175874 10300 175934 10880
rect 176610 10300 176670 10880
rect 177346 10300 177406 10880
rect 178082 10300 178142 10880
rect 178818 10300 178878 10880
rect 179554 10572 179614 10880
rect 180290 10300 180350 10880
rect 181026 10436 181086 10880
rect 181762 10300 181822 10880
rect 182498 10300 182558 10880
rect 183234 10300 183294 10880
rect 183970 10300 184030 10880
rect 184706 10300 184766 10880
rect 185442 10300 185502 10880
rect 186178 10300 186238 10880
rect 186914 10300 186974 10880
rect 187650 10300 187710 10880
rect 188386 10300 188446 10880
rect 189122 10300 189182 10880
rect 189858 10300 189918 10880
rect 190594 10436 190654 10880
rect 191330 10300 191390 10880
rect 192066 10300 192126 10880
rect 192802 10436 192862 10880
rect 193538 10300 193598 10880
rect 194274 10300 194334 10880
rect 195010 10300 195070 10880
rect 195746 10300 195806 10880
rect 196482 10300 196542 10880
rect 197218 10300 197278 10880
rect 197954 10300 198014 10880
rect 198690 10300 198750 10880
rect 199426 10300 199486 10880
rect 200162 10300 200222 10880
rect 200898 10300 200958 10880
rect 201634 10300 201694 10880
rect 202370 10436 202430 10880
rect 203106 10300 203166 10880
rect 205590 10300 205650 10880
rect 206326 10164 206386 10880
rect 207062 10164 207122 10880
rect 207798 10572 207858 10880
rect 208534 10164 208594 10880
rect 209270 10164 209330 10880
rect 210006 10436 210066 10880
rect 210742 10164 210802 10880
rect 103194 0 103254 370
rect 103930 0 103990 370
rect 104666 0 104726 370
rect 105402 0 105462 370
rect 106138 0 106198 370
rect 106874 0 106934 370
rect 107610 0 107670 370
rect 108346 0 108406 370
rect 109082 0 109142 370
rect 109818 0 109878 370
rect 110554 0 110614 370
rect 111290 0 111350 370
rect 112026 0 112086 370
rect 112762 0 112822 370
rect 113498 0 113558 370
rect 114234 0 114294 370
rect 114970 0 115030 370
rect 115706 0 115766 370
rect 116442 0 116502 370
rect 117178 0 117238 370
rect 117914 0 117974 444
rect 118650 0 118710 444
rect 119386 0 119446 444
rect 120122 0 120182 444
rect 120858 0 120918 444
rect 121594 0 121654 444
rect 122330 0 122390 444
rect 123066 0 123126 444
rect 123802 0 123862 370
rect 124538 0 124598 580
rect 125274 0 125334 580
rect 126010 0 126070 580
rect 126746 0 126806 370
rect 127482 0 127542 444
rect 128218 0 128278 370
rect 128954 0 129014 580
rect 129690 0 129750 308
rect 130426 0 130486 580
rect 131162 0 131222 580
rect 131898 0 131958 308
rect 132634 0 132694 308
rect 133370 0 133430 370
rect 134106 0 134166 580
rect 134842 0 134902 370
rect 137326 0 137386 1396
rect 138062 0 138122 580
rect 138798 0 138858 716
rect 139534 0 139594 988
rect 140270 0 140330 1804
rect 141006 0 141066 1396
rect 141742 0 141802 716
rect 142478 0 142538 716
rect 143214 0 143274 580
rect 143950 0 144010 444
rect 144686 0 144746 3164
rect 145422 0 145482 2756
rect 146158 0 146218 716
rect 146894 0 146954 308
rect 147630 0 147690 580
rect 148366 0 148426 716
rect 149102 0 149162 2892
rect 149838 0 149898 716
rect 150574 0 150634 1396
rect 151310 0 151370 580
rect 152046 0 152106 1396
rect 152782 0 152842 1260
rect 153518 0 153578 2892
rect 154254 0 154314 3300
rect 154990 0 155050 2892
rect 155726 0 155786 1396
rect 156462 0 156522 2756
rect 157198 0 157258 1396
rect 157934 0 157994 1260
rect 158670 0 158730 1124
rect 159406 0 159466 580
rect 160142 0 160202 1124
rect 160878 0 160938 308
rect 161614 0 161674 1124
rect 162350 0 162410 580
rect 163086 0 163146 580
rect 163822 0 163882 1124
rect 164558 0 164618 580
rect 165294 0 165354 1124
rect 166030 0 166090 1124
rect 166766 0 166826 1124
rect 167502 0 167562 308
rect 168238 0 168298 1396
rect 169936 1040 170256 9840
rect 203734 1040 204054 9840
rect 211478 9892 211538 10880
rect 212214 10164 212274 10880
rect 212950 10572 213010 10880
rect 213686 10164 213746 10880
rect 214422 10164 214482 10880
rect 215158 9620 215218 10880
rect 215894 10164 215954 10880
rect 216630 9892 216690 10880
rect 217366 10164 217426 10880
rect 218102 10572 218162 10880
rect 218838 10164 218898 10880
rect 219574 10164 219634 10880
rect 220310 10300 220370 10880
rect 221046 10436 221106 10880
rect 221782 9892 221842 10880
rect 222518 10164 222578 10880
rect 223254 10164 223314 10880
rect 223990 9484 224050 10880
rect 224726 8668 224786 10880
rect 225462 8668 225522 10880
rect 226198 8668 226258 10880
rect 226934 8668 226994 10880
rect 227670 9484 227730 10880
rect 228406 9484 228466 10880
rect 229142 8668 229202 10880
rect 229878 9484 229938 10880
rect 230614 8668 230674 10880
rect 231350 8668 231410 10880
rect 232086 9484 232146 10880
rect 232822 8668 232882 10880
rect 233558 9484 233618 10880
rect 234294 8668 234354 10880
rect 235030 8396 235090 10880
rect 235766 9484 235826 10880
rect 236502 9212 236562 10880
rect 237238 8668 237298 10880
rect 239722 10300 239782 10880
rect 240458 10300 240518 10880
rect 241194 10300 241254 10880
rect 241930 10300 241990 10880
rect 242666 10300 242726 10880
rect 243402 10300 243462 10880
rect 244138 10300 244198 10880
rect 244874 10300 244934 10880
rect 245610 10436 245670 10880
rect 246346 10300 246406 10880
rect 247082 10300 247142 10880
rect 247818 10300 247878 10880
rect 248554 10300 248614 10880
rect 249290 10300 249350 10880
rect 250026 10300 250086 10880
rect 250762 10300 250822 10880
rect 251498 10300 251558 10880
rect 252234 10300 252294 10880
rect 252970 10436 253030 10880
rect 253706 10300 253766 10880
rect 254442 10300 254502 10880
rect 255178 10300 255238 10880
rect 255914 10300 255974 10880
rect 256650 10300 256710 10880
rect 257386 10300 257446 10880
rect 258122 10300 258182 10880
rect 258858 10300 258918 10880
rect 259594 10300 259654 10880
rect 260330 10300 260390 10880
rect 261066 10436 261126 10880
rect 261802 10300 261862 10880
rect 262538 10300 262598 10880
rect 263274 10300 263334 10880
rect 264010 10300 264070 10880
rect 264746 10238 264806 10880
rect 265482 10436 265542 10880
rect 266218 10300 266278 10880
rect 266954 10238 267014 10880
rect 267690 10238 267750 10880
rect 268426 10238 268486 10880
rect 269162 10238 269222 10880
rect 269898 10238 269958 10880
rect 270634 10238 270694 10880
rect 271370 10238 271430 10880
rect 168974 0 169034 580
rect 171458 0 171518 580
rect 172194 0 172254 580
rect 172930 0 172990 580
rect 173666 0 173726 580
rect 174402 0 174462 580
rect 175138 0 175198 580
rect 175874 0 175934 444
rect 176610 0 176670 580
rect 177346 0 177406 580
rect 178082 0 178142 580
rect 178818 0 178878 580
rect 179554 0 179614 580
rect 180290 0 180350 580
rect 181026 0 181086 308
rect 181762 0 181822 444
rect 182498 0 182558 444
rect 183234 0 183294 444
rect 183970 0 184030 444
rect 184706 0 184766 444
rect 185442 0 185502 444
rect 186178 0 186238 370
rect 186914 0 186974 444
rect 187650 0 187710 444
rect 188386 0 188446 444
rect 189122 0 189182 444
rect 189858 0 189918 370
rect 190594 0 190654 444
rect 191330 0 191390 370
rect 192066 0 192126 308
rect 192802 0 192862 444
rect 193538 0 193598 444
rect 194274 0 194334 370
rect 195010 0 195070 444
rect 195746 0 195806 370
rect 196482 0 196542 444
rect 197218 0 197278 370
rect 197954 0 198014 370
rect 198690 0 198750 444
rect 199426 0 199486 370
rect 200162 0 200222 444
rect 200898 0 200958 370
rect 201634 0 201694 370
rect 202370 0 202430 444
rect 203106 0 203166 444
rect 205590 0 205650 852
rect 206326 0 206386 852
rect 207062 0 207122 852
rect 207798 0 207858 308
rect 208534 0 208594 852
rect 209270 0 209330 444
rect 210006 0 210066 1396
rect 210742 0 210802 2756
rect 211478 0 211538 3028
rect 212214 0 212274 1804
rect 212950 0 213010 308
rect 213686 0 213746 444
rect 214422 0 214482 308
rect 215158 0 215218 3980
rect 215894 0 215954 716
rect 216630 0 216690 2892
rect 217366 0 217426 3164
rect 218102 0 218162 1396
rect 218838 0 218898 3708
rect 219574 0 219634 1396
rect 220310 0 220370 308
rect 221046 0 221106 3164
rect 221782 0 221842 580
rect 222518 0 222578 1396
rect 223254 0 223314 3708
rect 223990 0 224050 1124
rect 224726 0 224786 716
rect 225462 0 225522 1124
rect 226198 0 226258 1396
rect 226934 0 226994 580
rect 227670 0 227730 1124
rect 228406 0 228466 580
rect 229142 0 229202 580
rect 229878 0 229938 1124
rect 230614 0 230674 1124
rect 231350 0 231410 580
rect 232086 0 232146 1124
rect 232822 0 232882 1124
rect 233558 0 233618 580
rect 234294 0 234354 580
rect 235030 0 235090 1124
rect 235766 0 235826 580
rect 236502 0 236562 1124
rect 237238 0 237298 1532
rect 237533 1040 237853 9840
rect 271331 1040 271651 9840
rect 239722 0 239782 580
rect 240458 0 240518 580
rect 241194 0 241254 580
rect 241930 0 241990 580
rect 242666 0 242726 370
rect 243402 0 243462 580
rect 244138 0 244198 580
rect 244874 0 244934 580
rect 245610 0 245670 370
rect 246346 0 246406 642
rect 247082 0 247142 580
rect 247818 0 247878 580
rect 248554 0 248614 370
rect 249290 0 249350 370
rect 250026 0 250086 580
rect 250762 0 250822 642
rect 251498 0 251558 370
rect 252234 0 252294 370
rect 252970 0 253030 444
rect 253706 0 253766 308
rect 254442 0 254502 580
rect 255178 0 255238 580
rect 255914 0 255974 642
rect 256650 0 256710 370
rect 257386 0 257446 370
rect 258122 0 258182 580
rect 258858 0 258918 642
rect 259594 0 259654 642
rect 260330 0 260390 642
rect 261066 0 261126 580
rect 261802 0 261862 642
rect 262538 0 262598 580
rect 263274 0 263334 580
rect 264010 0 264070 580
rect 264746 0 264806 580
rect 265482 0 265542 580
rect 266218 0 266278 580
rect 266954 0 267014 580
rect 267690 0 267750 580
rect 268426 0 268486 580
rect 269162 0 269222 580
rect 269898 0 269958 308
rect 270634 0 270694 580
rect 271370 0 271430 642
<< obsm4 >>
rect 938 10084 1454 10573
rect 1674 10084 2190 10573
rect 2410 10084 2926 10573
rect 938 9812 2926 10084
rect 3146 10084 3662 10573
rect 3882 10084 4398 10573
rect 4618 10084 5134 10573
rect 5354 10084 5870 10573
rect 6090 10084 6606 10573
rect 6826 10084 7342 10573
rect 7562 10084 8078 10573
rect 3146 9812 8078 10084
rect 8298 10084 8814 10573
rect 9034 10084 9550 10573
rect 9770 10084 10286 10573
rect 10506 10084 11022 10573
rect 11242 10084 11758 10573
rect 11978 10084 12494 10573
rect 12714 10084 13230 10573
rect 8298 9812 13230 10084
rect 13450 10084 13966 10573
rect 14186 10084 14702 10573
rect 14922 10084 15438 10573
rect 15658 10084 16174 10573
rect 16394 10084 16910 10573
rect 17130 10084 17646 10573
rect 17866 10084 18382 10573
rect 18602 10084 19118 10573
rect 13450 9812 19118 10084
rect 938 9132 19118 9812
rect 795 6820 19118 9132
rect 19338 9812 19854 10573
rect 20074 9812 20590 10573
rect 19338 8316 20590 9812
rect 20810 8588 21326 10573
rect 21546 8860 22062 10573
rect 22282 8860 22798 10573
rect 21546 8588 22798 8860
rect 20810 8316 22798 8588
rect 23018 8316 23534 10573
rect 23754 9132 24270 10573
rect 24490 9132 25006 10573
rect 23754 8316 25006 9132
rect 25226 9676 25742 10573
rect 25962 9676 26478 10573
rect 26698 9676 27214 10573
rect 25226 8588 27214 9676
rect 27434 8588 27950 10573
rect 28170 8588 28686 10573
rect 28906 9676 29422 10573
rect 29642 9676 30158 10573
rect 30378 9676 30894 10573
rect 28906 8588 30894 9676
rect 31114 10220 31630 10573
rect 31850 10220 32366 10573
rect 31114 9132 32366 10220
rect 32586 10220 34850 10573
rect 35070 10220 35586 10573
rect 35806 10220 36322 10573
rect 36542 10220 37058 10573
rect 37278 10220 37794 10573
rect 38014 10220 38530 10573
rect 38750 10220 39266 10573
rect 39486 10220 40002 10573
rect 40222 10220 40738 10573
rect 40958 10220 41474 10573
rect 41694 10220 42210 10573
rect 42430 10220 42946 10573
rect 43166 10220 43682 10573
rect 43902 10220 44418 10573
rect 44638 10220 45154 10573
rect 45374 10220 45890 10573
rect 46110 10220 46626 10573
rect 46846 10220 47362 10573
rect 47582 10220 48098 10573
rect 48318 10220 48834 10573
rect 49054 10220 49570 10573
rect 49790 10220 50306 10573
rect 50526 10220 51042 10573
rect 51262 10220 51778 10573
rect 51998 10492 52514 10573
rect 52734 10492 53250 10573
rect 51998 10220 53250 10492
rect 53470 10220 53986 10573
rect 54206 10220 54722 10573
rect 54942 10220 55458 10573
rect 55678 10220 56194 10573
rect 56414 10220 56930 10573
rect 57150 10220 57666 10573
rect 57886 10220 58402 10573
rect 58622 10220 59138 10573
rect 59358 10220 59874 10573
rect 60094 10220 60610 10573
rect 60830 10220 61346 10573
rect 61566 10220 62082 10573
rect 62302 10220 62818 10573
rect 63038 10220 63554 10573
rect 63774 10220 64290 10573
rect 64510 10220 65026 10573
rect 65246 10220 65762 10573
rect 65982 10220 66498 10573
rect 66718 10220 68982 10573
rect 32586 9920 68982 10220
rect 32586 9132 34662 9920
rect 31114 8588 34662 9132
rect 25226 8316 34662 8588
rect 19338 6820 34662 8316
rect 795 2836 34662 6820
rect 938 1340 19118 2836
rect 938 1068 4398 1340
rect 938 171 1454 1068
rect 1674 796 3662 1068
rect 1674 660 2926 796
rect 1674 171 2190 660
rect 2410 171 2926 660
rect 3146 171 3662 796
rect 3882 171 4398 1068
rect 4618 1068 6606 1340
rect 4618 171 5134 1068
rect 5354 796 6606 1068
rect 5354 171 5870 796
rect 6090 171 6606 796
rect 6826 1068 14702 1340
rect 6826 171 7342 1068
rect 7562 524 9550 1068
rect 7562 171 8078 524
rect 8298 388 9550 524
rect 8298 171 8814 388
rect 9034 171 9550 388
rect 9770 796 11758 1068
rect 9770 171 10286 796
rect 10506 171 11022 796
rect 11242 171 11758 796
rect 11978 171 12494 1068
rect 12714 660 13966 1068
rect 12714 171 13230 660
rect 13450 171 13966 660
rect 14186 171 14702 1068
rect 14922 1068 19118 1340
rect 14922 171 15438 1068
rect 15658 796 17646 1068
rect 15658 171 16174 796
rect 16394 171 16910 796
rect 17130 171 17646 796
rect 17866 388 19118 1068
rect 17866 171 18382 388
rect 18602 171 19118 388
rect 19338 1748 22798 2836
rect 19338 1612 22062 1748
rect 19338 171 19854 1612
rect 20074 1476 22062 1612
rect 20074 171 20590 1476
rect 20810 660 22062 1476
rect 20810 171 21326 660
rect 21546 171 22062 660
rect 22282 171 22798 1748
rect 23018 1340 25006 2836
rect 23018 171 23534 1340
rect 23754 171 24270 1340
rect 24490 171 25006 1340
rect 25226 1340 27214 2836
rect 25226 171 25742 1340
rect 25962 171 26478 1340
rect 26698 171 27214 1340
rect 27434 1612 34662 2836
rect 27434 1204 32366 1612
rect 27434 660 29422 1204
rect 27434 171 27950 660
rect 28170 388 29422 660
rect 28170 171 28686 388
rect 28906 171 29422 388
rect 29642 660 32366 1204
rect 29642 171 30158 660
rect 30378 171 30894 660
rect 31114 171 31630 660
rect 31850 171 32366 660
rect 32586 960 34662 1612
rect 35142 960 68460 9920
rect 68940 9540 68982 9920
rect 69202 9812 69718 10573
rect 69938 9812 70454 10573
rect 69202 9540 70454 9812
rect 70674 10084 71190 10573
rect 71410 10356 71926 10573
rect 72146 10356 72662 10573
rect 71410 10084 72662 10356
rect 70674 9540 72662 10084
rect 72882 9540 73398 10573
rect 68940 8996 73398 9540
rect 73618 9540 74134 10573
rect 74354 9540 74870 10573
rect 73618 8996 74870 9540
rect 75090 9540 75606 10573
rect 75826 9540 76342 10573
rect 76562 9812 77078 10573
rect 77298 9812 77814 10573
rect 76562 9540 77814 9812
rect 78034 9812 78550 10573
rect 78770 10084 79286 10573
rect 79506 10084 80022 10573
rect 78770 9812 80022 10084
rect 78034 9540 80022 9812
rect 80242 9812 80758 10573
rect 80978 10492 81494 10573
rect 81714 10492 82230 10573
rect 82450 10492 82966 10573
rect 80978 10084 82966 10492
rect 83186 10084 83702 10573
rect 83922 10084 84438 10573
rect 84658 10084 85174 10573
rect 85394 10084 85910 10573
rect 80978 9812 85910 10084
rect 86130 10492 86646 10573
rect 86866 10492 87382 10573
rect 86130 9812 87382 10492
rect 80242 9540 87382 9812
rect 75090 8996 87382 9540
rect 68940 8588 87382 8996
rect 87602 9132 88118 10573
rect 88338 9132 88854 10573
rect 87602 8588 88854 9132
rect 68940 8044 88854 8588
rect 89074 10220 89590 10573
rect 89810 10220 90326 10573
rect 89074 8588 90326 10220
rect 90546 9948 91062 10573
rect 91282 9948 91798 10573
rect 90546 9132 91798 9948
rect 92018 9676 92534 10573
rect 92754 9676 93270 10573
rect 93490 9676 94006 10573
rect 92018 9132 94006 9676
rect 90546 8588 94006 9132
rect 94226 8588 94742 10573
rect 94962 9676 95478 10573
rect 95698 9676 96214 10573
rect 96434 9676 96950 10573
rect 94962 8588 96950 9676
rect 97170 8588 97686 10573
rect 97906 9676 98422 10573
rect 98642 9676 99158 10573
rect 97906 8588 99158 9676
rect 99378 9676 99894 10573
rect 100114 9676 100630 10573
rect 99378 9132 100630 9676
rect 100850 10220 103114 10573
rect 103334 10220 103850 10573
rect 104070 10220 104586 10573
rect 104806 10220 105322 10573
rect 105542 10220 106058 10573
rect 106278 10220 106794 10573
rect 107014 10220 107530 10573
rect 107750 10220 108266 10573
rect 108486 10220 109002 10573
rect 109222 10220 109738 10573
rect 109958 10220 110474 10573
rect 110694 10220 111210 10573
rect 111430 10220 111946 10573
rect 112166 10220 112682 10573
rect 112902 10220 113418 10573
rect 113638 10220 114154 10573
rect 114374 10220 114890 10573
rect 115110 10220 115626 10573
rect 115846 10220 116362 10573
rect 116582 10220 117098 10573
rect 117318 10220 117834 10573
rect 118054 10220 118570 10573
rect 118790 10220 119306 10573
rect 119526 10220 120042 10573
rect 120262 10220 120778 10573
rect 120998 10220 121514 10573
rect 121734 10220 122250 10573
rect 122470 10220 122986 10573
rect 123206 10220 123722 10573
rect 123942 10220 124458 10573
rect 124678 10356 125194 10573
rect 125414 10356 125930 10573
rect 124678 10220 125930 10356
rect 126150 10220 126666 10573
rect 126886 10220 127402 10573
rect 127622 10220 128138 10573
rect 128358 10220 128874 10573
rect 129094 10220 129610 10573
rect 129830 10220 130346 10573
rect 130566 10220 131082 10573
rect 131302 10220 131818 10573
rect 132038 10220 132554 10573
rect 132774 10220 133290 10573
rect 133510 10220 134026 10573
rect 134246 10220 134762 10573
rect 134982 10220 137246 10573
rect 100850 9920 137246 10220
rect 100850 9132 102259 9920
rect 99378 8588 102259 9132
rect 89074 8044 102259 8588
rect 68940 3788 102259 8044
rect 68940 3108 97686 3788
rect 68940 1612 94006 3108
rect 68940 1476 91062 1612
rect 68940 1340 88118 1476
rect 68940 1068 76342 1340
rect 68940 960 71190 1068
rect 32586 932 71190 960
rect 32586 660 68982 932
rect 32586 171 34850 660
rect 35070 171 35586 660
rect 35806 171 36322 660
rect 36542 171 37058 660
rect 37278 171 37794 660
rect 38014 171 38530 660
rect 38750 388 40002 660
rect 38750 171 39266 388
rect 39486 171 40002 388
rect 40222 171 40738 660
rect 40958 171 41474 660
rect 41694 171 42210 660
rect 42430 171 42946 660
rect 43166 171 43682 660
rect 43902 171 44418 660
rect 44638 171 45154 660
rect 45374 171 45890 660
rect 46110 171 46626 660
rect 46846 171 47362 660
rect 47582 171 48098 660
rect 48318 171 48834 660
rect 49054 171 49570 660
rect 49790 171 50306 660
rect 50526 171 51042 660
rect 51262 171 51778 660
rect 51998 388 53250 660
rect 51998 171 52514 388
rect 52734 171 53250 388
rect 53470 171 53986 660
rect 54206 524 68982 660
rect 54206 450 55458 524
rect 54206 171 54722 450
rect 54942 171 55458 450
rect 55678 171 56194 524
rect 56414 171 56930 524
rect 57150 450 58402 524
rect 57150 171 57666 450
rect 57886 171 58402 450
rect 58622 450 59874 524
rect 58622 171 59138 450
rect 59358 171 59874 450
rect 60094 171 60610 524
rect 60830 171 61346 524
rect 61566 171 62082 524
rect 62302 171 62818 524
rect 63038 388 65762 524
rect 63038 171 63554 388
rect 63774 171 64290 388
rect 64510 171 65026 388
rect 65246 171 65762 388
rect 65982 171 66498 524
rect 66718 171 68982 524
rect 69202 171 69718 932
rect 69938 171 70454 932
rect 70674 171 71190 932
rect 71410 171 71926 1068
rect 72146 932 73398 1068
rect 72146 171 72662 932
rect 72882 171 73398 932
rect 73618 932 75606 1068
rect 73618 171 74134 932
rect 74354 171 74870 932
rect 75090 171 75606 932
rect 75826 171 76342 1068
rect 76562 1068 78550 1340
rect 76562 171 77078 1068
rect 77298 932 78550 1068
rect 77298 171 77814 932
rect 78034 171 78550 932
rect 78770 1068 81494 1340
rect 78770 171 79286 1068
rect 79506 932 80758 1068
rect 79506 171 80022 932
rect 80242 171 80758 932
rect 80978 171 81494 1068
rect 81714 1068 83702 1340
rect 81714 171 82230 1068
rect 82450 932 83702 1068
rect 82450 171 82966 932
rect 83186 171 83702 932
rect 83922 1068 88118 1340
rect 83922 171 84438 1068
rect 84658 388 85910 1068
rect 84658 171 85174 388
rect 85394 171 85910 388
rect 86130 932 88118 1068
rect 86130 171 86646 932
rect 86866 524 88118 932
rect 86866 171 87382 524
rect 87602 171 88118 524
rect 88338 1340 91062 1476
rect 88338 171 88854 1340
rect 89074 450 90326 1340
rect 89074 171 89590 450
rect 89810 171 90326 450
rect 90546 171 91062 1340
rect 91282 1340 94006 1612
rect 91282 171 91798 1340
rect 92018 660 93270 1340
rect 92018 171 92534 660
rect 92754 171 93270 660
rect 93490 171 94006 1340
rect 94226 2836 97686 3108
rect 94226 660 95478 2836
rect 94226 171 94742 660
rect 94962 171 95478 660
rect 95698 1612 96950 2836
rect 95698 171 96214 1612
rect 96434 171 96950 1612
rect 97170 171 97686 2836
rect 97906 3244 102259 3788
rect 97906 1612 100630 3244
rect 97906 171 98422 1612
rect 98642 932 100630 1612
rect 98642 171 99158 932
rect 99378 660 100630 932
rect 99378 171 99894 660
rect 100114 171 100630 660
rect 100850 960 102259 3244
rect 102739 960 136057 9920
rect 136537 9540 137246 9920
rect 137466 10220 137982 10573
rect 138202 10220 138718 10573
rect 137466 10084 138718 10220
rect 138938 10084 139454 10573
rect 137466 9812 139454 10084
rect 139674 10084 140190 10573
rect 140410 10084 140926 10573
rect 141146 10084 141662 10573
rect 141882 10220 142398 10573
rect 142618 10220 143134 10573
rect 141882 10084 143134 10220
rect 143354 10084 143870 10573
rect 144090 10084 144606 10573
rect 139674 9812 144606 10084
rect 144826 10084 145342 10573
rect 145562 10084 146078 10573
rect 146298 10084 146814 10573
rect 147034 10492 147550 10573
rect 147770 10492 148286 10573
rect 147034 10220 148286 10492
rect 148506 10220 149022 10573
rect 147034 10084 149022 10220
rect 149242 10084 149758 10573
rect 144826 9812 149758 10084
rect 149978 10084 150494 10573
rect 150714 10084 151230 10573
rect 151450 10084 151966 10573
rect 152186 10084 152702 10573
rect 152922 10084 153438 10573
rect 153658 10356 154174 10573
rect 154394 10356 154910 10573
rect 153658 10084 154910 10356
rect 149978 9812 154910 10084
rect 155130 9812 155646 10573
rect 137466 9540 155646 9812
rect 136537 8588 155646 9540
rect 155866 9404 156382 10573
rect 156602 9404 157118 10573
rect 155866 8588 157118 9404
rect 136537 8316 157118 8588
rect 157338 8316 157854 10573
rect 136537 8044 157854 8316
rect 158074 8316 158590 10573
rect 158810 8316 159326 10573
rect 158074 8044 159326 8316
rect 159546 8316 160062 10573
rect 160282 8316 160798 10573
rect 159546 8044 160798 8316
rect 161018 8316 161534 10573
rect 161754 8316 162270 10573
rect 161018 8044 162270 8316
rect 136537 7772 162270 8044
rect 162490 8316 163006 10573
rect 163226 8316 163742 10573
rect 162490 8044 163742 8316
rect 163962 8316 164478 10573
rect 164698 8316 165214 10573
rect 163962 8044 165214 8316
rect 165434 8316 165950 10573
rect 166170 8316 166686 10573
rect 166906 9676 167422 10573
rect 167642 9676 168158 10573
rect 166906 9132 168158 9676
rect 168378 9676 168894 10573
rect 169114 10220 171378 10573
rect 171598 10492 172114 10573
rect 172334 10492 172850 10573
rect 171598 10356 172850 10492
rect 173070 10356 173586 10573
rect 171598 10220 173586 10356
rect 173806 10220 174322 10573
rect 174542 10220 175058 10573
rect 175278 10220 175794 10573
rect 176014 10220 176530 10573
rect 176750 10220 177266 10573
rect 177486 10220 178002 10573
rect 178222 10220 178738 10573
rect 178958 10492 179474 10573
rect 179694 10492 180210 10573
rect 178958 10220 180210 10492
rect 180430 10356 180946 10573
rect 181166 10356 181682 10573
rect 180430 10220 181682 10356
rect 181902 10220 182418 10573
rect 182638 10220 183154 10573
rect 183374 10220 183890 10573
rect 184110 10220 184626 10573
rect 184846 10220 185362 10573
rect 185582 10220 186098 10573
rect 186318 10220 186834 10573
rect 187054 10220 187570 10573
rect 187790 10220 188306 10573
rect 188526 10220 189042 10573
rect 189262 10220 189778 10573
rect 189998 10356 190514 10573
rect 190734 10356 191250 10573
rect 189998 10220 191250 10356
rect 191470 10220 191986 10573
rect 192206 10356 192722 10573
rect 192942 10356 193458 10573
rect 192206 10220 193458 10356
rect 193678 10220 194194 10573
rect 194414 10220 194930 10573
rect 195150 10220 195666 10573
rect 195886 10220 196402 10573
rect 196622 10220 197138 10573
rect 197358 10220 197874 10573
rect 198094 10220 198610 10573
rect 198830 10220 199346 10573
rect 199566 10220 200082 10573
rect 200302 10220 200818 10573
rect 201038 10220 201554 10573
rect 201774 10356 202290 10573
rect 202510 10356 203026 10573
rect 201774 10220 203026 10356
rect 203246 10220 205510 10573
rect 205730 10220 206246 10573
rect 169114 10084 206246 10220
rect 206466 10084 206982 10573
rect 207202 10492 207718 10573
rect 207938 10492 208454 10573
rect 207202 10084 208454 10492
rect 208674 10084 209190 10573
rect 209410 10356 209926 10573
rect 210146 10356 210662 10573
rect 209410 10084 210662 10356
rect 210882 10084 211398 10573
rect 169114 9920 211398 10084
rect 169114 9676 169856 9920
rect 168378 9132 169856 9676
rect 166906 8316 169856 9132
rect 165434 8044 169856 8316
rect 162490 7772 169856 8044
rect 136537 3380 169856 7772
rect 136537 3244 154174 3380
rect 136537 1884 144606 3244
rect 136537 1476 140190 1884
rect 136537 960 137246 1476
rect 100850 660 137246 960
rect 100850 524 124458 660
rect 100850 450 117834 524
rect 100850 171 103114 450
rect 103334 171 103850 450
rect 104070 171 104586 450
rect 104806 171 105322 450
rect 105542 171 106058 450
rect 106278 171 106794 450
rect 107014 171 107530 450
rect 107750 171 108266 450
rect 108486 171 109002 450
rect 109222 171 109738 450
rect 109958 171 110474 450
rect 110694 171 111210 450
rect 111430 171 111946 450
rect 112166 171 112682 450
rect 112902 171 113418 450
rect 113638 171 114154 450
rect 114374 171 114890 450
rect 115110 171 115626 450
rect 115846 171 116362 450
rect 116582 171 117098 450
rect 117318 171 117834 450
rect 118054 171 118570 524
rect 118790 171 119306 524
rect 119526 171 120042 524
rect 120262 171 120778 524
rect 120998 171 121514 524
rect 121734 171 122250 524
rect 122470 171 122986 524
rect 123206 450 124458 524
rect 123206 171 123722 450
rect 123942 171 124458 450
rect 124678 171 125194 660
rect 125414 171 125930 660
rect 126150 524 128874 660
rect 126150 450 127402 524
rect 126150 171 126666 450
rect 126886 171 127402 450
rect 127622 450 128874 524
rect 127622 171 128138 450
rect 128358 171 128874 450
rect 129094 388 130346 660
rect 129094 171 129610 388
rect 129830 171 130346 388
rect 130566 171 131082 660
rect 131302 450 134026 660
rect 131302 388 133290 450
rect 131302 171 131818 388
rect 132038 171 132554 388
rect 132774 171 133290 388
rect 133510 171 134026 450
rect 134246 450 137246 660
rect 134246 171 134762 450
rect 134982 171 137246 450
rect 137466 1068 140190 1476
rect 137466 796 139454 1068
rect 137466 660 138718 796
rect 137466 171 137982 660
rect 138202 171 138718 660
rect 138938 171 139454 796
rect 139674 171 140190 1068
rect 140410 1476 144606 1884
rect 140410 171 140926 1476
rect 141146 796 144606 1476
rect 141146 171 141662 796
rect 141882 171 142398 796
rect 142618 660 144606 796
rect 142618 171 143134 660
rect 143354 524 144606 660
rect 143354 171 143870 524
rect 144090 171 144606 524
rect 144826 2972 154174 3244
rect 144826 2836 149022 2972
rect 144826 171 145342 2836
rect 145562 796 149022 2836
rect 145562 171 146078 796
rect 146298 660 148286 796
rect 146298 388 147550 660
rect 146298 171 146814 388
rect 147034 171 147550 388
rect 147770 171 148286 660
rect 148506 171 149022 796
rect 149242 1476 153438 2972
rect 149242 796 150494 1476
rect 149242 171 149758 796
rect 149978 171 150494 796
rect 150714 660 151966 1476
rect 150714 171 151230 660
rect 151450 171 151966 660
rect 152186 1340 153438 1476
rect 152186 171 152702 1340
rect 152922 171 153438 1340
rect 153658 171 154174 2972
rect 154394 2972 169856 3380
rect 154394 171 154910 2972
rect 155130 2836 169856 2972
rect 155130 1476 156382 2836
rect 155130 171 155646 1476
rect 155866 171 156382 1476
rect 156602 1476 169856 2836
rect 156602 171 157118 1476
rect 157338 1340 168158 1476
rect 157338 171 157854 1340
rect 158074 1204 168158 1340
rect 158074 171 158590 1204
rect 158810 660 160062 1204
rect 158810 171 159326 660
rect 159546 171 160062 660
rect 160282 388 161534 1204
rect 160282 171 160798 388
rect 161018 171 161534 388
rect 161754 660 163742 1204
rect 161754 171 162270 660
rect 162490 171 163006 660
rect 163226 171 163742 660
rect 163962 660 165214 1204
rect 163962 171 164478 660
rect 164698 171 165214 660
rect 165434 171 165950 1204
rect 166170 171 166686 1204
rect 166906 388 168158 1204
rect 166906 171 167422 388
rect 167642 171 168158 388
rect 168378 960 169856 1476
rect 170336 960 203654 9920
rect 204134 9812 211398 9920
rect 211618 10084 212134 10573
rect 212354 10492 212870 10573
rect 213090 10492 213606 10573
rect 212354 10084 213606 10492
rect 213826 10084 214342 10573
rect 214562 10084 215078 10573
rect 211618 9812 215078 10084
rect 204134 9540 215078 9812
rect 215298 10084 215814 10573
rect 216034 10084 216550 10573
rect 215298 9812 216550 10084
rect 216770 10084 217286 10573
rect 217506 10492 218022 10573
rect 218242 10492 218758 10573
rect 217506 10084 218758 10492
rect 218978 10084 219494 10573
rect 219714 10220 220230 10573
rect 220450 10356 220966 10573
rect 221186 10356 221702 10573
rect 220450 10220 221702 10356
rect 219714 10084 221702 10220
rect 216770 9812 221702 10084
rect 221922 10084 222438 10573
rect 222658 10084 223174 10573
rect 223394 10084 223910 10573
rect 221922 9812 223910 10084
rect 215298 9540 223910 9812
rect 204134 9404 223910 9540
rect 224130 9404 224646 10573
rect 204134 8588 224646 9404
rect 224866 8588 225382 10573
rect 225602 8588 226118 10573
rect 226338 8588 226854 10573
rect 227074 9404 227590 10573
rect 227810 9404 228326 10573
rect 228546 9404 229062 10573
rect 227074 8588 229062 9404
rect 229282 9404 229798 10573
rect 230018 9404 230534 10573
rect 229282 8588 230534 9404
rect 230754 8588 231270 10573
rect 231490 9404 232006 10573
rect 232226 9404 232742 10573
rect 231490 8588 232742 9404
rect 232962 9404 233478 10573
rect 233698 9404 234214 10573
rect 232962 8588 234214 9404
rect 234434 8588 234950 10573
rect 204134 8316 234950 8588
rect 235170 9404 235686 10573
rect 235906 9404 236422 10573
rect 235170 9132 236422 9404
rect 236642 9132 237158 10573
rect 235170 8588 237158 9132
rect 237378 10220 239642 10573
rect 239862 10220 240378 10573
rect 240598 10220 241114 10573
rect 241334 10220 241850 10573
rect 242070 10220 242586 10573
rect 242806 10220 243322 10573
rect 243542 10220 244058 10573
rect 244278 10220 244794 10573
rect 245014 10356 245530 10573
rect 245750 10356 246266 10573
rect 245014 10220 246266 10356
rect 246486 10220 247002 10573
rect 247222 10220 247738 10573
rect 247958 10220 248474 10573
rect 248694 10220 249210 10573
rect 249430 10220 249946 10573
rect 250166 10220 250682 10573
rect 250902 10220 251418 10573
rect 251638 10220 252154 10573
rect 252374 10356 252890 10573
rect 253110 10356 253626 10573
rect 252374 10220 253626 10356
rect 253846 10220 254362 10573
rect 254582 10220 255098 10573
rect 255318 10220 255834 10573
rect 256054 10220 256570 10573
rect 256790 10220 257306 10573
rect 257526 10220 258042 10573
rect 258262 10220 258778 10573
rect 258998 10220 259514 10573
rect 259734 10220 260250 10573
rect 260470 10356 260986 10573
rect 261206 10356 261722 10573
rect 260470 10220 261722 10356
rect 261942 10220 262458 10573
rect 262678 10220 263194 10573
rect 263414 10220 263930 10573
rect 264150 10220 264666 10573
rect 264886 10356 265402 10573
rect 265622 10356 266138 10573
rect 237378 10158 264666 10220
rect 264886 10220 266138 10356
rect 266358 10220 266874 10573
rect 264886 10158 266874 10220
rect 267094 10158 267610 10573
rect 267830 10158 268346 10573
rect 268566 10158 269082 10573
rect 269302 10158 269818 10573
rect 270038 10158 270554 10573
rect 270774 10158 271290 10573
rect 237378 9920 271370 10158
rect 237378 8588 237453 9920
rect 235170 8316 237453 8588
rect 204134 4060 237453 8316
rect 204134 3108 215078 4060
rect 204134 2836 211398 3108
rect 204134 1476 210662 2836
rect 204134 960 209926 1476
rect 168378 932 209926 960
rect 168378 660 205510 932
rect 168378 171 168894 660
rect 169114 171 171378 660
rect 171598 171 172114 660
rect 172334 171 172850 660
rect 173070 171 173586 660
rect 173806 171 174322 660
rect 174542 171 175058 660
rect 175278 524 176530 660
rect 175278 171 175794 524
rect 176014 171 176530 524
rect 176750 171 177266 660
rect 177486 171 178002 660
rect 178222 171 178738 660
rect 178958 171 179474 660
rect 179694 171 180210 660
rect 180430 524 205510 660
rect 180430 388 181682 524
rect 180430 171 180946 388
rect 181166 171 181682 388
rect 181902 171 182418 524
rect 182638 171 183154 524
rect 183374 171 183890 524
rect 184110 171 184626 524
rect 184846 171 185362 524
rect 185582 450 186834 524
rect 185582 171 186098 450
rect 186318 171 186834 450
rect 187054 171 187570 524
rect 187790 171 188306 524
rect 188526 171 189042 524
rect 189262 450 190514 524
rect 189262 171 189778 450
rect 189998 171 190514 450
rect 190734 450 192722 524
rect 190734 171 191250 450
rect 191470 388 192722 450
rect 191470 171 191986 388
rect 192206 171 192722 388
rect 192942 171 193458 524
rect 193678 450 194930 524
rect 193678 171 194194 450
rect 194414 171 194930 450
rect 195150 450 196402 524
rect 195150 171 195666 450
rect 195886 171 196402 450
rect 196622 450 198610 524
rect 196622 171 197138 450
rect 197358 171 197874 450
rect 198094 171 198610 450
rect 198830 450 200082 524
rect 198830 171 199346 450
rect 199566 171 200082 450
rect 200302 450 202290 524
rect 200302 171 200818 450
rect 201038 171 201554 450
rect 201774 171 202290 450
rect 202510 171 203026 524
rect 203246 171 205510 524
rect 205730 171 206246 932
rect 206466 171 206982 932
rect 207202 388 208454 932
rect 207202 171 207718 388
rect 207938 171 208454 388
rect 208674 524 209926 932
rect 208674 171 209190 524
rect 209410 171 209926 524
rect 210146 171 210662 1476
rect 210882 171 211398 2836
rect 211618 1884 215078 3108
rect 211618 171 212134 1884
rect 212354 524 215078 1884
rect 212354 388 213606 524
rect 212354 171 212870 388
rect 213090 171 213606 388
rect 213826 388 215078 524
rect 213826 171 214342 388
rect 214562 171 215078 388
rect 215298 3788 237453 4060
rect 215298 3244 218758 3788
rect 215298 2972 217286 3244
rect 215298 796 216550 2972
rect 215298 171 215814 796
rect 216034 171 216550 796
rect 216770 171 217286 2972
rect 217506 1476 218758 3244
rect 217506 171 218022 1476
rect 218242 171 218758 1476
rect 218978 3244 223174 3788
rect 218978 1476 220966 3244
rect 218978 171 219494 1476
rect 219714 388 220966 1476
rect 219714 171 220230 388
rect 220450 171 220966 388
rect 221186 1476 223174 3244
rect 221186 660 222438 1476
rect 221186 171 221702 660
rect 221922 171 222438 660
rect 222658 171 223174 1476
rect 223394 1612 237453 3788
rect 223394 1476 237158 1612
rect 223394 1204 226118 1476
rect 223394 171 223910 1204
rect 224130 796 225382 1204
rect 224130 171 224646 796
rect 224866 171 225382 796
rect 225602 171 226118 1204
rect 226338 1204 237158 1476
rect 226338 660 227590 1204
rect 226338 171 226854 660
rect 227074 171 227590 660
rect 227810 660 229798 1204
rect 227810 171 228326 660
rect 228546 171 229062 660
rect 229282 171 229798 660
rect 230018 171 230534 1204
rect 230754 660 232006 1204
rect 230754 171 231270 660
rect 231490 171 232006 660
rect 232226 171 232742 1204
rect 232962 660 234950 1204
rect 232962 171 233478 660
rect 233698 171 234214 660
rect 234434 171 234950 660
rect 235170 660 236422 1204
rect 235170 171 235686 660
rect 235906 171 236422 660
rect 236642 171 237158 1204
rect 237378 960 237453 1612
rect 237933 960 271251 9920
rect 237378 722 271370 960
rect 237378 660 246266 722
rect 237378 171 239642 660
rect 239862 171 240378 660
rect 240598 171 241114 660
rect 241334 171 241850 660
rect 242070 450 243322 660
rect 242070 171 242586 450
rect 242806 171 243322 450
rect 243542 171 244058 660
rect 244278 171 244794 660
rect 245014 450 246266 660
rect 246486 660 250682 722
rect 245014 171 245530 450
rect 245750 171 246266 450
rect 246486 171 247002 660
rect 247222 171 247738 660
rect 247958 450 249946 660
rect 247958 171 248474 450
rect 248694 171 249210 450
rect 249430 171 249946 450
rect 250166 171 250682 660
rect 250902 660 255834 722
rect 250902 524 254362 660
rect 250902 450 252890 524
rect 250902 171 251418 450
rect 251638 171 252154 450
rect 252374 171 252890 450
rect 253110 388 254362 524
rect 253110 171 253626 388
rect 253846 171 254362 388
rect 254582 171 255098 660
rect 255318 171 255834 660
rect 256054 660 258778 722
rect 256054 450 258042 660
rect 256054 171 256570 450
rect 256790 171 257306 450
rect 257526 171 258042 450
rect 258262 171 258778 660
rect 258998 171 259514 722
rect 259734 171 260250 722
rect 260470 660 261722 722
rect 260470 171 260986 660
rect 261206 171 261722 660
rect 261942 660 271290 722
rect 261942 171 262458 660
rect 262678 171 263194 660
rect 263414 171 263930 660
rect 264150 171 264666 660
rect 264886 171 265402 660
rect 265622 171 266138 660
rect 266358 171 266874 660
rect 267094 171 267610 660
rect 267830 171 268346 660
rect 268566 171 269082 660
rect 269302 388 270554 660
rect 269302 171 269818 388
rect 270038 171 270554 388
rect 270774 171 271290 660
<< labels >>
rlabel metal3 s 270554 9558 272504 9618 6 addr[0]
port 1 nsew signal input
rlabel metal3 s 272210 9422 272504 9482 6 addr[1]
port 2 nsew signal input
rlabel metal3 s 268070 9286 272504 9346 6 addr[2]
port 3 nsew signal input
rlabel metal3 s 268806 9150 272504 9210 6 addr[3]
port 4 nsew signal input
rlabel metal3 s 268714 9014 272504 9074 6 addr[4]
port 5 nsew signal input
rlabel metal3 s 272026 8878 272504 8938 6 k_one
port 6 nsew signal output
rlabel metal3 s 271830 8742 272504 8802 6 k_zero
port 7 nsew signal output
rlabel metal3 s 272304 8606 272504 8666 6 spine_iw[0]
port 8 nsew signal input
rlabel metal3 s 262366 7246 272504 7306 6 spine_iw[10]
port 9 nsew signal input
rlabel metal3 s 263286 7110 272504 7170 6 spine_iw[11]
port 10 nsew signal input
rlabel metal3 s 267978 6974 272504 7034 6 spine_iw[12]
port 11 nsew signal input
rlabel metal3 s 267978 6838 272504 6898 6 spine_iw[13]
port 12 nsew signal input
rlabel metal3 s 271014 6702 272504 6762 6 spine_iw[14]
port 13 nsew signal input
rlabel metal3 s 272118 6566 272504 6626 6 spine_iw[15]
port 14 nsew signal input
rlabel metal3 s 271934 6430 272504 6490 6 spine_iw[16]
port 15 nsew signal input
rlabel metal3 s 271382 6294 272504 6354 6 spine_iw[17]
port 16 nsew signal input
rlabel metal3 s 270542 6158 272504 6218 6 spine_iw[18]
port 17 nsew signal input
rlabel metal3 s 271750 6022 272504 6082 6 spine_iw[19]
port 18 nsew signal input
rlabel metal3 s 268346 8470 272504 8530 6 spine_iw[1]
port 19 nsew signal input
rlabel metal3 s 271198 5886 272504 5946 6 spine_iw[20]
port 20 nsew signal input
rlabel metal3 s 270910 5750 272504 5810 6 spine_iw[21]
port 21 nsew signal input
rlabel metal3 s 270726 5614 272504 5674 6 spine_iw[22]
port 22 nsew signal input
rlabel metal3 s 271842 5478 272504 5538 6 spine_iw[23]
port 23 nsew signal input
rlabel metal3 s 271842 5342 272504 5402 6 spine_iw[24]
port 24 nsew signal input
rlabel metal3 s 269082 5206 272504 5266 6 spine_iw[25]
port 25 nsew signal input
rlabel metal3 s 268530 5070 272504 5130 6 spine_iw[26]
port 26 nsew signal input
rlabel metal3 s 272026 4934 272504 4994 6 spine_iw[27]
port 27 nsew signal input
rlabel metal3 s 268990 4798 272504 4858 6 spine_iw[28]
port 28 nsew signal input
rlabel metal3 s 268346 4662 272504 4722 6 spine_iw[29]
port 29 nsew signal input
rlabel metal3 s 268070 8334 272504 8394 6 spine_iw[2]
port 30 nsew signal input
rlabel metal3 s 272304 4526 272504 4586 6 spine_iw[30]
port 31 nsew signal input
rlabel metal3 s 272014 8198 272504 8258 6 spine_iw[3]
port 32 nsew signal input
rlabel metal3 s 272210 8062 272504 8122 6 spine_iw[4]
port 33 nsew signal input
rlabel metal3 s 272210 7926 272504 7986 6 spine_iw[5]
port 34 nsew signal input
rlabel metal3 s 264942 7790 272504 7850 6 spine_iw[6]
port 35 nsew signal input
rlabel metal3 s 271842 7654 272504 7714 6 spine_iw[7]
port 36 nsew signal input
rlabel metal3 s 271830 7518 272504 7578 6 spine_iw[8]
port 37 nsew signal input
rlabel metal3 s 272026 7382 272504 7442 6 spine_iw[9]
port 38 nsew signal input
rlabel metal3 s 271830 4390 272504 4450 6 spine_ow[0]
port 39 nsew signal output
rlabel metal3 s 267978 3030 272504 3090 6 spine_ow[10]
port 40 nsew signal output
rlabel metal3 s 258766 2894 272504 2954 6 spine_ow[11]
port 41 nsew signal output
rlabel metal3 s 271290 2758 272504 2818 6 spine_ow[12]
port 42 nsew signal output
rlabel metal3 s 267978 2622 272504 2682 6 spine_ow[13]
port 43 nsew signal output
rlabel metal3 s 268438 2486 272504 2546 6 spine_ow[14]
port 44 nsew signal output
rlabel metal3 s 248474 2350 272504 2410 6 spine_ow[15]
port 45 nsew signal output
rlabel metal3 s 271830 2214 272504 2274 6 spine_ow[16]
port 46 nsew signal output
rlabel metal3 s 272026 2078 272504 2138 6 spine_ow[17]
port 47 nsew signal output
rlabel metal3 s 272118 1942 272504 2002 6 spine_ow[18]
port 48 nsew signal output
rlabel metal3 s 268898 1806 272504 1866 6 spine_ow[19]
port 49 nsew signal output
rlabel metal3 s 271842 4254 272504 4314 6 spine_ow[1]
port 50 nsew signal output
rlabel metal3 s 269622 1670 272504 1730 6 spine_ow[20]
port 51 nsew signal output
rlabel metal3 s 272210 1534 272504 1594 6 spine_ow[21]
port 52 nsew signal output
rlabel metal3 s 258778 1398 272504 1458 6 spine_ow[22]
port 53 nsew signal output
rlabel metal3 s 272026 1262 272504 1322 6 spine_ow[23]
port 54 nsew signal output
rlabel metal3 s 271830 1126 272504 1186 6 spine_ow[24]
port 55 nsew signal output
rlabel metal3 s 272198 990 272504 1050 6 spine_ow[25]
port 56 nsew signal output
rlabel metal3 s 271830 4118 272504 4178 6 spine_ow[2]
port 57 nsew signal output
rlabel metal3 s 272014 3982 272504 4042 6 spine_ow[3]
port 58 nsew signal output
rlabel metal3 s 272210 3846 272504 3906 6 spine_ow[4]
port 59 nsew signal output
rlabel metal3 s 268070 3710 272504 3770 6 spine_ow[5]
port 60 nsew signal output
rlabel metal3 s 272210 3574 272504 3634 6 spine_ow[6]
port 61 nsew signal output
rlabel metal3 s 272014 3438 272504 3498 6 spine_ow[7]
port 62 nsew signal output
rlabel metal3 s 271830 3302 272504 3362 6 spine_ow[8]
port 63 nsew signal output
rlabel metal3 s 271842 3166 272504 3226 6 spine_ow[9]
port 64 nsew signal output
rlabel metal4 s 32446 0 32506 1532 6 um_ena[0]
port 65 nsew signal output
rlabel metal4 s 203106 0 203166 444 6 um_ena[10]
port 66 nsew signal output
rlabel metal4 s 203106 10300 203166 10880 6 um_ena[11]
port 67 nsew signal output
rlabel metal4 s 237238 0 237298 1532 6 um_ena[12]
port 68 nsew signal output
rlabel metal4 s 237238 8668 237298 10880 6 um_ena[13]
port 69 nsew signal output
rlabel metal4 s 271370 0 271430 642 6 um_ena[14]
port 70 nsew signal output
rlabel metal4 s 271370 10238 271430 10880 6 um_ena[15]
port 71 nsew signal output
rlabel metal4 s 32446 9212 32506 10880 6 um_ena[1]
port 72 nsew signal output
rlabel metal4 s 66578 0 66638 444 6 um_ena[2]
port 73 nsew signal output
rlabel metal4 s 66578 10300 66638 10880 6 um_ena[3]
port 74 nsew signal output
rlabel metal4 s 100710 0 100770 3164 6 um_ena[4]
port 75 nsew signal output
rlabel metal4 s 100710 9212 100770 10880 6 um_ena[5]
port 76 nsew signal output
rlabel metal4 s 134842 0 134902 370 6 um_ena[6]
port 77 nsew signal output
rlabel metal4 s 134842 10300 134902 10880 6 um_ena[7]
port 78 nsew signal output
rlabel metal4 s 168974 0 169034 580 6 um_ena[8]
port 79 nsew signal output
rlabel metal4 s 168974 9756 169034 10880 6 um_ena[9]
port 80 nsew signal output
rlabel metal4 s 31710 0 31770 580 6 um_iw[0]
port 81 nsew signal output
rlabel metal4 s 92614 9756 92674 10880 6 um_iw[100]
port 82 nsew signal output
rlabel metal4 s 91878 9212 91938 10880 6 um_iw[101]
port 83 nsew signal output
rlabel metal4 s 91142 10028 91202 10880 6 um_iw[102]
port 84 nsew signal output
rlabel metal4 s 90406 8668 90466 10880 6 um_iw[103]
port 85 nsew signal output
rlabel metal4 s 89670 10300 89730 10880 6 um_iw[104]
port 86 nsew signal output
rlabel metal4 s 88934 8124 88994 10880 6 um_iw[105]
port 87 nsew signal output
rlabel metal4 s 88198 9212 88258 10880 6 um_iw[106]
port 88 nsew signal output
rlabel metal4 s 87462 8668 87522 10880 6 um_iw[107]
port 89 nsew signal output
rlabel metal4 s 134106 0 134166 580 6 um_iw[108]
port 90 nsew signal output
rlabel metal4 s 133370 0 133430 370 6 um_iw[109]
port 91 nsew signal output
rlabel metal4 s 24350 0 24410 1260 6 um_iw[10]
port 92 nsew signal output
rlabel metal4 s 132634 0 132694 308 6 um_iw[110]
port 93 nsew signal output
rlabel metal4 s 131898 0 131958 308 6 um_iw[111]
port 94 nsew signal output
rlabel metal4 s 131162 0 131222 580 6 um_iw[112]
port 95 nsew signal output
rlabel metal4 s 130426 0 130486 580 6 um_iw[113]
port 96 nsew signal output
rlabel metal4 s 129690 0 129750 308 6 um_iw[114]
port 97 nsew signal output
rlabel metal4 s 128954 0 129014 580 6 um_iw[115]
port 98 nsew signal output
rlabel metal4 s 128218 0 128278 370 6 um_iw[116]
port 99 nsew signal output
rlabel metal4 s 127482 0 127542 444 6 um_iw[117]
port 100 nsew signal output
rlabel metal4 s 126746 0 126806 370 6 um_iw[118]
port 101 nsew signal output
rlabel metal4 s 126010 0 126070 580 6 um_iw[119]
port 102 nsew signal output
rlabel metal4 s 23614 0 23674 1260 6 um_iw[11]
port 103 nsew signal output
rlabel metal4 s 125274 0 125334 580 6 um_iw[120]
port 104 nsew signal output
rlabel metal4 s 124538 0 124598 580 6 um_iw[121]
port 105 nsew signal output
rlabel metal4 s 123802 0 123862 370 6 um_iw[122]
port 106 nsew signal output
rlabel metal4 s 123066 0 123126 444 6 um_iw[123]
port 107 nsew signal output
rlabel metal4 s 122330 0 122390 444 6 um_iw[124]
port 108 nsew signal output
rlabel metal4 s 121594 0 121654 444 6 um_iw[125]
port 109 nsew signal output
rlabel metal4 s 134106 10300 134166 10880 6 um_iw[126]
port 110 nsew signal output
rlabel metal4 s 133370 10300 133430 10880 6 um_iw[127]
port 111 nsew signal output
rlabel metal4 s 132634 10300 132694 10880 6 um_iw[128]
port 112 nsew signal output
rlabel metal4 s 131898 10300 131958 10880 6 um_iw[129]
port 113 nsew signal output
rlabel metal4 s 22878 0 22938 2756 6 um_iw[12]
port 114 nsew signal output
rlabel metal4 s 131162 10300 131222 10880 6 um_iw[130]
port 115 nsew signal output
rlabel metal4 s 130426 10300 130486 10880 6 um_iw[131]
port 116 nsew signal output
rlabel metal4 s 129690 10300 129750 10880 6 um_iw[132]
port 117 nsew signal output
rlabel metal4 s 128954 10300 129014 10880 6 um_iw[133]
port 118 nsew signal output
rlabel metal4 s 128218 10300 128278 10880 6 um_iw[134]
port 119 nsew signal output
rlabel metal4 s 127482 10300 127542 10880 6 um_iw[135]
port 120 nsew signal output
rlabel metal4 s 126746 10300 126806 10880 6 um_iw[136]
port 121 nsew signal output
rlabel metal4 s 126010 10300 126070 10880 6 um_iw[137]
port 122 nsew signal output
rlabel metal4 s 125274 10436 125334 10880 6 um_iw[138]
port 123 nsew signal output
rlabel metal4 s 124538 10300 124598 10880 6 um_iw[139]
port 124 nsew signal output
rlabel metal4 s 22142 0 22202 1668 6 um_iw[13]
port 125 nsew signal output
rlabel metal4 s 123802 10300 123862 10880 6 um_iw[140]
port 126 nsew signal output
rlabel metal4 s 123066 10300 123126 10880 6 um_iw[141]
port 127 nsew signal output
rlabel metal4 s 122330 10300 122390 10880 6 um_iw[142]
port 128 nsew signal output
rlabel metal4 s 121594 10300 121654 10880 6 um_iw[143]
port 129 nsew signal output
rlabel metal4 s 168238 0 168298 1396 6 um_iw[144]
port 130 nsew signal output
rlabel metal4 s 167502 0 167562 308 6 um_iw[145]
port 131 nsew signal output
rlabel metal4 s 166766 0 166826 1124 6 um_iw[146]
port 132 nsew signal output
rlabel metal4 s 166030 0 166090 1124 6 um_iw[147]
port 133 nsew signal output
rlabel metal4 s 165294 0 165354 1124 6 um_iw[148]
port 134 nsew signal output
rlabel metal4 s 164558 0 164618 580 6 um_iw[149]
port 135 nsew signal output
rlabel metal4 s 21406 0 21466 580 6 um_iw[14]
port 136 nsew signal output
rlabel metal4 s 163822 0 163882 1124 6 um_iw[150]
port 137 nsew signal output
rlabel metal4 s 163086 0 163146 580 6 um_iw[151]
port 138 nsew signal output
rlabel metal4 s 162350 0 162410 580 6 um_iw[152]
port 139 nsew signal output
rlabel metal4 s 161614 0 161674 1124 6 um_iw[153]
port 140 nsew signal output
rlabel metal4 s 160878 0 160938 308 6 um_iw[154]
port 141 nsew signal output
rlabel metal4 s 160142 0 160202 1124 6 um_iw[155]
port 142 nsew signal output
rlabel metal4 s 159406 0 159466 580 6 um_iw[156]
port 143 nsew signal output
rlabel metal4 s 158670 0 158730 1124 6 um_iw[157]
port 144 nsew signal output
rlabel metal4 s 157934 0 157994 1260 6 um_iw[158]
port 145 nsew signal output
rlabel metal4 s 157198 0 157258 1396 6 um_iw[159]
port 146 nsew signal output
rlabel metal4 s 20670 0 20730 1396 6 um_iw[15]
port 147 nsew signal output
rlabel metal4 s 156462 0 156522 2756 6 um_iw[160]
port 148 nsew signal output
rlabel metal4 s 155726 0 155786 1396 6 um_iw[161]
port 149 nsew signal output
rlabel metal4 s 168238 9212 168298 10880 6 um_iw[162]
port 150 nsew signal output
rlabel metal4 s 167502 9756 167562 10880 6 um_iw[163]
port 151 nsew signal output
rlabel metal4 s 166766 8396 166826 10880 6 um_iw[164]
port 152 nsew signal output
rlabel metal4 s 166030 8396 166090 10880 6 um_iw[165]
port 153 nsew signal output
rlabel metal4 s 165294 8124 165354 10880 6 um_iw[166]
port 154 nsew signal output
rlabel metal4 s 164558 8396 164618 10880 6 um_iw[167]
port 155 nsew signal output
rlabel metal4 s 163822 8124 163882 10880 6 um_iw[168]
port 156 nsew signal output
rlabel metal4 s 163086 8396 163146 10880 6 um_iw[169]
port 157 nsew signal output
rlabel metal4 s 19934 0 19994 1532 6 um_iw[16]
port 158 nsew signal output
rlabel metal4 s 162350 7852 162410 10880 6 um_iw[170]
port 159 nsew signal output
rlabel metal4 s 161614 8396 161674 10880 6 um_iw[171]
port 160 nsew signal output
rlabel metal4 s 160878 8124 160938 10880 6 um_iw[172]
port 161 nsew signal output
rlabel metal4 s 160142 8396 160202 10880 6 um_iw[173]
port 162 nsew signal output
rlabel metal4 s 159406 8124 159466 10880 6 um_iw[174]
port 163 nsew signal output
rlabel metal4 s 158670 8396 158730 10880 6 um_iw[175]
port 164 nsew signal output
rlabel metal4 s 157934 8124 157994 10880 6 um_iw[176]
port 165 nsew signal output
rlabel metal4 s 157198 8396 157258 10880 6 um_iw[177]
port 166 nsew signal output
rlabel metal4 s 156462 9484 156522 10880 6 um_iw[178]
port 167 nsew signal output
rlabel metal4 s 155726 8668 155786 10880 6 um_iw[179]
port 168 nsew signal output
rlabel metal4 s 19198 0 19258 2756 6 um_iw[17]
port 169 nsew signal output
rlabel metal4 s 202370 0 202430 444 6 um_iw[180]
port 170 nsew signal output
rlabel metal4 s 201634 0 201694 370 6 um_iw[181]
port 171 nsew signal output
rlabel metal4 s 200898 0 200958 370 6 um_iw[182]
port 172 nsew signal output
rlabel metal4 s 200162 0 200222 444 6 um_iw[183]
port 173 nsew signal output
rlabel metal4 s 199426 0 199486 370 6 um_iw[184]
port 174 nsew signal output
rlabel metal4 s 198690 0 198750 444 6 um_iw[185]
port 175 nsew signal output
rlabel metal4 s 197954 0 198014 370 6 um_iw[186]
port 176 nsew signal output
rlabel metal4 s 197218 0 197278 370 6 um_iw[187]
port 177 nsew signal output
rlabel metal4 s 196482 0 196542 444 6 um_iw[188]
port 178 nsew signal output
rlabel metal4 s 195746 0 195806 370 6 um_iw[189]
port 179 nsew signal output
rlabel metal4 s 31710 10300 31770 10880 6 um_iw[18]
port 180 nsew signal output
rlabel metal4 s 195010 0 195070 444 6 um_iw[190]
port 181 nsew signal output
rlabel metal4 s 194274 0 194334 370 6 um_iw[191]
port 182 nsew signal output
rlabel metal4 s 193538 0 193598 444 6 um_iw[192]
port 183 nsew signal output
rlabel metal4 s 192802 0 192862 444 6 um_iw[193]
port 184 nsew signal output
rlabel metal4 s 192066 0 192126 308 6 um_iw[194]
port 185 nsew signal output
rlabel metal4 s 191330 0 191390 370 6 um_iw[195]
port 186 nsew signal output
rlabel metal4 s 190594 0 190654 444 6 um_iw[196]
port 187 nsew signal output
rlabel metal4 s 189858 0 189918 370 6 um_iw[197]
port 188 nsew signal output
rlabel metal4 s 202370 10436 202430 10880 6 um_iw[198]
port 189 nsew signal output
rlabel metal4 s 201634 10300 201694 10880 6 um_iw[199]
port 190 nsew signal output
rlabel metal4 s 30974 8668 31034 10880 6 um_iw[19]
port 191 nsew signal output
rlabel metal4 s 30974 0 31034 580 6 um_iw[1]
port 192 nsew signal output
rlabel metal4 s 200898 10300 200958 10880 6 um_iw[200]
port 193 nsew signal output
rlabel metal4 s 200162 10300 200222 10880 6 um_iw[201]
port 194 nsew signal output
rlabel metal4 s 199426 10300 199486 10880 6 um_iw[202]
port 195 nsew signal output
rlabel metal4 s 198690 10300 198750 10880 6 um_iw[203]
port 196 nsew signal output
rlabel metal4 s 197954 10300 198014 10880 6 um_iw[204]
port 197 nsew signal output
rlabel metal4 s 197218 10300 197278 10880 6 um_iw[205]
port 198 nsew signal output
rlabel metal4 s 196482 10300 196542 10880 6 um_iw[206]
port 199 nsew signal output
rlabel metal4 s 195746 10300 195806 10880 6 um_iw[207]
port 200 nsew signal output
rlabel metal4 s 195010 10300 195070 10880 6 um_iw[208]
port 201 nsew signal output
rlabel metal4 s 194274 10300 194334 10880 6 um_iw[209]
port 202 nsew signal output
rlabel metal4 s 30238 9756 30298 10880 6 um_iw[20]
port 203 nsew signal output
rlabel metal4 s 193538 10300 193598 10880 6 um_iw[210]
port 204 nsew signal output
rlabel metal4 s 192802 10436 192862 10880 6 um_iw[211]
port 205 nsew signal output
rlabel metal4 s 192066 10300 192126 10880 6 um_iw[212]
port 206 nsew signal output
rlabel metal4 s 191330 10300 191390 10880 6 um_iw[213]
port 207 nsew signal output
rlabel metal4 s 190594 10436 190654 10880 6 um_iw[214]
port 208 nsew signal output
rlabel metal4 s 189858 10300 189918 10880 6 um_iw[215]
port 209 nsew signal output
rlabel metal4 s 236502 0 236562 1124 6 um_iw[216]
port 210 nsew signal output
rlabel metal4 s 235766 0 235826 580 6 um_iw[217]
port 211 nsew signal output
rlabel metal4 s 235030 0 235090 1124 6 um_iw[218]
port 212 nsew signal output
rlabel metal4 s 234294 0 234354 580 6 um_iw[219]
port 213 nsew signal output
rlabel metal4 s 29502 9756 29562 10880 6 um_iw[21]
port 214 nsew signal output
rlabel metal4 s 233558 0 233618 580 6 um_iw[220]
port 215 nsew signal output
rlabel metal4 s 232822 0 232882 1124 6 um_iw[221]
port 216 nsew signal output
rlabel metal4 s 232086 0 232146 1124 6 um_iw[222]
port 217 nsew signal output
rlabel metal4 s 231350 0 231410 580 6 um_iw[223]
port 218 nsew signal output
rlabel metal4 s 230614 0 230674 1124 6 um_iw[224]
port 219 nsew signal output
rlabel metal4 s 229878 0 229938 1124 6 um_iw[225]
port 220 nsew signal output
rlabel metal4 s 229142 0 229202 580 6 um_iw[226]
port 221 nsew signal output
rlabel metal4 s 228406 0 228466 580 6 um_iw[227]
port 222 nsew signal output
rlabel metal4 s 227670 0 227730 1124 6 um_iw[228]
port 223 nsew signal output
rlabel metal4 s 226934 0 226994 580 6 um_iw[229]
port 224 nsew signal output
rlabel metal4 s 28766 8668 28826 10880 6 um_iw[22]
port 225 nsew signal output
rlabel metal4 s 226198 0 226258 1396 6 um_iw[230]
port 226 nsew signal output
rlabel metal4 s 225462 0 225522 1124 6 um_iw[231]
port 227 nsew signal output
rlabel metal4 s 224726 0 224786 716 6 um_iw[232]
port 228 nsew signal output
rlabel metal4 s 223990 0 224050 1124 6 um_iw[233]
port 229 nsew signal output
rlabel metal4 s 236502 9212 236562 10880 6 um_iw[234]
port 230 nsew signal output
rlabel metal4 s 235766 9484 235826 10880 6 um_iw[235]
port 231 nsew signal output
rlabel metal4 s 235030 8396 235090 10880 6 um_iw[236]
port 232 nsew signal output
rlabel metal4 s 234294 8668 234354 10880 6 um_iw[237]
port 233 nsew signal output
rlabel metal4 s 233558 9484 233618 10880 6 um_iw[238]
port 234 nsew signal output
rlabel metal4 s 232822 8668 232882 10880 6 um_iw[239]
port 235 nsew signal output
rlabel metal4 s 28030 8668 28090 10880 6 um_iw[23]
port 236 nsew signal output
rlabel metal4 s 232086 9484 232146 10880 6 um_iw[240]
port 237 nsew signal output
rlabel metal4 s 231350 8668 231410 10880 6 um_iw[241]
port 238 nsew signal output
rlabel metal4 s 230614 8668 230674 10880 6 um_iw[242]
port 239 nsew signal output
rlabel metal4 s 229878 9484 229938 10880 6 um_iw[243]
port 240 nsew signal output
rlabel metal4 s 229142 8668 229202 10880 6 um_iw[244]
port 241 nsew signal output
rlabel metal4 s 228406 9484 228466 10880 6 um_iw[245]
port 242 nsew signal output
rlabel metal4 s 227670 9484 227730 10880 6 um_iw[246]
port 243 nsew signal output
rlabel metal4 s 226934 8668 226994 10880 6 um_iw[247]
port 244 nsew signal output
rlabel metal4 s 226198 8668 226258 10880 6 um_iw[248]
port 245 nsew signal output
rlabel metal4 s 225462 8668 225522 10880 6 um_iw[249]
port 246 nsew signal output
rlabel metal4 s 27294 8668 27354 10880 6 um_iw[24]
port 247 nsew signal output
rlabel metal4 s 224726 8668 224786 10880 6 um_iw[250]
port 248 nsew signal output
rlabel metal4 s 223990 9484 224050 10880 6 um_iw[251]
port 249 nsew signal output
rlabel metal4 s 270634 0 270694 580 6 um_iw[252]
port 250 nsew signal output
rlabel metal4 s 269898 0 269958 308 6 um_iw[253]
port 251 nsew signal output
rlabel metal4 s 269162 0 269222 580 6 um_iw[254]
port 252 nsew signal output
rlabel metal4 s 268426 0 268486 580 6 um_iw[255]
port 253 nsew signal output
rlabel metal4 s 267690 0 267750 580 6 um_iw[256]
port 254 nsew signal output
rlabel metal4 s 266954 0 267014 580 6 um_iw[257]
port 255 nsew signal output
rlabel metal4 s 266218 0 266278 580 6 um_iw[258]
port 256 nsew signal output
rlabel metal4 s 265482 0 265542 580 6 um_iw[259]
port 257 nsew signal output
rlabel metal4 s 26558 9756 26618 10880 6 um_iw[25]
port 258 nsew signal output
rlabel metal4 s 264746 0 264806 580 6 um_iw[260]
port 259 nsew signal output
rlabel metal4 s 264010 0 264070 580 6 um_iw[261]
port 260 nsew signal output
rlabel metal4 s 263274 0 263334 580 6 um_iw[262]
port 261 nsew signal output
rlabel metal4 s 262538 0 262598 580 6 um_iw[263]
port 262 nsew signal output
rlabel metal4 s 261802 0 261862 642 6 um_iw[264]
port 263 nsew signal output
rlabel metal4 s 261066 0 261126 580 6 um_iw[265]
port 264 nsew signal output
rlabel metal4 s 260330 0 260390 642 6 um_iw[266]
port 265 nsew signal output
rlabel metal4 s 259594 0 259654 642 6 um_iw[267]
port 266 nsew signal output
rlabel metal4 s 258858 0 258918 642 6 um_iw[268]
port 267 nsew signal output
rlabel metal4 s 258122 0 258182 580 6 um_iw[269]
port 268 nsew signal output
rlabel metal4 s 25822 9756 25882 10880 6 um_iw[26]
port 269 nsew signal output
rlabel metal4 s 270634 10238 270694 10880 6 um_iw[270]
port 270 nsew signal output
rlabel metal4 s 269898 10238 269958 10880 6 um_iw[271]
port 271 nsew signal output
rlabel metal4 s 269162 10238 269222 10880 6 um_iw[272]
port 272 nsew signal output
rlabel metal4 s 268426 10238 268486 10880 6 um_iw[273]
port 273 nsew signal output
rlabel metal4 s 267690 10238 267750 10880 6 um_iw[274]
port 274 nsew signal output
rlabel metal4 s 266954 10238 267014 10880 6 um_iw[275]
port 275 nsew signal output
rlabel metal4 s 266218 10300 266278 10880 6 um_iw[276]
port 276 nsew signal output
rlabel metal4 s 265482 10436 265542 10880 6 um_iw[277]
port 277 nsew signal output
rlabel metal4 s 264746 10238 264806 10880 6 um_iw[278]
port 278 nsew signal output
rlabel metal4 s 264010 10300 264070 10880 6 um_iw[279]
port 279 nsew signal output
rlabel metal4 s 25086 8396 25146 10880 6 um_iw[27]
port 280 nsew signal output
rlabel metal4 s 263274 10300 263334 10880 6 um_iw[280]
port 281 nsew signal output
rlabel metal4 s 262538 10300 262598 10880 6 um_iw[281]
port 282 nsew signal output
rlabel metal4 s 261802 10300 261862 10880 6 um_iw[282]
port 283 nsew signal output
rlabel metal4 s 261066 10436 261126 10880 6 um_iw[283]
port 284 nsew signal output
rlabel metal4 s 260330 10300 260390 10880 6 um_iw[284]
port 285 nsew signal output
rlabel metal4 s 259594 10300 259654 10880 6 um_iw[285]
port 286 nsew signal output
rlabel metal4 s 258858 10300 258918 10880 6 um_iw[286]
port 287 nsew signal output
rlabel metal4 s 258122 10300 258182 10880 6 um_iw[287]
port 288 nsew signal output
rlabel metal4 s 24350 9212 24410 10880 6 um_iw[28]
port 289 nsew signal output
rlabel metal4 s 23614 8396 23674 10880 6 um_iw[29]
port 290 nsew signal output
rlabel metal4 s 30238 0 30298 580 6 um_iw[2]
port 291 nsew signal output
rlabel metal4 s 22878 8396 22938 10880 6 um_iw[30]
port 292 nsew signal output
rlabel metal4 s 22142 8940 22202 10880 6 um_iw[31]
port 293 nsew signal output
rlabel metal4 s 21406 8668 21466 10880 6 um_iw[32]
port 294 nsew signal output
rlabel metal4 s 20670 8396 20730 10880 6 um_iw[33]
port 295 nsew signal output
rlabel metal4 s 19934 9892 19994 10880 6 um_iw[34]
port 296 nsew signal output
rlabel metal4 s 19198 6900 19258 10880 6 um_iw[35]
port 297 nsew signal output
rlabel metal4 s 65842 0 65902 444 6 um_iw[36]
port 298 nsew signal output
rlabel metal4 s 65106 0 65166 308 6 um_iw[37]
port 299 nsew signal output
rlabel metal4 s 64370 0 64430 308 6 um_iw[38]
port 300 nsew signal output
rlabel metal4 s 63634 0 63694 308 6 um_iw[39]
port 301 nsew signal output
rlabel metal4 s 29502 0 29562 1124 6 um_iw[3]
port 302 nsew signal output
rlabel metal4 s 62898 0 62958 444 6 um_iw[40]
port 303 nsew signal output
rlabel metal4 s 62162 0 62222 444 6 um_iw[41]
port 304 nsew signal output
rlabel metal4 s 61426 0 61486 444 6 um_iw[42]
port 305 nsew signal output
rlabel metal4 s 60690 0 60750 444 6 um_iw[43]
port 306 nsew signal output
rlabel metal4 s 59954 0 60014 444 6 um_iw[44]
port 307 nsew signal output
rlabel metal4 s 59218 0 59278 370 6 um_iw[45]
port 308 nsew signal output
rlabel metal4 s 58482 0 58542 444 6 um_iw[46]
port 309 nsew signal output
rlabel metal4 s 57746 0 57806 370 6 um_iw[47]
port 310 nsew signal output
rlabel metal4 s 57010 0 57070 444 6 um_iw[48]
port 311 nsew signal output
rlabel metal4 s 56274 0 56334 444 6 um_iw[49]
port 312 nsew signal output
rlabel metal4 s 28766 0 28826 308 6 um_iw[4]
port 313 nsew signal output
rlabel metal4 s 55538 0 55598 444 6 um_iw[50]
port 314 nsew signal output
rlabel metal4 s 54802 0 54862 370 6 um_iw[51]
port 315 nsew signal output
rlabel metal4 s 54066 0 54126 580 6 um_iw[52]
port 316 nsew signal output
rlabel metal4 s 53330 0 53390 580 6 um_iw[53]
port 317 nsew signal output
rlabel metal4 s 65842 10300 65902 10880 6 um_iw[54]
port 318 nsew signal output
rlabel metal4 s 65106 10300 65166 10880 6 um_iw[55]
port 319 nsew signal output
rlabel metal4 s 64370 10300 64430 10880 6 um_iw[56]
port 320 nsew signal output
rlabel metal4 s 63634 10300 63694 10880 6 um_iw[57]
port 321 nsew signal output
rlabel metal4 s 62898 10300 62958 10880 6 um_iw[58]
port 322 nsew signal output
rlabel metal4 s 62162 10300 62222 10880 6 um_iw[59]
port 323 nsew signal output
rlabel metal4 s 28030 0 28090 580 6 um_iw[5]
port 324 nsew signal output
rlabel metal4 s 61426 10300 61486 10880 6 um_iw[60]
port 325 nsew signal output
rlabel metal4 s 60690 10300 60750 10880 6 um_iw[61]
port 326 nsew signal output
rlabel metal4 s 59954 10300 60014 10880 6 um_iw[62]
port 327 nsew signal output
rlabel metal4 s 59218 10300 59278 10880 6 um_iw[63]
port 328 nsew signal output
rlabel metal4 s 58482 10300 58542 10880 6 um_iw[64]
port 329 nsew signal output
rlabel metal4 s 57746 10300 57806 10880 6 um_iw[65]
port 330 nsew signal output
rlabel metal4 s 57010 10300 57070 10880 6 um_iw[66]
port 331 nsew signal output
rlabel metal4 s 56274 10300 56334 10880 6 um_iw[67]
port 332 nsew signal output
rlabel metal4 s 55538 10300 55598 10880 6 um_iw[68]
port 333 nsew signal output
rlabel metal4 s 54802 10300 54862 10880 6 um_iw[69]
port 334 nsew signal output
rlabel metal4 s 27294 0 27354 2756 6 um_iw[6]
port 335 nsew signal output
rlabel metal4 s 54066 10300 54126 10880 6 um_iw[70]
port 336 nsew signal output
rlabel metal4 s 53330 10300 53390 10880 6 um_iw[71]
port 337 nsew signal output
rlabel metal4 s 99974 0 100034 580 6 um_iw[72]
port 338 nsew signal output
rlabel metal4 s 99238 0 99298 852 6 um_iw[73]
port 339 nsew signal output
rlabel metal4 s 98502 0 98562 1532 6 um_iw[74]
port 340 nsew signal output
rlabel metal4 s 97766 0 97826 3708 6 um_iw[75]
port 341 nsew signal output
rlabel metal4 s 97030 0 97090 2756 6 um_iw[76]
port 342 nsew signal output
rlabel metal4 s 96294 0 96354 1532 6 um_iw[77]
port 343 nsew signal output
rlabel metal4 s 95558 0 95618 2756 6 um_iw[78]
port 344 nsew signal output
rlabel metal4 s 94822 0 94882 580 6 um_iw[79]
port 345 nsew signal output
rlabel metal4 s 26558 0 26618 1260 6 um_iw[7]
port 346 nsew signal output
rlabel metal4 s 94086 0 94146 3028 6 um_iw[80]
port 347 nsew signal output
rlabel metal4 s 93350 0 93410 1260 6 um_iw[81]
port 348 nsew signal output
rlabel metal4 s 92614 0 92674 580 6 um_iw[82]
port 349 nsew signal output
rlabel metal4 s 91878 0 91938 1260 6 um_iw[83]
port 350 nsew signal output
rlabel metal4 s 91142 0 91202 1532 6 um_iw[84]
port 351 nsew signal output
rlabel metal4 s 90406 0 90466 1260 6 um_iw[85]
port 352 nsew signal output
rlabel metal4 s 89670 0 89730 370 6 um_iw[86]
port 353 nsew signal output
rlabel metal4 s 88934 0 88994 1260 6 um_iw[87]
port 354 nsew signal output
rlabel metal4 s 88198 0 88258 1396 6 um_iw[88]
port 355 nsew signal output
rlabel metal4 s 87462 0 87522 444 6 um_iw[89]
port 356 nsew signal output
rlabel metal4 s 25822 0 25882 1260 6 um_iw[8]
port 357 nsew signal output
rlabel metal4 s 99974 9756 100034 10880 6 um_iw[90]
port 358 nsew signal output
rlabel metal4 s 99238 8668 99298 10880 6 um_iw[91]
port 359 nsew signal output
rlabel metal4 s 98502 9756 98562 10880 6 um_iw[92]
port 360 nsew signal output
rlabel metal4 s 97766 8668 97826 10880 6 um_iw[93]
port 361 nsew signal output
rlabel metal4 s 97030 8668 97090 10880 6 um_iw[94]
port 362 nsew signal output
rlabel metal4 s 96294 9756 96354 10880 6 um_iw[95]
port 363 nsew signal output
rlabel metal4 s 95558 9756 95618 10880 6 um_iw[96]
port 364 nsew signal output
rlabel metal4 s 94822 8668 94882 10880 6 um_iw[97]
port 365 nsew signal output
rlabel metal4 s 94086 8668 94146 10880 6 um_iw[98]
port 366 nsew signal output
rlabel metal4 s 93350 9756 93410 10880 6 um_iw[99]
port 367 nsew signal output
rlabel metal4 s 25086 0 25146 2756 6 um_iw[9]
port 368 nsew signal output
rlabel metal4 s 798 0 858 2756 6 um_k_zero[0]
port 369 nsew signal output
rlabel metal4 s 171458 0 171518 580 6 um_k_zero[10]
port 370 nsew signal output
rlabel metal4 s 171458 10300 171518 10880 6 um_k_zero[11]
port 371 nsew signal output
rlabel metal4 s 205590 0 205650 852 6 um_k_zero[12]
port 372 nsew signal output
rlabel metal4 s 205590 10300 205650 10880 6 um_k_zero[13]
port 373 nsew signal output
rlabel metal4 s 239722 0 239782 580 6 um_k_zero[14]
port 374 nsew signal output
rlabel metal4 s 239722 10300 239782 10880 6 um_k_zero[15]
port 375 nsew signal output
rlabel metal4 s 798 9212 858 10880 6 um_k_zero[1]
port 376 nsew signal output
rlabel metal4 s 34930 0 34990 580 6 um_k_zero[2]
port 377 nsew signal output
rlabel metal4 s 34930 10300 34990 10880 6 um_k_zero[3]
port 378 nsew signal output
rlabel metal4 s 69062 0 69122 852 6 um_k_zero[4]
port 379 nsew signal output
rlabel metal4 s 69062 9620 69122 10880 6 um_k_zero[5]
port 380 nsew signal output
rlabel metal4 s 103194 0 103254 370 6 um_k_zero[6]
port 381 nsew signal output
rlabel metal4 s 103194 10300 103254 10880 6 um_k_zero[7]
port 382 nsew signal output
rlabel metal4 s 137326 0 137386 1396 6 um_k_zero[8]
port 383 nsew signal output
rlabel metal4 s 137326 9620 137386 10880 6 um_k_zero[9]
port 384 nsew signal output
rlabel metal4 s 18462 0 18522 308 6 um_ow[0]
port 385 nsew signal input
rlabel metal4 s 83782 0 83842 1260 6 um_ow[100]
port 386 nsew signal input
rlabel metal4 s 83046 0 83106 852 6 um_ow[101]
port 387 nsew signal input
rlabel metal4 s 82310 0 82370 988 6 um_ow[102]
port 388 nsew signal input
rlabel metal4 s 81574 0 81634 1260 6 um_ow[103]
port 389 nsew signal input
rlabel metal4 s 80838 0 80898 988 6 um_ow[104]
port 390 nsew signal input
rlabel metal4 s 80102 0 80162 852 6 um_ow[105]
port 391 nsew signal input
rlabel metal4 s 79366 0 79426 988 6 um_ow[106]
port 392 nsew signal input
rlabel metal4 s 78630 0 78690 1260 6 um_ow[107]
port 393 nsew signal input
rlabel metal4 s 77894 0 77954 852 6 um_ow[108]
port 394 nsew signal input
rlabel metal4 s 77158 0 77218 988 6 um_ow[109]
port 395 nsew signal input
rlabel metal4 s 11102 0 11162 716 6 um_ow[10]
port 396 nsew signal input
rlabel metal4 s 76422 0 76482 1260 6 um_ow[110]
port 397 nsew signal input
rlabel metal4 s 75686 0 75746 988 6 um_ow[111]
port 398 nsew signal input
rlabel metal4 s 74950 0 75010 852 6 um_ow[112]
port 399 nsew signal input
rlabel metal4 s 74214 0 74274 852 6 um_ow[113]
port 400 nsew signal input
rlabel metal4 s 73478 0 73538 988 6 um_ow[114]
port 401 nsew signal input
rlabel metal4 s 72742 0 72802 852 6 um_ow[115]
port 402 nsew signal input
rlabel metal4 s 72006 0 72066 988 6 um_ow[116]
port 403 nsew signal input
rlabel metal4 s 71270 0 71330 988 6 um_ow[117]
port 404 nsew signal input
rlabel metal4 s 70534 0 70594 852 6 um_ow[118]
port 405 nsew signal input
rlabel metal4 s 69798 0 69858 852 6 um_ow[119]
port 406 nsew signal input
rlabel metal4 s 10366 0 10426 716 6 um_ow[11]
port 407 nsew signal input
rlabel metal4 s 86726 10572 86786 10880 6 um_ow[120]
port 408 nsew signal input
rlabel metal4 s 85990 9892 86050 10880 6 um_ow[121]
port 409 nsew signal input
rlabel metal4 s 85254 10164 85314 10880 6 um_ow[122]
port 410 nsew signal input
rlabel metal4 s 84518 10164 84578 10880 6 um_ow[123]
port 411 nsew signal input
rlabel metal4 s 83782 10164 83842 10880 6 um_ow[124]
port 412 nsew signal input
rlabel metal4 s 83046 10164 83106 10880 6 um_ow[125]
port 413 nsew signal input
rlabel metal4 s 82310 10572 82370 10880 6 um_ow[126]
port 414 nsew signal input
rlabel metal4 s 81574 10572 81634 10880 6 um_ow[127]
port 415 nsew signal input
rlabel metal4 s 80838 9892 80898 10880 6 um_ow[128]
port 416 nsew signal input
rlabel metal4 s 80102 9620 80162 10880 6 um_ow[129]
port 417 nsew signal input
rlabel metal4 s 9630 0 9690 988 6 um_ow[12]
port 418 nsew signal input
rlabel metal4 s 79366 10164 79426 10880 6 um_ow[130]
port 419 nsew signal input
rlabel metal4 s 78630 9892 78690 10880 6 um_ow[131]
port 420 nsew signal input
rlabel metal4 s 77894 9620 77954 10880 6 um_ow[132]
port 421 nsew signal input
rlabel metal4 s 77158 9892 77218 10880 6 um_ow[133]
port 422 nsew signal input
rlabel metal4 s 76422 9620 76482 10880 6 um_ow[134]
port 423 nsew signal input
rlabel metal4 s 75686 9620 75746 10880 6 um_ow[135]
port 424 nsew signal input
rlabel metal4 s 74950 9076 75010 10880 6 um_ow[136]
port 425 nsew signal input
rlabel metal4 s 74214 9620 74274 10880 6 um_ow[137]
port 426 nsew signal input
rlabel metal4 s 73478 9076 73538 10880 6 um_ow[138]
port 427 nsew signal input
rlabel metal4 s 72742 9620 72802 10880 6 um_ow[139]
port 428 nsew signal input
rlabel metal4 s 8894 0 8954 308 6 um_ow[13]
port 429 nsew signal input
rlabel metal4 s 72006 10436 72066 10880 6 um_ow[140]
port 430 nsew signal input
rlabel metal4 s 71270 10164 71330 10880 6 um_ow[141]
port 431 nsew signal input
rlabel metal4 s 70534 9620 70594 10880 6 um_ow[142]
port 432 nsew signal input
rlabel metal4 s 69798 9892 69858 10880 6 um_ow[143]
port 433 nsew signal input
rlabel metal4 s 120858 0 120918 444 6 um_ow[144]
port 434 nsew signal input
rlabel metal4 s 120122 0 120182 444 6 um_ow[145]
port 435 nsew signal input
rlabel metal4 s 119386 0 119446 444 6 um_ow[146]
port 436 nsew signal input
rlabel metal4 s 118650 0 118710 444 6 um_ow[147]
port 437 nsew signal input
rlabel metal4 s 117914 0 117974 444 6 um_ow[148]
port 438 nsew signal input
rlabel metal4 s 117178 0 117238 370 6 um_ow[149]
port 439 nsew signal input
rlabel metal4 s 8158 0 8218 444 6 um_ow[14]
port 440 nsew signal input
rlabel metal4 s 116442 0 116502 370 6 um_ow[150]
port 441 nsew signal input
rlabel metal4 s 115706 0 115766 370 6 um_ow[151]
port 442 nsew signal input
rlabel metal4 s 114970 0 115030 370 6 um_ow[152]
port 443 nsew signal input
rlabel metal4 s 114234 0 114294 370 6 um_ow[153]
port 444 nsew signal input
rlabel metal4 s 113498 0 113558 370 6 um_ow[154]
port 445 nsew signal input
rlabel metal4 s 112762 0 112822 370 6 um_ow[155]
port 446 nsew signal input
rlabel metal4 s 112026 0 112086 370 6 um_ow[156]
port 447 nsew signal input
rlabel metal4 s 111290 0 111350 370 6 um_ow[157]
port 448 nsew signal input
rlabel metal4 s 110554 0 110614 370 6 um_ow[158]
port 449 nsew signal input
rlabel metal4 s 109818 0 109878 370 6 um_ow[159]
port 450 nsew signal input
rlabel metal4 s 7422 0 7482 988 6 um_ow[15]
port 451 nsew signal input
rlabel metal4 s 109082 0 109142 370 6 um_ow[160]
port 452 nsew signal input
rlabel metal4 s 108346 0 108406 370 6 um_ow[161]
port 453 nsew signal input
rlabel metal4 s 107610 0 107670 370 6 um_ow[162]
port 454 nsew signal input
rlabel metal4 s 106874 0 106934 370 6 um_ow[163]
port 455 nsew signal input
rlabel metal4 s 106138 0 106198 370 6 um_ow[164]
port 456 nsew signal input
rlabel metal4 s 105402 0 105462 370 6 um_ow[165]
port 457 nsew signal input
rlabel metal4 s 104666 0 104726 370 6 um_ow[166]
port 458 nsew signal input
rlabel metal4 s 103930 0 103990 370 6 um_ow[167]
port 459 nsew signal input
rlabel metal4 s 120858 10300 120918 10880 6 um_ow[168]
port 460 nsew signal input
rlabel metal4 s 120122 10300 120182 10880 6 um_ow[169]
port 461 nsew signal input
rlabel metal4 s 6686 0 6746 1260 6 um_ow[16]
port 462 nsew signal input
rlabel metal4 s 119386 10300 119446 10880 6 um_ow[170]
port 463 nsew signal input
rlabel metal4 s 118650 10300 118710 10880 6 um_ow[171]
port 464 nsew signal input
rlabel metal4 s 117914 10300 117974 10880 6 um_ow[172]
port 465 nsew signal input
rlabel metal4 s 117178 10300 117238 10880 6 um_ow[173]
port 466 nsew signal input
rlabel metal4 s 116442 10300 116502 10880 6 um_ow[174]
port 467 nsew signal input
rlabel metal4 s 115706 10300 115766 10880 6 um_ow[175]
port 468 nsew signal input
rlabel metal4 s 114970 10300 115030 10880 6 um_ow[176]
port 469 nsew signal input
rlabel metal4 s 114234 10300 114294 10880 6 um_ow[177]
port 470 nsew signal input
rlabel metal4 s 113498 10300 113558 10880 6 um_ow[178]
port 471 nsew signal input
rlabel metal4 s 112762 10300 112822 10880 6 um_ow[179]
port 472 nsew signal input
rlabel metal4 s 5950 0 6010 716 6 um_ow[17]
port 473 nsew signal input
rlabel metal4 s 112026 10300 112086 10880 6 um_ow[180]
port 474 nsew signal input
rlabel metal4 s 111290 10300 111350 10880 6 um_ow[181]
port 475 nsew signal input
rlabel metal4 s 110554 10300 110614 10880 6 um_ow[182]
port 476 nsew signal input
rlabel metal4 s 109818 10300 109878 10880 6 um_ow[183]
port 477 nsew signal input
rlabel metal4 s 109082 10300 109142 10880 6 um_ow[184]
port 478 nsew signal input
rlabel metal4 s 108346 10300 108406 10880 6 um_ow[185]
port 479 nsew signal input
rlabel metal4 s 107610 10300 107670 10880 6 um_ow[186]
port 480 nsew signal input
rlabel metal4 s 106874 10300 106934 10880 6 um_ow[187]
port 481 nsew signal input
rlabel metal4 s 106138 10300 106198 10880 6 um_ow[188]
port 482 nsew signal input
rlabel metal4 s 105402 10300 105462 10880 6 um_ow[189]
port 483 nsew signal input
rlabel metal4 s 5214 0 5274 988 6 um_ow[18]
port 484 nsew signal input
rlabel metal4 s 104666 10300 104726 10880 6 um_ow[190]
port 485 nsew signal input
rlabel metal4 s 103930 10300 103990 10880 6 um_ow[191]
port 486 nsew signal input
rlabel metal4 s 154990 0 155050 2892 6 um_ow[192]
port 487 nsew signal input
rlabel metal4 s 154254 0 154314 3300 6 um_ow[193]
port 488 nsew signal input
rlabel metal4 s 153518 0 153578 2892 6 um_ow[194]
port 489 nsew signal input
rlabel metal4 s 152782 0 152842 1260 6 um_ow[195]
port 490 nsew signal input
rlabel metal4 s 152046 0 152106 1396 6 um_ow[196]
port 491 nsew signal input
rlabel metal4 s 151310 0 151370 580 6 um_ow[197]
port 492 nsew signal input
rlabel metal4 s 150574 0 150634 1396 6 um_ow[198]
port 493 nsew signal input
rlabel metal4 s 149838 0 149898 716 6 um_ow[199]
port 494 nsew signal input
rlabel metal4 s 4478 0 4538 1260 6 um_ow[19]
port 495 nsew signal input
rlabel metal4 s 17726 0 17786 988 6 um_ow[1]
port 496 nsew signal input
rlabel metal4 s 149102 0 149162 2892 6 um_ow[200]
port 497 nsew signal input
rlabel metal4 s 148366 0 148426 716 6 um_ow[201]
port 498 nsew signal input
rlabel metal4 s 147630 0 147690 580 6 um_ow[202]
port 499 nsew signal input
rlabel metal4 s 146894 0 146954 308 6 um_ow[203]
port 500 nsew signal input
rlabel metal4 s 146158 0 146218 716 6 um_ow[204]
port 501 nsew signal input
rlabel metal4 s 145422 0 145482 2756 6 um_ow[205]
port 502 nsew signal input
rlabel metal4 s 144686 0 144746 3164 6 um_ow[206]
port 503 nsew signal input
rlabel metal4 s 143950 0 144010 444 6 um_ow[207]
port 504 nsew signal input
rlabel metal4 s 143214 0 143274 580 6 um_ow[208]
port 505 nsew signal input
rlabel metal4 s 142478 0 142538 716 6 um_ow[209]
port 506 nsew signal input
rlabel metal4 s 3742 0 3802 988 6 um_ow[20]
port 507 nsew signal input
rlabel metal4 s 141742 0 141802 716 6 um_ow[210]
port 508 nsew signal input
rlabel metal4 s 141006 0 141066 1396 6 um_ow[211]
port 509 nsew signal input
rlabel metal4 s 140270 0 140330 1804 6 um_ow[212]
port 510 nsew signal input
rlabel metal4 s 139534 0 139594 988 6 um_ow[213]
port 511 nsew signal input
rlabel metal4 s 138798 0 138858 716 6 um_ow[214]
port 512 nsew signal input
rlabel metal4 s 138062 0 138122 580 6 um_ow[215]
port 513 nsew signal input
rlabel metal4 s 154990 9892 155050 10880 6 um_ow[216]
port 514 nsew signal input
rlabel metal4 s 154254 10436 154314 10880 6 um_ow[217]
port 515 nsew signal input
rlabel metal4 s 153518 10164 153578 10880 6 um_ow[218]
port 516 nsew signal input
rlabel metal4 s 152782 10164 152842 10880 6 um_ow[219]
port 517 nsew signal input
rlabel metal4 s 3006 0 3066 716 6 um_ow[21]
port 518 nsew signal input
rlabel metal4 s 152046 10164 152106 10880 6 um_ow[220]
port 519 nsew signal input
rlabel metal4 s 151310 10164 151370 10880 6 um_ow[221]
port 520 nsew signal input
rlabel metal4 s 150574 10164 150634 10880 6 um_ow[222]
port 521 nsew signal input
rlabel metal4 s 149838 9892 149898 10880 6 um_ow[223]
port 522 nsew signal input
rlabel metal4 s 149102 10164 149162 10880 6 um_ow[224]
port 523 nsew signal input
rlabel metal4 s 148366 10300 148426 10880 6 um_ow[225]
port 524 nsew signal input
rlabel metal4 s 147630 10572 147690 10880 6 um_ow[226]
port 525 nsew signal input
rlabel metal4 s 146894 10164 146954 10880 6 um_ow[227]
port 526 nsew signal input
rlabel metal4 s 146158 10164 146218 10880 6 um_ow[228]
port 527 nsew signal input
rlabel metal4 s 145422 10164 145482 10880 6 um_ow[229]
port 528 nsew signal input
rlabel metal4 s 2270 0 2330 580 6 um_ow[22]
port 529 nsew signal input
rlabel metal4 s 144686 9892 144746 10880 6 um_ow[230]
port 530 nsew signal input
rlabel metal4 s 143950 10164 144010 10880 6 um_ow[231]
port 531 nsew signal input
rlabel metal4 s 143214 10164 143274 10880 6 um_ow[232]
port 532 nsew signal input
rlabel metal4 s 142478 10300 142538 10880 6 um_ow[233]
port 533 nsew signal input
rlabel metal4 s 141742 10164 141802 10880 6 um_ow[234]
port 534 nsew signal input
rlabel metal4 s 141006 10164 141066 10880 6 um_ow[235]
port 535 nsew signal input
rlabel metal4 s 140270 10164 140330 10880 6 um_ow[236]
port 536 nsew signal input
rlabel metal4 s 139534 9892 139594 10880 6 um_ow[237]
port 537 nsew signal input
rlabel metal4 s 138798 10164 138858 10880 6 um_ow[238]
port 538 nsew signal input
rlabel metal4 s 138062 10300 138122 10880 6 um_ow[239]
port 539 nsew signal input
rlabel metal4 s 1534 0 1594 988 6 um_ow[23]
port 540 nsew signal input
rlabel metal4 s 189122 0 189182 444 6 um_ow[240]
port 541 nsew signal input
rlabel metal4 s 188386 0 188446 444 6 um_ow[241]
port 542 nsew signal input
rlabel metal4 s 187650 0 187710 444 6 um_ow[242]
port 543 nsew signal input
rlabel metal4 s 186914 0 186974 444 6 um_ow[243]
port 544 nsew signal input
rlabel metal4 s 186178 0 186238 370 6 um_ow[244]
port 545 nsew signal input
rlabel metal4 s 185442 0 185502 444 6 um_ow[245]
port 546 nsew signal input
rlabel metal4 s 184706 0 184766 444 6 um_ow[246]
port 547 nsew signal input
rlabel metal4 s 183970 0 184030 444 6 um_ow[247]
port 548 nsew signal input
rlabel metal4 s 183234 0 183294 444 6 um_ow[248]
port 549 nsew signal input
rlabel metal4 s 182498 0 182558 444 6 um_ow[249]
port 550 nsew signal input
rlabel metal4 s 18462 10164 18522 10880 6 um_ow[24]
port 551 nsew signal input
rlabel metal4 s 181762 0 181822 444 6 um_ow[250]
port 552 nsew signal input
rlabel metal4 s 181026 0 181086 308 6 um_ow[251]
port 553 nsew signal input
rlabel metal4 s 180290 0 180350 580 6 um_ow[252]
port 554 nsew signal input
rlabel metal4 s 179554 0 179614 580 6 um_ow[253]
port 555 nsew signal input
rlabel metal4 s 178818 0 178878 580 6 um_ow[254]
port 556 nsew signal input
rlabel metal4 s 178082 0 178142 580 6 um_ow[255]
port 557 nsew signal input
rlabel metal4 s 177346 0 177406 580 6 um_ow[256]
port 558 nsew signal input
rlabel metal4 s 176610 0 176670 580 6 um_ow[257]
port 559 nsew signal input
rlabel metal4 s 175874 0 175934 444 6 um_ow[258]
port 560 nsew signal input
rlabel metal4 s 175138 0 175198 580 6 um_ow[259]
port 561 nsew signal input
rlabel metal4 s 17726 10164 17786 10880 6 um_ow[25]
port 562 nsew signal input
rlabel metal4 s 174402 0 174462 580 6 um_ow[260]
port 563 nsew signal input
rlabel metal4 s 173666 0 173726 580 6 um_ow[261]
port 564 nsew signal input
rlabel metal4 s 172930 0 172990 580 6 um_ow[262]
port 565 nsew signal input
rlabel metal4 s 172194 0 172254 580 6 um_ow[263]
port 566 nsew signal input
rlabel metal4 s 189122 10300 189182 10880 6 um_ow[264]
port 567 nsew signal input
rlabel metal4 s 188386 10300 188446 10880 6 um_ow[265]
port 568 nsew signal input
rlabel metal4 s 187650 10300 187710 10880 6 um_ow[266]
port 569 nsew signal input
rlabel metal4 s 186914 10300 186974 10880 6 um_ow[267]
port 570 nsew signal input
rlabel metal4 s 186178 10300 186238 10880 6 um_ow[268]
port 571 nsew signal input
rlabel metal4 s 185442 10300 185502 10880 6 um_ow[269]
port 572 nsew signal input
rlabel metal4 s 16990 10164 17050 10880 6 um_ow[26]
port 573 nsew signal input
rlabel metal4 s 184706 10300 184766 10880 6 um_ow[270]
port 574 nsew signal input
rlabel metal4 s 183970 10300 184030 10880 6 um_ow[271]
port 575 nsew signal input
rlabel metal4 s 183234 10300 183294 10880 6 um_ow[272]
port 576 nsew signal input
rlabel metal4 s 182498 10300 182558 10880 6 um_ow[273]
port 577 nsew signal input
rlabel metal4 s 181762 10300 181822 10880 6 um_ow[274]
port 578 nsew signal input
rlabel metal4 s 181026 10436 181086 10880 6 um_ow[275]
port 579 nsew signal input
rlabel metal4 s 180290 10300 180350 10880 6 um_ow[276]
port 580 nsew signal input
rlabel metal4 s 179554 10572 179614 10880 6 um_ow[277]
port 581 nsew signal input
rlabel metal4 s 178818 10300 178878 10880 6 um_ow[278]
port 582 nsew signal input
rlabel metal4 s 178082 10300 178142 10880 6 um_ow[279]
port 583 nsew signal input
rlabel metal4 s 16254 10164 16314 10880 6 um_ow[27]
port 584 nsew signal input
rlabel metal4 s 177346 10300 177406 10880 6 um_ow[280]
port 585 nsew signal input
rlabel metal4 s 176610 10300 176670 10880 6 um_ow[281]
port 586 nsew signal input
rlabel metal4 s 175874 10300 175934 10880 6 um_ow[282]
port 587 nsew signal input
rlabel metal4 s 175138 10300 175198 10880 6 um_ow[283]
port 588 nsew signal input
rlabel metal4 s 174402 10300 174462 10880 6 um_ow[284]
port 589 nsew signal input
rlabel metal4 s 173666 10300 173726 10880 6 um_ow[285]
port 590 nsew signal input
rlabel metal4 s 172930 10436 172990 10880 6 um_ow[286]
port 591 nsew signal input
rlabel metal4 s 172194 10572 172254 10880 6 um_ow[287]
port 592 nsew signal input
rlabel metal4 s 223254 0 223314 3708 6 um_ow[288]
port 593 nsew signal input
rlabel metal4 s 222518 0 222578 1396 6 um_ow[289]
port 594 nsew signal input
rlabel metal4 s 15518 10164 15578 10880 6 um_ow[28]
port 595 nsew signal input
rlabel metal4 s 221782 0 221842 580 6 um_ow[290]
port 596 nsew signal input
rlabel metal4 s 221046 0 221106 3164 6 um_ow[291]
port 597 nsew signal input
rlabel metal4 s 220310 0 220370 308 6 um_ow[292]
port 598 nsew signal input
rlabel metal4 s 219574 0 219634 1396 6 um_ow[293]
port 599 nsew signal input
rlabel metal4 s 218838 0 218898 3708 6 um_ow[294]
port 600 nsew signal input
rlabel metal4 s 218102 0 218162 1396 6 um_ow[295]
port 601 nsew signal input
rlabel metal4 s 217366 0 217426 3164 6 um_ow[296]
port 602 nsew signal input
rlabel metal4 s 216630 0 216690 2892 6 um_ow[297]
port 603 nsew signal input
rlabel metal4 s 215894 0 215954 716 6 um_ow[298]
port 604 nsew signal input
rlabel metal4 s 215158 0 215218 3980 6 um_ow[299]
port 605 nsew signal input
rlabel metal4 s 14782 10164 14842 10880 6 um_ow[29]
port 606 nsew signal input
rlabel metal4 s 16990 0 17050 716 6 um_ow[2]
port 607 nsew signal input
rlabel metal4 s 214422 0 214482 308 6 um_ow[300]
port 608 nsew signal input
rlabel metal4 s 213686 0 213746 444 6 um_ow[301]
port 609 nsew signal input
rlabel metal4 s 212950 0 213010 308 6 um_ow[302]
port 610 nsew signal input
rlabel metal4 s 212214 0 212274 1804 6 um_ow[303]
port 611 nsew signal input
rlabel metal4 s 211478 0 211538 3028 6 um_ow[304]
port 612 nsew signal input
rlabel metal4 s 210742 0 210802 2756 6 um_ow[305]
port 613 nsew signal input
rlabel metal4 s 210006 0 210066 1396 6 um_ow[306]
port 614 nsew signal input
rlabel metal4 s 209270 0 209330 444 6 um_ow[307]
port 615 nsew signal input
rlabel metal4 s 208534 0 208594 852 6 um_ow[308]
port 616 nsew signal input
rlabel metal4 s 207798 0 207858 308 6 um_ow[309]
port 617 nsew signal input
rlabel metal4 s 14046 10164 14106 10880 6 um_ow[30]
port 618 nsew signal input
rlabel metal4 s 207062 0 207122 852 6 um_ow[310]
port 619 nsew signal input
rlabel metal4 s 206326 0 206386 852 6 um_ow[311]
port 620 nsew signal input
rlabel metal4 s 223254 10164 223314 10880 6 um_ow[312]
port 621 nsew signal input
rlabel metal4 s 222518 10164 222578 10880 6 um_ow[313]
port 622 nsew signal input
rlabel metal4 s 221782 9892 221842 10880 6 um_ow[314]
port 623 nsew signal input
rlabel metal4 s 221046 10436 221106 10880 6 um_ow[315]
port 624 nsew signal input
rlabel metal4 s 220310 10300 220370 10880 6 um_ow[316]
port 625 nsew signal input
rlabel metal4 s 219574 10164 219634 10880 6 um_ow[317]
port 626 nsew signal input
rlabel metal4 s 218838 10164 218898 10880 6 um_ow[318]
port 627 nsew signal input
rlabel metal4 s 218102 10572 218162 10880 6 um_ow[319]
port 628 nsew signal input
rlabel metal4 s 13310 9892 13370 10880 6 um_ow[31]
port 629 nsew signal input
rlabel metal4 s 217366 10164 217426 10880 6 um_ow[320]
port 630 nsew signal input
rlabel metal4 s 216630 9892 216690 10880 6 um_ow[321]
port 631 nsew signal input
rlabel metal4 s 215894 10164 215954 10880 6 um_ow[322]
port 632 nsew signal input
rlabel metal4 s 215158 9620 215218 10880 6 um_ow[323]
port 633 nsew signal input
rlabel metal4 s 214422 10164 214482 10880 6 um_ow[324]
port 634 nsew signal input
rlabel metal4 s 213686 10164 213746 10880 6 um_ow[325]
port 635 nsew signal input
rlabel metal4 s 212950 10572 213010 10880 6 um_ow[326]
port 636 nsew signal input
rlabel metal4 s 212214 10164 212274 10880 6 um_ow[327]
port 637 nsew signal input
rlabel metal4 s 211478 9892 211538 10880 6 um_ow[328]
port 638 nsew signal input
rlabel metal4 s 210742 10164 210802 10880 6 um_ow[329]
port 639 nsew signal input
rlabel metal4 s 12574 10164 12634 10880 6 um_ow[32]
port 640 nsew signal input
rlabel metal4 s 210006 10436 210066 10880 6 um_ow[330]
port 641 nsew signal input
rlabel metal4 s 209270 10164 209330 10880 6 um_ow[331]
port 642 nsew signal input
rlabel metal4 s 208534 10164 208594 10880 6 um_ow[332]
port 643 nsew signal input
rlabel metal4 s 207798 10572 207858 10880 6 um_ow[333]
port 644 nsew signal input
rlabel metal4 s 207062 10164 207122 10880 6 um_ow[334]
port 645 nsew signal input
rlabel metal4 s 206326 10164 206386 10880 6 um_ow[335]
port 646 nsew signal input
rlabel metal4 s 257386 0 257446 370 6 um_ow[336]
port 647 nsew signal input
rlabel metal4 s 256650 0 256710 370 6 um_ow[337]
port 648 nsew signal input
rlabel metal4 s 255914 0 255974 642 6 um_ow[338]
port 649 nsew signal input
rlabel metal4 s 255178 0 255238 580 6 um_ow[339]
port 650 nsew signal input
rlabel metal4 s 11838 10164 11898 10880 6 um_ow[33]
port 651 nsew signal input
rlabel metal4 s 254442 0 254502 580 6 um_ow[340]
port 652 nsew signal input
rlabel metal4 s 253706 0 253766 308 6 um_ow[341]
port 653 nsew signal input
rlabel metal4 s 252970 0 253030 444 6 um_ow[342]
port 654 nsew signal input
rlabel metal4 s 252234 0 252294 370 6 um_ow[343]
port 655 nsew signal input
rlabel metal4 s 251498 0 251558 370 6 um_ow[344]
port 656 nsew signal input
rlabel metal4 s 250762 0 250822 642 6 um_ow[345]
port 657 nsew signal input
rlabel metal4 s 250026 0 250086 580 6 um_ow[346]
port 658 nsew signal input
rlabel metal4 s 249290 0 249350 370 6 um_ow[347]
port 659 nsew signal input
rlabel metal4 s 248554 0 248614 370 6 um_ow[348]
port 660 nsew signal input
rlabel metal4 s 247818 0 247878 580 6 um_ow[349]
port 661 nsew signal input
rlabel metal4 s 11102 10164 11162 10880 6 um_ow[34]
port 662 nsew signal input
rlabel metal4 s 247082 0 247142 580 6 um_ow[350]
port 663 nsew signal input
rlabel metal4 s 246346 0 246406 642 6 um_ow[351]
port 664 nsew signal input
rlabel metal4 s 245610 0 245670 370 6 um_ow[352]
port 665 nsew signal input
rlabel metal4 s 244874 0 244934 580 6 um_ow[353]
port 666 nsew signal input
rlabel metal4 s 244138 0 244198 580 6 um_ow[354]
port 667 nsew signal input
rlabel metal4 s 243402 0 243462 580 6 um_ow[355]
port 668 nsew signal input
rlabel metal4 s 242666 0 242726 370 6 um_ow[356]
port 669 nsew signal input
rlabel metal4 s 241930 0 241990 580 6 um_ow[357]
port 670 nsew signal input
rlabel metal4 s 241194 0 241254 580 6 um_ow[358]
port 671 nsew signal input
rlabel metal4 s 240458 0 240518 580 6 um_ow[359]
port 672 nsew signal input
rlabel metal4 s 10366 10164 10426 10880 6 um_ow[35]
port 673 nsew signal input
rlabel metal4 s 257386 10300 257446 10880 6 um_ow[360]
port 674 nsew signal input
rlabel metal4 s 256650 10300 256710 10880 6 um_ow[361]
port 675 nsew signal input
rlabel metal4 s 255914 10300 255974 10880 6 um_ow[362]
port 676 nsew signal input
rlabel metal4 s 255178 10300 255238 10880 6 um_ow[363]
port 677 nsew signal input
rlabel metal4 s 254442 10300 254502 10880 6 um_ow[364]
port 678 nsew signal input
rlabel metal4 s 253706 10300 253766 10880 6 um_ow[365]
port 679 nsew signal input
rlabel metal4 s 252970 10436 253030 10880 6 um_ow[366]
port 680 nsew signal input
rlabel metal4 s 252234 10300 252294 10880 6 um_ow[367]
port 681 nsew signal input
rlabel metal4 s 251498 10300 251558 10880 6 um_ow[368]
port 682 nsew signal input
rlabel metal4 s 250762 10300 250822 10880 6 um_ow[369]
port 683 nsew signal input
rlabel metal4 s 9630 10164 9690 10880 6 um_ow[36]
port 684 nsew signal input
rlabel metal4 s 250026 10300 250086 10880 6 um_ow[370]
port 685 nsew signal input
rlabel metal4 s 249290 10300 249350 10880 6 um_ow[371]
port 686 nsew signal input
rlabel metal4 s 248554 10300 248614 10880 6 um_ow[372]
port 687 nsew signal input
rlabel metal4 s 247818 10300 247878 10880 6 um_ow[373]
port 688 nsew signal input
rlabel metal4 s 247082 10300 247142 10880 6 um_ow[374]
port 689 nsew signal input
rlabel metal4 s 246346 10300 246406 10880 6 um_ow[375]
port 690 nsew signal input
rlabel metal4 s 245610 10436 245670 10880 6 um_ow[376]
port 691 nsew signal input
rlabel metal4 s 244874 10300 244934 10880 6 um_ow[377]
port 692 nsew signal input
rlabel metal4 s 244138 10300 244198 10880 6 um_ow[378]
port 693 nsew signal input
rlabel metal4 s 243402 10300 243462 10880 6 um_ow[379]
port 694 nsew signal input
rlabel metal4 s 8894 10164 8954 10880 6 um_ow[37]
port 695 nsew signal input
rlabel metal4 s 242666 10300 242726 10880 6 um_ow[380]
port 696 nsew signal input
rlabel metal4 s 241930 10300 241990 10880 6 um_ow[381]
port 697 nsew signal input
rlabel metal4 s 241194 10300 241254 10880 6 um_ow[382]
port 698 nsew signal input
rlabel metal4 s 240458 10300 240518 10880 6 um_ow[383]
port 699 nsew signal input
rlabel metal4 s 8158 9892 8218 10880 6 um_ow[38]
port 700 nsew signal input
rlabel metal4 s 7422 10164 7482 10880 6 um_ow[39]
port 701 nsew signal input
rlabel metal4 s 16254 0 16314 716 6 um_ow[3]
port 702 nsew signal input
rlabel metal4 s 6686 10164 6746 10880 6 um_ow[40]
port 703 nsew signal input
rlabel metal4 s 5950 10164 6010 10880 6 um_ow[41]
port 704 nsew signal input
rlabel metal4 s 5214 10164 5274 10880 6 um_ow[42]
port 705 nsew signal input
rlabel metal4 s 4478 10164 4538 10880 6 um_ow[43]
port 706 nsew signal input
rlabel metal4 s 3742 10164 3802 10880 6 um_ow[44]
port 707 nsew signal input
rlabel metal4 s 3006 9892 3066 10880 6 um_ow[45]
port 708 nsew signal input
rlabel metal4 s 2270 10164 2330 10880 6 um_ow[46]
port 709 nsew signal input
rlabel metal4 s 1534 10164 1594 10880 6 um_ow[47]
port 710 nsew signal input
rlabel metal4 s 52594 0 52654 308 6 um_ow[48]
port 711 nsew signal input
rlabel metal4 s 51858 0 51918 580 6 um_ow[49]
port 712 nsew signal input
rlabel metal4 s 15518 0 15578 988 6 um_ow[4]
port 713 nsew signal input
rlabel metal4 s 51122 0 51182 580 6 um_ow[50]
port 714 nsew signal input
rlabel metal4 s 50386 0 50446 580 6 um_ow[51]
port 715 nsew signal input
rlabel metal4 s 49650 0 49710 580 6 um_ow[52]
port 716 nsew signal input
rlabel metal4 s 48914 0 48974 580 6 um_ow[53]
port 717 nsew signal input
rlabel metal4 s 48178 0 48238 580 6 um_ow[54]
port 718 nsew signal input
rlabel metal4 s 47442 0 47502 580 6 um_ow[55]
port 719 nsew signal input
rlabel metal4 s 46706 0 46766 580 6 um_ow[56]
port 720 nsew signal input
rlabel metal4 s 45970 0 46030 580 6 um_ow[57]
port 721 nsew signal input
rlabel metal4 s 45234 0 45294 580 6 um_ow[58]
port 722 nsew signal input
rlabel metal4 s 44498 0 44558 580 6 um_ow[59]
port 723 nsew signal input
rlabel metal4 s 14782 0 14842 1260 6 um_ow[5]
port 724 nsew signal input
rlabel metal4 s 43762 0 43822 580 6 um_ow[60]
port 725 nsew signal input
rlabel metal4 s 43026 0 43086 580 6 um_ow[61]
port 726 nsew signal input
rlabel metal4 s 42290 0 42350 580 6 um_ow[62]
port 727 nsew signal input
rlabel metal4 s 41554 0 41614 580 6 um_ow[63]
port 728 nsew signal input
rlabel metal4 s 40818 0 40878 580 6 um_ow[64]
port 729 nsew signal input
rlabel metal4 s 40082 0 40142 580 6 um_ow[65]
port 730 nsew signal input
rlabel metal4 s 39346 0 39406 308 6 um_ow[66]
port 731 nsew signal input
rlabel metal4 s 38610 0 38670 580 6 um_ow[67]
port 732 nsew signal input
rlabel metal4 s 37874 0 37934 580 6 um_ow[68]
port 733 nsew signal input
rlabel metal4 s 37138 0 37198 580 6 um_ow[69]
port 734 nsew signal input
rlabel metal4 s 14046 0 14106 988 6 um_ow[6]
port 735 nsew signal input
rlabel metal4 s 36402 0 36462 580 6 um_ow[70]
port 736 nsew signal input
rlabel metal4 s 35666 0 35726 580 6 um_ow[71]
port 737 nsew signal input
rlabel metal4 s 52594 10572 52654 10880 6 um_ow[72]
port 738 nsew signal input
rlabel metal4 s 51858 10300 51918 10880 6 um_ow[73]
port 739 nsew signal input
rlabel metal4 s 51122 10300 51182 10880 6 um_ow[74]
port 740 nsew signal input
rlabel metal4 s 50386 10300 50446 10880 6 um_ow[75]
port 741 nsew signal input
rlabel metal4 s 49650 10300 49710 10880 6 um_ow[76]
port 742 nsew signal input
rlabel metal4 s 48914 10300 48974 10880 6 um_ow[77]
port 743 nsew signal input
rlabel metal4 s 48178 10300 48238 10880 6 um_ow[78]
port 744 nsew signal input
rlabel metal4 s 47442 10300 47502 10880 6 um_ow[79]
port 745 nsew signal input
rlabel metal4 s 13310 0 13370 580 6 um_ow[7]
port 746 nsew signal input
rlabel metal4 s 46706 10300 46766 10880 6 um_ow[80]
port 747 nsew signal input
rlabel metal4 s 45970 10300 46030 10880 6 um_ow[81]
port 748 nsew signal input
rlabel metal4 s 45234 10300 45294 10880 6 um_ow[82]
port 749 nsew signal input
rlabel metal4 s 44498 10300 44558 10880 6 um_ow[83]
port 750 nsew signal input
rlabel metal4 s 43762 10300 43822 10880 6 um_ow[84]
port 751 nsew signal input
rlabel metal4 s 43026 10300 43086 10880 6 um_ow[85]
port 752 nsew signal input
rlabel metal4 s 42290 10300 42350 10880 6 um_ow[86]
port 753 nsew signal input
rlabel metal4 s 41554 10300 41614 10880 6 um_ow[87]
port 754 nsew signal input
rlabel metal4 s 40818 10300 40878 10880 6 um_ow[88]
port 755 nsew signal input
rlabel metal4 s 40082 10300 40142 10880 6 um_ow[89]
port 756 nsew signal input
rlabel metal4 s 12574 0 12634 988 6 um_ow[8]
port 757 nsew signal input
rlabel metal4 s 39346 10300 39406 10880 6 um_ow[90]
port 758 nsew signal input
rlabel metal4 s 38610 10300 38670 10880 6 um_ow[91]
port 759 nsew signal input
rlabel metal4 s 37874 10300 37934 10880 6 um_ow[92]
port 760 nsew signal input
rlabel metal4 s 37138 10300 37198 10880 6 um_ow[93]
port 761 nsew signal input
rlabel metal4 s 36402 10300 36462 10880 6 um_ow[94]
port 762 nsew signal input
rlabel metal4 s 35666 10300 35726 10880 6 um_ow[95]
port 763 nsew signal input
rlabel metal4 s 86726 0 86786 852 6 um_ow[96]
port 764 nsew signal input
rlabel metal4 s 85990 0 86050 988 6 um_ow[97]
port 765 nsew signal input
rlabel metal4 s 85254 0 85314 308 6 um_ow[98]
port 766 nsew signal input
rlabel metal4 s 84518 0 84578 988 6 um_ow[99]
port 767 nsew signal input
rlabel metal4 s 11838 0 11898 988 6 um_ow[9]
port 768 nsew signal input
rlabel metal4 s 34742 1040 35062 9840 6 vccd1
port 769 nsew power bidirectional
rlabel metal4 s 102339 1040 102659 9840 6 vccd1
port 769 nsew power bidirectional
rlabel metal4 s 169936 1040 170256 9840 6 vccd1
port 769 nsew power bidirectional
rlabel metal4 s 237533 1040 237853 9840 6 vccd1
port 769 nsew power bidirectional
rlabel metal4 s 68540 1040 68860 9840 6 vssd1
port 770 nsew ground bidirectional
rlabel metal4 s 136137 1040 136457 9840 6 vssd1
port 770 nsew ground bidirectional
rlabel metal4 s 203734 1040 204054 9840 6 vssd1
port 770 nsew ground bidirectional
rlabel metal4 s 271331 1040 271651 9840 6 vssd1
port 770 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 272600 11000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5064396
string GDS_FILE /home/uri/p/tinytapeout-03p5-gds/openlane/tt_mux/runs/23_06_01_20_50/results/signoff/tt_mux.magic.gds
string GDS_START 281990
<< end >>

