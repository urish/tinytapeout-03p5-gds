magic
tech sky130A
magscale 1 2
timestamp 1684932508
<< metal1 >>
rect 282730 190476 282736 190528
rect 282788 190516 282794 190528
rect 293862 190516 293868 190528
rect 282788 190488 293868 190516
rect 282788 190476 282794 190488
rect 293862 190476 293868 190488
rect 293920 190476 293926 190528
rect 296714 189252 296720 189304
rect 296772 189292 296778 189304
rect 300946 189292 300952 189304
rect 296772 189264 300952 189292
rect 296772 189252 296778 189264
rect 300946 189252 300952 189264
rect 301004 189252 301010 189304
rect 283282 187620 283288 187672
rect 283340 187660 283346 187672
rect 285674 187660 285680 187672
rect 283340 187632 285680 187660
rect 283340 187620 283346 187632
rect 285674 187620 285680 187632
rect 285732 187620 285738 187672
rect 298002 185648 298008 185700
rect 298060 185688 298066 185700
rect 300854 185688 300860 185700
rect 298060 185660 300860 185688
rect 298060 185648 298066 185660
rect 300854 185648 300860 185660
rect 300912 185648 300918 185700
rect 282546 184356 282552 184408
rect 282604 184396 282610 184408
rect 285582 184396 285588 184408
rect 282604 184368 285588 184396
rect 282604 184356 282610 184368
rect 285582 184356 285588 184368
rect 285640 184356 285646 184408
rect 292574 184152 292580 184204
rect 292632 184192 292638 184204
rect 300854 184192 300860 184204
rect 292632 184164 300860 184192
rect 292632 184152 292638 184164
rect 300854 184152 300860 184164
rect 300912 184152 300918 184204
rect 288342 182792 288348 182844
rect 288400 182832 288406 182844
rect 300854 182832 300860 182844
rect 288400 182804 300860 182832
rect 288400 182792 288406 182804
rect 300854 182792 300860 182804
rect 300912 182792 300918 182844
rect 282362 181432 282368 181484
rect 282420 181472 282426 181484
rect 300854 181472 300860 181484
rect 282420 181444 300860 181472
rect 282420 181432 282426 181444
rect 300854 181432 300860 181444
rect 300912 181432 300918 181484
rect 281810 179324 281816 179376
rect 281868 179364 281874 179376
rect 301774 179364 301780 179376
rect 281868 179336 301780 179364
rect 281868 179324 281874 179336
rect 301774 179324 301780 179336
rect 301832 179324 301838 179376
rect 249702 178508 249708 178560
rect 249760 178548 249766 178560
rect 251174 178548 251180 178560
rect 249760 178520 251180 178548
rect 249760 178508 249766 178520
rect 251174 178508 251180 178520
rect 251232 178508 251238 178560
rect 289906 177284 289912 177336
rect 289964 177324 289970 177336
rect 300854 177324 300860 177336
rect 289964 177296 300860 177324
rect 289964 177284 289970 177296
rect 300854 177284 300860 177296
rect 300912 177284 300918 177336
rect 249702 156612 249708 156664
rect 249760 156652 249766 156664
rect 261478 156652 261484 156664
rect 249760 156624 261484 156652
rect 249760 156612 249766 156624
rect 261478 156612 261484 156624
rect 261536 156612 261542 156664
rect 261478 148316 261484 148368
rect 261536 148356 261542 148368
rect 266998 148356 267004 148368
rect 261536 148328 267004 148356
rect 261536 148316 261542 148328
rect 266998 148316 267004 148328
rect 267056 148316 267062 148368
rect 266998 68960 267004 69012
rect 267056 69000 267062 69012
rect 282178 69000 282184 69012
rect 267056 68972 282184 69000
rect 267056 68960 267062 68972
rect 282178 68960 282184 68972
rect 282236 68960 282242 69012
<< via1 >>
rect 282736 190476 282788 190528
rect 293868 190476 293920 190528
rect 296720 189252 296772 189304
rect 300952 189252 301004 189304
rect 283288 187620 283340 187672
rect 285680 187620 285732 187672
rect 298008 185648 298060 185700
rect 300860 185648 300912 185700
rect 282552 184356 282604 184408
rect 285588 184356 285640 184408
rect 292580 184152 292632 184204
rect 300860 184152 300912 184204
rect 288348 182792 288400 182844
rect 300860 182792 300912 182844
rect 282368 181432 282420 181484
rect 300860 181432 300912 181484
rect 281816 179324 281868 179376
rect 301780 179324 301832 179376
rect 249708 178508 249760 178560
rect 251180 178508 251232 178560
rect 289912 177284 289964 177336
rect 300860 177284 300912 177336
rect 249708 156612 249760 156664
rect 261484 156612 261536 156664
rect 261484 148316 261536 148368
rect 267004 148316 267056 148368
rect 267004 68960 267056 69012
rect 282184 68960 282236 69012
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 701049 8156 703520
rect 6182 701040 6238 701049
rect 6182 700975 6238 700984
rect 8114 701040 8170 701049
rect 8114 700975 8170 700984
rect 6196 254289 6224 700975
rect 24320 700369 24348 703520
rect 72988 701049 73016 703520
rect 72974 701040 73030 701049
rect 72974 700975 73030 700984
rect 24306 700360 24362 700369
rect 24306 700295 24362 700304
rect 35162 700360 35218 700369
rect 35162 700295 35218 700304
rect 35176 671401 35204 700295
rect 35162 671392 35218 671401
rect 35162 671327 35218 671336
rect 42798 671392 42854 671401
rect 42798 671327 42854 671336
rect 6182 254280 6238 254289
rect 6182 254215 6238 254224
rect 2778 241088 2834 241097
rect 2778 241023 2834 241032
rect 2792 136785 2820 241023
rect 42812 191049 42840 671327
rect 89180 214577 89208 703520
rect 137848 701049 137876 703520
rect 137834 701040 137890 701049
rect 137834 700975 137890 700984
rect 154132 214713 154160 703520
rect 202800 701049 202828 703520
rect 202786 701040 202842 701049
rect 202786 700975 202842 700984
rect 154118 214704 154174 214713
rect 154118 214639 154174 214648
rect 89166 214568 89222 214577
rect 89166 214503 89222 214512
rect 218992 213217 219020 703520
rect 267660 701049 267688 703520
rect 267646 701040 267702 701049
rect 267646 700975 267702 700984
rect 283852 699825 283880 703520
rect 332520 701049 332548 703520
rect 332506 701040 332562 701049
rect 332506 700975 332562 700984
rect 348804 700369 348832 703520
rect 397472 701049 397500 703520
rect 397458 701040 397514 701049
rect 397458 700975 397514 700984
rect 295246 700360 295302 700369
rect 295246 700295 295302 700304
rect 348790 700360 348846 700369
rect 348790 700295 348846 700304
rect 283838 699816 283894 699825
rect 283838 699751 283894 699760
rect 218978 213208 219034 213217
rect 218978 213143 219034 213152
rect 290462 213208 290518 213217
rect 290462 213143 290518 213152
rect 282918 191720 282974 191729
rect 282918 191655 282974 191664
rect 9678 191040 9734 191049
rect 9678 190975 9734 190984
rect 42798 191040 42854 191049
rect 42798 190975 42854 190984
rect 9692 190454 9720 190975
rect 282736 190528 282788 190534
rect 282736 190470 282788 190476
rect 9600 190426 9720 190454
rect 9600 175273 9628 190426
rect 9770 189136 9826 189145
rect 9770 189071 9826 189080
rect 9784 180794 9812 189071
rect 282748 185745 282776 190470
rect 282826 186416 282882 186425
rect 282932 186402 282960 191655
rect 287058 190768 287114 190777
rect 287058 190703 287114 190712
rect 285678 189136 285734 189145
rect 285678 189071 285734 189080
rect 285692 187678 285720 189071
rect 287072 188329 287100 190703
rect 289726 189680 289782 189689
rect 289726 189615 289782 189624
rect 289740 188329 289768 189615
rect 287058 188320 287114 188329
rect 287058 188255 287114 188264
rect 289726 188320 289782 188329
rect 289726 188255 289782 188264
rect 283288 187672 283340 187678
rect 283286 187640 283288 187649
rect 285680 187672 285732 187678
rect 283340 187640 283342 187649
rect 285680 187614 285732 187620
rect 283286 187575 283342 187584
rect 286966 187368 287022 187377
rect 286966 187303 287022 187312
rect 282882 186374 282960 186402
rect 282826 186351 282882 186360
rect 284022 186144 284078 186153
rect 284022 186079 284078 186088
rect 282734 185736 282790 185745
rect 282734 185671 282790 185680
rect 284036 185065 284064 186079
rect 284022 185056 284078 185065
rect 284022 184991 284078 185000
rect 282552 184408 282604 184414
rect 282550 184376 282552 184385
rect 285588 184408 285640 184414
rect 282604 184376 282606 184385
rect 282550 184311 282606 184320
rect 282918 184376 282974 184385
rect 282918 184311 282974 184320
rect 285586 184376 285588 184385
rect 285640 184376 285642 184385
rect 285586 184311 285642 184320
rect 282932 182730 282960 184311
rect 285586 183696 285642 183705
rect 285586 183631 285642 183640
rect 282748 182702 282960 182730
rect 282368 181484 282420 181490
rect 282368 181426 282420 181432
rect 281814 180976 281870 180985
rect 281814 180911 281870 180920
rect 9784 180766 9904 180794
rect 9586 175264 9642 175273
rect 9586 175199 9642 175208
rect 2778 136776 2834 136785
rect 2778 136711 2834 136720
rect 2792 45529 2820 136711
rect 9876 68513 9904 180766
rect 281828 179382 281856 180911
rect 282380 180849 282408 181426
rect 282748 181121 282776 182702
rect 282918 182608 282974 182617
rect 282918 182543 282974 182552
rect 282734 181112 282790 181121
rect 282734 181047 282790 181056
rect 282366 180840 282422 180849
rect 282366 180775 282422 180784
rect 281816 179376 281868 179382
rect 251178 179344 251234 179353
rect 251178 179279 251234 179288
rect 281814 179344 281816 179353
rect 281868 179344 281870 179353
rect 281814 179279 281870 179288
rect 251192 178566 251220 179279
rect 282826 178800 282882 178809
rect 282826 178735 282882 178744
rect 249708 178560 249760 178566
rect 249708 178502 249760 178508
rect 251180 178560 251232 178566
rect 251180 178502 251232 178508
rect 11702 157448 11758 157457
rect 11702 157383 11758 157392
rect 11716 148345 11744 157383
rect 249720 156670 249748 178502
rect 280894 176080 280950 176089
rect 280894 176015 280950 176024
rect 280908 161474 280936 176015
rect 280816 161446 280936 161474
rect 249708 156664 249760 156670
rect 249708 156606 249760 156612
rect 261484 156664 261536 156670
rect 261484 156606 261536 156612
rect 261496 148374 261524 156606
rect 261484 148368 261536 148374
rect 11702 148336 11758 148345
rect 267004 148368 267056 148374
rect 261484 148310 261536 148316
rect 262862 148336 262918 148345
rect 11702 148271 11758 148280
rect 267004 148310 267056 148316
rect 262862 148271 262918 148280
rect 262876 70825 262904 148271
rect 262862 70816 262918 70825
rect 262862 70751 262918 70760
rect 265070 70816 265126 70825
rect 265070 70751 265126 70760
rect 9862 68504 9918 68513
rect 9862 68439 9918 68448
rect 265084 67153 265112 70751
rect 267016 69018 267044 148310
rect 267004 69012 267056 69018
rect 267004 68954 267056 68960
rect 280816 67561 280844 161446
rect 282840 69601 282868 178735
rect 282932 177449 282960 182543
rect 283010 182200 283066 182209
rect 283010 182135 283066 182144
rect 283024 180169 283052 182135
rect 283562 181248 283618 181257
rect 283562 181183 283618 181192
rect 283010 180160 283066 180169
rect 283010 180095 283066 180104
rect 282918 177440 282974 177449
rect 282918 177375 282974 177384
rect 282826 69592 282882 69601
rect 282826 69527 282882 69536
rect 282184 69012 282236 69018
rect 282184 68954 282236 68960
rect 282196 67697 282224 68954
rect 282182 67688 282238 67697
rect 282182 67623 282238 67632
rect 283576 67561 283604 181183
rect 285600 156641 285628 183631
rect 286980 177313 287008 187303
rect 288438 183560 288494 183569
rect 288438 183495 288494 183504
rect 288346 183152 288402 183161
rect 288346 183087 288402 183096
rect 288360 182850 288388 183087
rect 288348 182844 288400 182850
rect 288348 182786 288400 182792
rect 287058 182608 287114 182617
rect 287058 182543 287114 182552
rect 287072 178809 287100 182543
rect 287058 178800 287114 178809
rect 287058 178735 287114 178744
rect 286966 177304 287022 177313
rect 286966 177239 287022 177248
rect 288452 176089 288480 183495
rect 289910 179480 289966 179489
rect 289910 179415 289966 179424
rect 289924 177342 289952 179415
rect 289912 177336 289964 177342
rect 289912 177278 289964 177284
rect 288438 176080 288494 176089
rect 288438 176015 288494 176024
rect 285586 156632 285642 156641
rect 285586 156567 285642 156576
rect 280802 67552 280858 67561
rect 280802 67487 280858 67496
rect 283562 67552 283618 67561
rect 283562 67487 283618 67496
rect 265070 67144 265126 67153
rect 265070 67079 265126 67088
rect 290476 66881 290504 213143
rect 293868 190528 293920 190534
rect 293868 190470 293920 190476
rect 292946 185736 293002 185745
rect 292946 185671 293002 185680
rect 292960 185473 292988 185671
rect 293880 185609 293908 190470
rect 293866 185600 293922 185609
rect 293866 185535 293922 185544
rect 292946 185464 293002 185473
rect 292946 185399 293002 185408
rect 292486 184920 292542 184929
rect 292486 184855 292542 184864
rect 292026 180160 292082 180169
rect 292026 180095 292082 180104
rect 292040 178945 292068 180095
rect 292026 178936 292082 178945
rect 292026 178871 292082 178880
rect 292500 174593 292528 184855
rect 293222 184784 293278 184793
rect 293222 184719 293278 184728
rect 292578 184376 292634 184385
rect 292578 184311 292634 184320
rect 292592 184210 292620 184311
rect 292580 184204 292632 184210
rect 292580 184146 292632 184152
rect 292592 183705 292620 184146
rect 292578 183696 292634 183705
rect 292578 183631 292634 183640
rect 292486 174584 292542 174593
rect 292486 174519 292542 174528
rect 293236 68921 293264 184719
rect 295260 180305 295288 700295
rect 295982 214704 296038 214713
rect 295982 214639 296038 214648
rect 295246 180296 295302 180305
rect 295246 180231 295302 180240
rect 295996 178673 296024 214639
rect 413664 213353 413692 703520
rect 462332 701049 462360 703520
rect 462318 701040 462374 701049
rect 462318 700975 462374 700984
rect 301502 213344 301558 213353
rect 301502 213279 301558 213288
rect 413650 213344 413706 213353
rect 413650 213279 413706 213288
rect 298834 213208 298890 213217
rect 298834 213143 298890 213152
rect 298848 210361 298876 213143
rect 298834 210352 298890 210361
rect 298834 210287 298890 210296
rect 301516 192545 301544 213279
rect 478524 213217 478552 703520
rect 527192 701049 527220 703520
rect 543476 701049 543504 703520
rect 527178 701040 527234 701049
rect 527178 700975 527234 700984
rect 543462 701040 543518 701049
rect 543462 700975 543518 700984
rect 543476 700369 543504 700975
rect 559668 700505 559696 703520
rect 559654 700496 559710 700505
rect 559654 700431 559710 700440
rect 582378 700496 582434 700505
rect 582378 700431 582434 700440
rect 543462 700360 543518 700369
rect 543462 700295 543518 700304
rect 580446 700360 580502 700369
rect 580446 700295 580502 700304
rect 580460 697241 580488 700295
rect 580446 697232 580502 697241
rect 580446 697167 580502 697176
rect 580906 697232 580962 697241
rect 580906 697167 580962 697176
rect 580920 683913 580948 697167
rect 580906 683904 580962 683913
rect 580906 683839 580962 683848
rect 580920 644065 580948 683839
rect 580906 644056 580962 644065
rect 580906 643991 580962 644000
rect 580920 630873 580948 643991
rect 580906 630864 580962 630873
rect 580906 630799 580962 630808
rect 580920 591025 580948 630799
rect 580906 591016 580962 591025
rect 580906 590951 580962 590960
rect 580920 577697 580948 590951
rect 580906 577688 580962 577697
rect 580906 577623 580962 577632
rect 580920 537849 580948 577623
rect 580906 537840 580962 537849
rect 580906 537775 580962 537784
rect 580920 524521 580948 537775
rect 580906 524512 580962 524521
rect 580906 524447 580962 524456
rect 580920 484673 580948 524447
rect 580906 484664 580962 484673
rect 580906 484599 580962 484608
rect 580920 471481 580948 484599
rect 580906 471472 580962 471481
rect 580906 471407 580962 471416
rect 580920 431633 580948 471407
rect 580906 431624 580962 431633
rect 580906 431559 580962 431568
rect 580920 418305 580948 431559
rect 580906 418296 580962 418305
rect 580906 418231 580962 418240
rect 580920 378457 580948 418231
rect 580906 378448 580962 378457
rect 580906 378383 580962 378392
rect 580920 365129 580948 378383
rect 580906 365120 580962 365129
rect 580906 365055 580962 365064
rect 580920 325281 580948 365055
rect 580906 325272 580962 325281
rect 580906 325207 580962 325216
rect 580920 312089 580948 325207
rect 580906 312080 580962 312089
rect 580906 312015 580962 312024
rect 580920 272241 580948 312015
rect 580906 272232 580962 272241
rect 580906 272167 580962 272176
rect 580920 258913 580948 272167
rect 580906 258904 580962 258913
rect 580906 258839 580962 258848
rect 478510 213208 478566 213217
rect 478510 213143 478566 213152
rect 301502 192536 301558 192545
rect 301502 192471 301558 192480
rect 296718 192128 296774 192137
rect 296718 192063 296774 192072
rect 296732 189310 296760 192063
rect 300306 190904 300362 190913
rect 300306 190839 300362 190848
rect 296720 189304 296772 189310
rect 296626 189272 296682 189281
rect 296720 189246 296772 189252
rect 296626 189207 296682 189216
rect 296640 186017 296668 189207
rect 299754 187096 299810 187105
rect 299754 187031 299810 187040
rect 296626 186008 296682 186017
rect 296626 185943 296682 185952
rect 296640 180849 296668 185943
rect 299768 185745 299796 187031
rect 298006 185736 298062 185745
rect 298006 185671 298008 185680
rect 298060 185671 298062 185680
rect 299754 185736 299810 185745
rect 299754 185671 299810 185680
rect 298008 185642 298060 185648
rect 300320 183705 300348 190839
rect 300766 190768 300822 190777
rect 300766 190703 300822 190712
rect 300780 189145 300808 190703
rect 300952 189304 301004 189310
rect 300952 189246 301004 189252
rect 300766 189136 300822 189145
rect 300766 189071 300822 189080
rect 300858 185736 300914 185745
rect 300858 185671 300860 185680
rect 300912 185671 300914 185680
rect 300860 185642 300912 185648
rect 300858 184376 300914 184385
rect 300858 184311 300914 184320
rect 300872 184210 300900 184311
rect 300860 184204 300912 184210
rect 300860 184146 300912 184152
rect 300306 183696 300362 183705
rect 300306 183631 300362 183640
rect 300858 183152 300914 183161
rect 300858 183087 300914 183096
rect 300872 182850 300900 183087
rect 300860 182844 300912 182850
rect 300860 182786 300912 182792
rect 300860 181484 300912 181490
rect 300860 181426 300912 181432
rect 300872 180849 300900 181426
rect 300964 181121 300992 189246
rect 302330 189136 302386 189145
rect 302330 189071 302386 189080
rect 302344 188465 302372 189071
rect 302330 188456 302386 188465
rect 302330 188391 302386 188400
rect 302238 182200 302294 182209
rect 302238 182135 302294 182144
rect 300950 181112 301006 181121
rect 300950 181047 301006 181056
rect 301778 180976 301834 180985
rect 301778 180911 301834 180920
rect 296626 180840 296682 180849
rect 296626 180775 296682 180784
rect 300858 180840 300914 180849
rect 300858 180775 300914 180784
rect 301792 179382 301820 180911
rect 301780 179376 301832 179382
rect 301780 179318 301832 179324
rect 302252 178945 302280 182135
rect 302330 180296 302386 180305
rect 302330 180231 302386 180240
rect 302238 178936 302294 178945
rect 302238 178871 302294 178880
rect 295982 178664 296038 178673
rect 295982 178599 296038 178608
rect 296166 178120 296222 178129
rect 296166 178055 296222 178064
rect 296180 158001 296208 178055
rect 300860 177336 300912 177342
rect 300860 177278 300912 177284
rect 296166 157992 296222 158001
rect 296166 157927 296222 157936
rect 300872 68921 300900 177278
rect 302344 171134 302372 180231
rect 335358 178664 335414 178673
rect 335358 178599 335414 178608
rect 302344 171106 302648 171134
rect 302620 156913 302648 171106
rect 306378 157992 306434 158001
rect 306378 157927 306434 157936
rect 302606 156904 302662 156913
rect 302606 156839 302662 156848
rect 304998 156496 305054 156505
rect 304998 156431 305054 156440
rect 304906 72448 304962 72457
rect 304906 72383 304962 72392
rect 293222 68912 293278 68921
rect 293222 68847 293278 68856
rect 300858 68912 300914 68921
rect 300858 68847 300914 68856
rect 304920 67561 304948 72383
rect 305012 68921 305040 156431
rect 306392 72457 306420 157927
rect 306378 72448 306434 72457
rect 306378 72383 306434 72392
rect 304998 68912 305054 68921
rect 304998 68847 305054 68856
rect 335372 68513 335400 178599
rect 573638 174584 573694 174593
rect 573638 174519 573694 174528
rect 573652 161474 573680 174519
rect 573376 161446 573680 161474
rect 335358 68504 335414 68513
rect 335358 68439 335414 68448
rect 304906 67552 304962 67561
rect 304906 67487 304962 67496
rect 290462 66872 290518 66881
rect 290462 66807 290518 66816
rect 2778 45520 2834 45529
rect 2778 45455 2834 45464
rect 2792 44305 2820 45455
rect 2778 44296 2834 44305
rect 2778 44231 2834 44240
rect 3422 44296 3478 44305
rect 3422 44231 3478 44240
rect 3436 24177 3464 44231
rect 3422 24168 3478 24177
rect 3422 24103 3478 24112
rect 273258 24168 273314 24177
rect 273258 24103 273314 24112
rect 273272 20233 273300 24103
rect 573376 20505 573404 161446
rect 580920 152697 580948 258839
rect 580906 152688 580962 152697
rect 580906 152623 580962 152632
rect 580920 139369 580948 152623
rect 580906 139360 580962 139369
rect 580906 139295 580962 139304
rect 580920 112849 580948 139295
rect 580906 112840 580962 112849
rect 580906 112775 580962 112784
rect 580920 99521 580948 112775
rect 580906 99512 580962 99521
rect 580906 99447 580962 99456
rect 580920 73001 580948 99447
rect 580906 72992 580962 73001
rect 580906 72927 580962 72936
rect 580920 59673 580948 72927
rect 582392 68241 582420 700431
rect 582378 68232 582434 68241
rect 582378 68167 582434 68176
rect 580906 59664 580962 59673
rect 580906 59599 580962 59608
rect 580920 33153 580948 59599
rect 580906 33144 580962 33153
rect 580906 33079 580962 33088
rect 573362 20496 573418 20505
rect 573362 20431 573418 20440
rect 273258 20224 273314 20233
rect 273258 20159 273314 20168
rect 278686 20224 278742 20233
rect 278686 20159 278742 20168
rect 2778 19544 2834 19553
rect 2778 19479 2834 19488
rect 277306 19544 277362 19553
rect 277306 19479 277362 19488
rect 2792 6497 2820 19479
rect 277320 19009 277348 19479
rect 278700 19417 278728 20159
rect 580920 19825 580948 33079
rect 580906 19816 580962 19825
rect 580906 19751 580962 19760
rect 278686 19408 278742 19417
rect 278686 19343 278742 19352
rect 277306 19000 277362 19009
rect 277306 18935 277362 18944
rect 2778 6488 2834 6497
rect 2778 6423 2834 6432
rect 579802 3496 579858 3505
rect 579802 3431 579858 3440
rect 579816 480 579844 3431
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 6182 700984 6238 701040
rect 8114 700984 8170 701040
rect 72974 700984 73030 701040
rect 24306 700304 24362 700360
rect 35162 700304 35218 700360
rect 35162 671336 35218 671392
rect 42798 671336 42854 671392
rect 6182 254224 6238 254280
rect 2778 241032 2834 241088
rect 137834 700984 137890 701040
rect 202786 700984 202842 701040
rect 154118 214648 154174 214704
rect 89166 214512 89222 214568
rect 267646 700984 267702 701040
rect 332506 700984 332562 701040
rect 397458 700984 397514 701040
rect 295246 700304 295302 700360
rect 348790 700304 348846 700360
rect 283838 699760 283894 699816
rect 218978 213152 219034 213208
rect 290462 213152 290518 213208
rect 282918 191664 282974 191720
rect 9678 190984 9734 191040
rect 42798 190984 42854 191040
rect 9770 189080 9826 189136
rect 282826 186360 282882 186416
rect 287058 190712 287114 190768
rect 285678 189080 285734 189136
rect 289726 189624 289782 189680
rect 287058 188264 287114 188320
rect 289726 188264 289782 188320
rect 283286 187620 283288 187640
rect 283288 187620 283340 187640
rect 283340 187620 283342 187640
rect 283286 187584 283342 187620
rect 286966 187312 287022 187368
rect 284022 186088 284078 186144
rect 282734 185680 282790 185736
rect 284022 185000 284078 185056
rect 282550 184356 282552 184376
rect 282552 184356 282604 184376
rect 282604 184356 282606 184376
rect 282550 184320 282606 184356
rect 282918 184320 282974 184376
rect 285586 184356 285588 184376
rect 285588 184356 285640 184376
rect 285640 184356 285642 184376
rect 285586 184320 285642 184356
rect 285586 183640 285642 183696
rect 281814 180920 281870 180976
rect 9586 175208 9642 175264
rect 2778 136720 2834 136776
rect 282918 182552 282974 182608
rect 282734 181056 282790 181112
rect 282366 180784 282422 180840
rect 251178 179288 251234 179344
rect 281814 179324 281816 179344
rect 281816 179324 281868 179344
rect 281868 179324 281870 179344
rect 281814 179288 281870 179324
rect 282826 178744 282882 178800
rect 11702 157392 11758 157448
rect 280894 176024 280950 176080
rect 11702 148280 11758 148336
rect 262862 148280 262918 148336
rect 262862 70760 262918 70816
rect 265070 70760 265126 70816
rect 9862 68448 9918 68504
rect 283010 182144 283066 182200
rect 283562 181192 283618 181248
rect 283010 180104 283066 180160
rect 282918 177384 282974 177440
rect 282826 69536 282882 69592
rect 282182 67632 282238 67688
rect 288438 183504 288494 183560
rect 288346 183096 288402 183152
rect 287058 182552 287114 182608
rect 287058 178744 287114 178800
rect 286966 177248 287022 177304
rect 289910 179424 289966 179480
rect 288438 176024 288494 176080
rect 285586 156576 285642 156632
rect 280802 67496 280858 67552
rect 283562 67496 283618 67552
rect 265070 67088 265126 67144
rect 292946 185680 293002 185736
rect 293866 185544 293922 185600
rect 292946 185408 293002 185464
rect 292486 184864 292542 184920
rect 292026 180104 292082 180160
rect 292026 178880 292082 178936
rect 293222 184728 293278 184784
rect 292578 184320 292634 184376
rect 292578 183640 292634 183696
rect 292486 174528 292542 174584
rect 295982 214648 296038 214704
rect 295246 180240 295302 180296
rect 462318 700984 462374 701040
rect 301502 213288 301558 213344
rect 413650 213288 413706 213344
rect 298834 213152 298890 213208
rect 298834 210296 298890 210352
rect 527178 700984 527234 701040
rect 543462 700984 543518 701040
rect 559654 700440 559710 700496
rect 582378 700440 582434 700496
rect 543462 700304 543518 700360
rect 580446 700304 580502 700360
rect 580446 697176 580502 697232
rect 580906 697176 580962 697232
rect 580906 683848 580962 683904
rect 580906 644000 580962 644056
rect 580906 630808 580962 630864
rect 580906 590960 580962 591016
rect 580906 577632 580962 577688
rect 580906 537784 580962 537840
rect 580906 524456 580962 524512
rect 580906 484608 580962 484664
rect 580906 471416 580962 471472
rect 580906 431568 580962 431624
rect 580906 418240 580962 418296
rect 580906 378392 580962 378448
rect 580906 365064 580962 365120
rect 580906 325216 580962 325272
rect 580906 312024 580962 312080
rect 580906 272176 580962 272232
rect 580906 258848 580962 258904
rect 478510 213152 478566 213208
rect 301502 192480 301558 192536
rect 296718 192072 296774 192128
rect 300306 190848 300362 190904
rect 296626 189216 296682 189272
rect 299754 187040 299810 187096
rect 296626 185952 296682 186008
rect 298006 185700 298062 185736
rect 298006 185680 298008 185700
rect 298008 185680 298060 185700
rect 298060 185680 298062 185700
rect 299754 185680 299810 185736
rect 300766 190712 300822 190768
rect 300766 189080 300822 189136
rect 300858 185700 300914 185736
rect 300858 185680 300860 185700
rect 300860 185680 300912 185700
rect 300912 185680 300914 185700
rect 300858 184320 300914 184376
rect 300306 183640 300362 183696
rect 300858 183096 300914 183152
rect 302330 189080 302386 189136
rect 302330 188400 302386 188456
rect 302238 182144 302294 182200
rect 300950 181056 301006 181112
rect 301778 180920 301834 180976
rect 296626 180784 296682 180840
rect 300858 180784 300914 180840
rect 302330 180240 302386 180296
rect 302238 178880 302294 178936
rect 295982 178608 296038 178664
rect 296166 178064 296222 178120
rect 296166 157936 296222 157992
rect 335358 178608 335414 178664
rect 306378 157936 306434 157992
rect 302606 156848 302662 156904
rect 304998 156440 305054 156496
rect 304906 72392 304962 72448
rect 293222 68856 293278 68912
rect 300858 68856 300914 68912
rect 306378 72392 306434 72448
rect 304998 68856 305054 68912
rect 573638 174528 573694 174584
rect 335358 68448 335414 68504
rect 304906 67496 304962 67552
rect 290462 66816 290518 66872
rect 2778 45464 2834 45520
rect 2778 44240 2834 44296
rect 3422 44240 3478 44296
rect 3422 24112 3478 24168
rect 273258 24112 273314 24168
rect 580906 152632 580962 152688
rect 580906 139304 580962 139360
rect 580906 112784 580962 112840
rect 580906 99456 580962 99512
rect 580906 72936 580962 72992
rect 582378 68176 582434 68232
rect 580906 59608 580962 59664
rect 580906 33088 580962 33144
rect 573362 20440 573418 20496
rect 273258 20168 273314 20224
rect 278686 20168 278742 20224
rect 2778 19488 2834 19544
rect 277306 19488 277362 19544
rect 580906 19760 580962 19816
rect 278686 19352 278742 19408
rect 277306 18944 277362 19000
rect 2778 6432 2834 6488
rect 579802 3440 579858 3496
<< metal3 >>
rect 6177 701042 6243 701045
rect 8109 701042 8175 701045
rect 72969 701042 73035 701045
rect 137829 701042 137895 701045
rect 202781 701042 202847 701045
rect 267641 701042 267707 701045
rect 332501 701042 332567 701045
rect 397453 701042 397519 701045
rect 462313 701042 462379 701045
rect 6177 701040 462379 701042
rect 6177 700984 6182 701040
rect 6238 700984 8114 701040
rect 8170 700984 72974 701040
rect 73030 700984 137834 701040
rect 137890 700984 202786 701040
rect 202842 700984 267646 701040
rect 267702 700984 332506 701040
rect 332562 700984 397458 701040
rect 397514 700984 462318 701040
rect 462374 700984 462379 701040
rect 6177 700982 462379 700984
rect 6177 700979 6243 700982
rect 8109 700979 8175 700982
rect 72969 700979 73035 700982
rect 137829 700979 137895 700982
rect 202781 700979 202847 700982
rect 267641 700979 267707 700982
rect 332501 700979 332567 700982
rect 397453 700979 397519 700982
rect 462313 700979 462379 700982
rect 527173 701042 527239 701045
rect 543457 701042 543523 701045
rect 527173 701040 543523 701042
rect 527173 700984 527178 701040
rect 527234 700984 543462 701040
rect 543518 700984 543523 701040
rect 527173 700982 543523 700984
rect 527173 700979 527239 700982
rect 543457 700979 543523 700982
rect 559649 700498 559715 700501
rect 582373 700498 582439 700501
rect 559649 700496 582439 700498
rect 559649 700440 559654 700496
rect 559710 700440 582378 700496
rect 582434 700440 582439 700496
rect 559649 700438 582439 700440
rect 559649 700435 559715 700438
rect 582373 700435 582439 700438
rect 24301 700362 24367 700365
rect 35157 700362 35223 700365
rect 24301 700360 35223 700362
rect 24301 700304 24306 700360
rect 24362 700304 35162 700360
rect 35218 700304 35223 700360
rect 24301 700302 35223 700304
rect 24301 700299 24367 700302
rect 35157 700299 35223 700302
rect 295241 700362 295307 700365
rect 348785 700362 348851 700365
rect 295241 700360 348851 700362
rect 295241 700304 295246 700360
rect 295302 700304 348790 700360
rect 348846 700304 348851 700360
rect 295241 700302 348851 700304
rect 295241 700299 295307 700302
rect 348785 700299 348851 700302
rect 543457 700362 543523 700365
rect 580441 700362 580507 700365
rect 543457 700360 580507 700362
rect 543457 700304 543462 700360
rect 543518 700304 580446 700360
rect 580502 700304 580507 700360
rect 543457 700302 580507 700304
rect 543457 700299 543523 700302
rect 580441 700299 580507 700302
rect 283833 699818 283899 699821
rect 284334 699818 284340 699820
rect 283833 699816 284340 699818
rect 283833 699760 283838 699816
rect 283894 699760 284340 699816
rect 283833 699758 284340 699760
rect 283833 699755 283899 699758
rect 284334 699756 284340 699758
rect 284404 699756 284410 699820
rect -960 697220 480 697460
rect 580441 697234 580507 697237
rect 580901 697234 580967 697237
rect 583520 697234 584960 697324
rect 580441 697232 584960 697234
rect 580441 697176 580446 697232
rect 580502 697176 580906 697232
rect 580962 697176 584960 697232
rect 580441 697174 584960 697176
rect 580441 697171 580507 697174
rect 580901 697171 580967 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 9806 684314 9812 684316
rect -960 684254 9812 684314
rect -960 684164 480 684254
rect 9806 684252 9812 684254
rect 9876 684252 9882 684316
rect 580901 683906 580967 683909
rect 583520 683906 584960 683996
rect 580901 683904 584960 683906
rect 580901 683848 580906 683904
rect 580962 683848 584960 683904
rect 580901 683846 584960 683848
rect 580901 683843 580967 683846
rect 583520 683756 584960 683846
rect 35157 671394 35223 671397
rect 42793 671394 42859 671397
rect 35157 671392 42859 671394
rect -960 671258 480 671348
rect 35157 671336 35162 671392
rect 35218 671336 42798 671392
rect 42854 671336 42859 671392
rect 35157 671334 42859 671336
rect 35157 671331 35223 671334
rect 42793 671331 42859 671334
rect 3366 671258 3372 671260
rect -960 671198 3372 671258
rect -960 671108 480 671198
rect 3366 671196 3372 671198
rect 3436 671196 3442 671260
rect 574686 670652 574692 670716
rect 574756 670714 574762 670716
rect 583520 670714 584960 670804
rect 574756 670654 584960 670714
rect 574756 670652 574762 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 291142 658202 291148 658204
rect -960 658142 291148 658202
rect -960 658052 480 658142
rect 291142 658140 291148 658142
rect 291212 658140 291218 658204
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580901 644058 580967 644061
rect 583520 644058 584960 644148
rect 580901 644056 584960 644058
rect 580901 644000 580906 644056
rect 580962 644000 584960 644056
rect 580901 643998 584960 644000
rect 580901 643995 580967 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 8886 632090 8892 632092
rect -960 632030 8892 632090
rect -960 631940 480 632030
rect 8886 632028 8892 632030
rect 8956 632028 8962 632092
rect 580901 630866 580967 630869
rect 583520 630866 584960 630956
rect 580901 630864 584960 630866
rect 580901 630808 580906 630864
rect 580962 630808 584960 630864
rect 580901 630806 584960 630808
rect 580901 630803 580967 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 4654 619170 4660 619172
rect -960 619110 4660 619170
rect -960 619020 480 619110
rect 4654 619108 4660 619110
rect 4724 619108 4730 619172
rect 575974 617476 575980 617540
rect 576044 617538 576050 617540
rect 583520 617538 584960 617628
rect 576044 617478 584960 617538
rect 576044 617476 576050 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 288382 606114 288388 606116
rect -960 606054 288388 606114
rect -960 605964 480 606054
rect 288382 606052 288388 606054
rect 288452 606052 288458 606116
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580901 591018 580967 591021
rect 583520 591018 584960 591108
rect 580901 591016 584960 591018
rect 580901 590960 580906 591016
rect 580962 590960 584960 591016
rect 580901 590958 584960 590960
rect 580901 590955 580967 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 7414 580002 7420 580004
rect -960 579942 7420 580002
rect -960 579852 480 579942
rect 7414 579940 7420 579942
rect 7484 579940 7490 580004
rect 580901 577690 580967 577693
rect 583520 577690 584960 577780
rect 580901 577688 584960 577690
rect 580901 577632 580906 577688
rect 580962 577632 584960 577688
rect 580901 577630 584960 577632
rect 580901 577627 580967 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 282126 566946 282132 566948
rect -960 566886 282132 566946
rect -960 566796 480 566886
rect 282126 566884 282132 566886
rect 282196 566884 282202 566948
rect 578734 564300 578740 564364
rect 578804 564362 578810 564364
rect 583520 564362 584960 564452
rect 578804 564302 584960 564362
rect 578804 564300 578810 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 17902 553890 17908 553892
rect -960 553830 17908 553890
rect -960 553740 480 553830
rect 17902 553828 17908 553830
rect 17972 553828 17978 553892
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580901 537842 580967 537845
rect 583520 537842 584960 537932
rect 580901 537840 584960 537842
rect 580901 537784 580906 537840
rect 580962 537784 584960 537840
rect 580901 537782 584960 537784
rect 580901 537779 580967 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2814 527914 2820 527916
rect -960 527854 2820 527914
rect -960 527764 480 527854
rect 2814 527852 2820 527854
rect 2884 527852 2890 527916
rect 580901 524514 580967 524517
rect 583520 524514 584960 524604
rect 580901 524512 584960 524514
rect 580901 524456 580906 524512
rect 580962 524456 584960 524512
rect 580901 524454 584960 524456
rect 580901 524451 580967 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 4838 514858 4844 514860
rect -960 514798 4844 514858
rect -960 514708 480 514798
rect 4838 514796 4844 514798
rect 4908 514796 4914 514860
rect 574870 511260 574876 511324
rect 574940 511322 574946 511324
rect 583520 511322 584960 511412
rect 574940 511262 584960 511322
rect 574940 511260 574946 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 12382 501802 12388 501804
rect -960 501742 12388 501802
rect -960 501652 480 501742
rect 12382 501740 12388 501742
rect 12452 501740 12458 501804
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580901 484666 580967 484669
rect 583520 484666 584960 484756
rect 580901 484664 584960 484666
rect 580901 484608 580906 484664
rect 580962 484608 584960 484664
rect 580901 484606 584960 484608
rect 580901 484603 580967 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 1894 475690 1900 475692
rect -960 475630 1900 475690
rect -960 475540 480 475630
rect 1894 475628 1900 475630
rect 1964 475628 1970 475692
rect 580901 471474 580967 471477
rect 583520 471474 584960 471564
rect 580901 471472 584960 471474
rect 580901 471416 580906 471472
rect 580962 471416 584960 471472
rect 580901 471414 584960 471416
rect 580901 471411 580967 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 13854 462634 13860 462636
rect -960 462574 13860 462634
rect -960 462484 480 462574
rect 13854 462572 13860 462574
rect 13924 462572 13930 462636
rect 578918 458084 578924 458148
rect 578988 458146 578994 458148
rect 583520 458146 584960 458236
rect 578988 458086 584960 458146
rect 578988 458084 578994 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 11094 449578 11100 449580
rect -960 449518 11100 449578
rect -960 449428 480 449518
rect 11094 449516 11100 449518
rect 11164 449516 11170 449580
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580901 431626 580967 431629
rect 583520 431626 584960 431716
rect 580901 431624 584960 431626
rect 580901 431568 580906 431624
rect 580962 431568 584960 431624
rect 580901 431566 584960 431568
rect 580901 431563 580967 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 9070 423602 9076 423604
rect -960 423542 9076 423602
rect -960 423452 480 423542
rect 9070 423540 9076 423542
rect 9140 423540 9146 423604
rect 580901 418298 580967 418301
rect 583520 418298 584960 418388
rect 580901 418296 584960 418298
rect 580901 418240 580906 418296
rect 580962 418240 584960 418296
rect 580901 418238 584960 418240
rect 580901 418235 580967 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 6126 410546 6132 410548
rect -960 410486 6132 410546
rect -960 410396 480 410486
rect 6126 410484 6132 410486
rect 6196 410484 6202 410548
rect 577446 404908 577452 404972
rect 577516 404970 577522 404972
rect 583520 404970 584960 405060
rect 577516 404910 584960 404970
rect 577516 404908 577522 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 15142 397490 15148 397492
rect -960 397430 15148 397490
rect -960 397340 480 397430
rect 15142 397428 15148 397430
rect 15212 397428 15218 397492
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580901 378450 580967 378453
rect 583520 378450 584960 378540
rect 580901 378448 584960 378450
rect 580901 378392 580906 378448
rect 580962 378392 584960 378448
rect 580901 378390 584960 378392
rect 580901 378387 580967 378390
rect 583520 378300 584960 378390
rect 54 371588 60 371652
rect 124 371588 130 371652
rect 62 371514 122 371588
rect 62 371468 674 371514
rect -960 371454 674 371468
rect -960 371378 480 371454
rect 614 371378 674 371454
rect -960 371318 674 371378
rect -960 371228 480 371318
rect 580901 365122 580967 365125
rect 583520 365122 584960 365212
rect 580901 365120 584960 365122
rect 580901 365064 580906 365120
rect 580962 365064 584960 365120
rect 580901 365062 584960 365064
rect 580901 365059 580967 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 9806 358458 9812 358460
rect -960 358398 9812 358458
rect -960 358308 480 358398
rect 9806 358396 9812 358398
rect 9876 358396 9882 358460
rect 577630 351868 577636 351932
rect 577700 351930 577706 351932
rect 583520 351930 584960 352020
rect 577700 351870 584960 351930
rect 577700 351868 577706 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3550 345402 3556 345404
rect -960 345342 3556 345402
rect -960 345252 480 345342
rect 3550 345340 3556 345342
rect 3620 345340 3626 345404
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580901 325274 580967 325277
rect 583520 325274 584960 325364
rect 580901 325272 584960 325274
rect 580901 325216 580906 325272
rect 580962 325216 584960 325272
rect 580901 325214 584960 325216
rect 580901 325211 580967 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 7598 319290 7604 319292
rect -960 319230 7604 319290
rect -960 319140 480 319230
rect 7598 319228 7604 319230
rect 7668 319228 7674 319292
rect 580901 312082 580967 312085
rect 583520 312082 584960 312172
rect 580901 312080 584960 312082
rect 580901 312024 580906 312080
rect 580962 312024 584960 312080
rect 580901 312022 584960 312024
rect 580901 312019 580967 312022
rect 583520 311932 584960 312022
rect 3366 306988 3372 307052
rect 3436 307050 3442 307052
rect 16614 307050 16620 307052
rect 3436 306990 16620 307050
rect 3436 306988 3442 306990
rect 16614 306988 16620 306990
rect 16684 306988 16690 307052
rect -960 306234 480 306324
rect 3734 306234 3740 306236
rect -960 306174 3740 306234
rect -960 306084 480 306174
rect 3734 306172 3740 306174
rect 3804 306172 3810 306236
rect 580206 298692 580212 298756
rect 580276 298754 580282 298756
rect 583520 298754 584960 298844
rect 580276 298694 584960 298754
rect 580276 298692 580282 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 2078 293178 2084 293180
rect -960 293118 2084 293178
rect -960 293028 480 293118
rect 2078 293116 2084 293118
rect 2148 293116 2154 293180
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580901 272234 580967 272237
rect 583520 272234 584960 272324
rect 580901 272232 584960 272234
rect 580901 272176 580906 272232
rect 580962 272176 584960 272232
rect 580901 272174 584960 272176
rect 580901 272171 580967 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3366 267202 3372 267204
rect -960 267142 3372 267202
rect -960 267052 480 267142
rect 3366 267140 3372 267142
rect 3436 267140 3442 267204
rect 580901 258906 580967 258909
rect 583520 258906 584960 258996
rect 580901 258904 584960 258906
rect 580901 258848 580906 258904
rect 580962 258848 584960 258904
rect 580901 258846 584960 258848
rect 580901 258843 580967 258846
rect 583520 258756 584960 258846
rect 3734 256668 3740 256732
rect 3804 256730 3810 256732
rect 6310 256730 6316 256732
rect 3804 256670 6316 256730
rect 3804 256668 3810 256670
rect 6310 256668 6316 256670
rect 6380 256668 6386 256732
rect -960 254146 480 254236
rect 2998 254220 3004 254284
rect 3068 254282 3074 254284
rect 6177 254282 6243 254285
rect 3068 254280 6243 254282
rect 3068 254224 6182 254280
rect 6238 254224 6243 254280
rect 3068 254222 6243 254224
rect 3068 254220 3074 254222
rect 3006 254146 3066 254220
rect 6177 254219 6243 254222
rect -960 254086 3066 254146
rect -960 253996 480 254086
rect 576158 245516 576164 245580
rect 576228 245578 576234 245580
rect 583520 245578 584960 245668
rect 576228 245518 584960 245578
rect 576228 245516 576234 245518
rect 583520 245428 584960 245518
rect 1158 242796 1164 242860
rect 1228 242858 1234 242860
rect 2814 242858 2820 242860
rect 1228 242798 2820 242858
rect 1228 242796 1234 242798
rect 2814 242796 2820 242798
rect 2884 242796 2890 242860
rect -960 241090 480 241180
rect 2773 241090 2839 241093
rect -960 241088 2839 241090
rect -960 241032 2778 241088
rect 2834 241032 2839 241088
rect -960 241030 2839 241032
rect -960 240940 480 241030
rect 2773 241027 2839 241030
rect 580574 232324 580580 232388
rect 580644 232386 580650 232388
rect 583520 232386 584960 232476
rect 580644 232326 584960 232386
rect 580644 232324 580650 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580758 218996 580764 219060
rect 580828 219058 580834 219060
rect 583520 219058 584960 219148
rect 580828 218998 584960 219058
rect 580828 218996 580834 218998
rect 583520 218908 584960 218998
rect -960 214828 480 215068
rect 154113 214706 154179 214709
rect 295977 214706 296043 214709
rect 154113 214704 296043 214706
rect 154113 214648 154118 214704
rect 154174 214648 295982 214704
rect 296038 214648 296043 214704
rect 154113 214646 296043 214648
rect 154113 214643 154179 214646
rect 295977 214643 296043 214646
rect 89161 214570 89227 214573
rect 285622 214570 285628 214572
rect 89161 214568 285628 214570
rect 89161 214512 89166 214568
rect 89222 214512 285628 214568
rect 89161 214510 285628 214512
rect 89161 214507 89227 214510
rect 285622 214508 285628 214510
rect 285692 214508 285698 214572
rect 10174 213828 10180 213892
rect 10244 213890 10250 213892
rect 12382 213890 12388 213892
rect 10244 213830 12388 213890
rect 10244 213828 10250 213830
rect 12382 213828 12388 213830
rect 12452 213828 12458 213892
rect 9438 213692 9444 213756
rect 9508 213754 9514 213756
rect 11094 213754 11100 213756
rect 9508 213694 11100 213754
rect 9508 213692 9514 213694
rect 11094 213692 11100 213694
rect 11164 213692 11170 213756
rect 6678 213556 6684 213620
rect 6748 213618 6754 213620
rect 13854 213618 13860 213620
rect 6748 213558 13860 213618
rect 6748 213556 6754 213558
rect 13854 213556 13860 213558
rect 13924 213556 13930 213620
rect 5390 213420 5396 213484
rect 5460 213482 5466 213484
rect 15142 213482 15148 213484
rect 5460 213422 15148 213482
rect 5460 213420 5466 213422
rect 15142 213420 15148 213422
rect 15212 213420 15218 213484
rect 2630 213284 2636 213348
rect 2700 213346 2706 213348
rect 17902 213346 17908 213348
rect 2700 213286 17908 213346
rect 2700 213284 2706 213286
rect 17902 213284 17908 213286
rect 17972 213284 17978 213348
rect 301497 213346 301563 213349
rect 413645 213346 413711 213349
rect 301497 213344 413711 213346
rect 301497 213288 301502 213344
rect 301558 213288 413650 213344
rect 413706 213288 413711 213344
rect 301497 213286 413711 213288
rect 301497 213283 301563 213286
rect 413645 213283 413711 213286
rect 974 213148 980 213212
rect 1044 213210 1050 213212
rect 16614 213210 16620 213212
rect 1044 213150 16620 213210
rect 1044 213148 1050 213150
rect 16614 213148 16620 213150
rect 16684 213148 16690 213212
rect 218973 213210 219039 213213
rect 290457 213210 290523 213213
rect 218973 213208 290523 213210
rect 218973 213152 218978 213208
rect 219034 213152 290462 213208
rect 290518 213152 290523 213208
rect 218973 213150 290523 213152
rect 218973 213147 219039 213150
rect 290457 213147 290523 213150
rect 298829 213210 298895 213213
rect 478505 213210 478571 213213
rect 298829 213208 478571 213210
rect 298829 213152 298834 213208
rect 298890 213152 478510 213208
rect 478566 213152 478571 213208
rect 298829 213150 478571 213152
rect 298829 213147 298895 213150
rect 478505 213147 478571 213150
rect 288198 210292 288204 210356
rect 288268 210354 288274 210356
rect 298829 210354 298895 210357
rect 288268 210352 298895 210354
rect 288268 210296 298834 210352
rect 298890 210296 298895 210352
rect 288268 210294 298895 210296
rect 288268 210292 288274 210294
rect 298829 210291 298895 210294
rect 583520 205580 584960 205820
rect -960 201922 480 202012
rect 2998 201922 3004 201924
rect -960 201862 3004 201922
rect -960 201772 480 201862
rect 2998 201860 3004 201862
rect 3068 201860 3074 201924
rect 8150 196012 8156 196076
rect 8220 196074 8226 196076
rect 9806 196074 9812 196076
rect 8220 196014 9812 196074
rect 8220 196012 8226 196014
rect 9806 196012 9812 196014
rect 9876 196012 9882 196076
rect 7966 194516 7972 194580
rect 8036 194578 8042 194580
rect 10174 194578 10180 194580
rect 8036 194518 10180 194578
rect 8036 194516 8042 194518
rect 10174 194516 10180 194518
rect 10244 194516 10250 194580
rect 289670 192476 289676 192540
rect 289740 192538 289746 192540
rect 301497 192538 301563 192541
rect 289740 192536 301563 192538
rect 289740 192480 301502 192536
rect 301558 192480 301563 192536
rect 289740 192478 301563 192480
rect 289740 192476 289746 192478
rect 301497 192475 301563 192478
rect 580574 192476 580580 192540
rect 580644 192538 580650 192540
rect 583520 192538 584960 192628
rect 580644 192478 584960 192538
rect 580644 192476 580650 192478
rect 583520 192388 584960 192478
rect 282862 192204 282868 192268
rect 282932 192266 282938 192268
rect 298134 192266 298140 192268
rect 282932 192206 298140 192266
rect 282932 192204 282938 192206
rect 298134 192204 298140 192206
rect 298204 192204 298210 192268
rect 284518 192068 284524 192132
rect 284588 192130 284594 192132
rect 296713 192130 296779 192133
rect 284588 192128 296779 192130
rect 284588 192072 296718 192128
rect 296774 192072 296779 192128
rect 284588 192070 296779 192072
rect 284588 192068 284594 192070
rect 296713 192067 296779 192070
rect 281022 191932 281028 191996
rect 281092 191994 281098 191996
rect 295190 191994 295196 191996
rect 281092 191934 295196 191994
rect 281092 191932 281098 191934
rect 295190 191932 295196 191934
rect 295260 191932 295266 191996
rect 297950 191858 297956 191860
rect 287010 191798 297956 191858
rect 282913 191722 282979 191725
rect 287010 191722 287070 191798
rect 297950 191796 297956 191798
rect 298020 191796 298026 191860
rect 282913 191720 287070 191722
rect 282913 191664 282918 191720
rect 282974 191664 287070 191720
rect 282913 191662 287070 191664
rect 282913 191659 282979 191662
rect 282126 191524 282132 191588
rect 282196 191586 282202 191588
rect 286174 191586 286180 191588
rect 282196 191526 286180 191586
rect 282196 191524 282202 191526
rect 286174 191524 286180 191526
rect 286244 191524 286250 191588
rect 9673 191042 9739 191045
rect 42793 191042 42859 191045
rect 9673 191040 42859 191042
rect 9673 190984 9678 191040
rect 9734 190984 42798 191040
rect 42854 190984 42859 191040
rect 9673 190982 42859 190984
rect 9673 190979 9739 190982
rect 42793 190979 42859 190982
rect 295190 190844 295196 190908
rect 295260 190906 295266 190908
rect 300301 190906 300367 190909
rect 295260 190904 300367 190906
rect 295260 190848 300306 190904
rect 300362 190848 300367 190904
rect 295260 190846 300367 190848
rect 295260 190844 295266 190846
rect 300301 190843 300367 190846
rect 287053 190770 287119 190773
rect 300761 190770 300827 190773
rect 287053 190768 300827 190770
rect 287053 190712 287058 190768
rect 287114 190712 300766 190768
rect 300822 190712 300827 190768
rect 287053 190710 300827 190712
rect 287053 190707 287119 190710
rect 300761 190707 300827 190710
rect 283966 190572 283972 190636
rect 284036 190634 284042 190636
rect 296294 190634 296300 190636
rect 284036 190574 296300 190634
rect 284036 190572 284042 190574
rect 296294 190572 296300 190574
rect 296364 190572 296370 190636
rect 300894 190498 300900 190500
rect 286366 190438 300900 190498
rect 285438 190300 285444 190364
rect 285508 190362 285514 190364
rect 286366 190362 286426 190438
rect 300894 190436 300900 190438
rect 300964 190436 300970 190500
rect 285508 190302 286426 190362
rect 285508 190300 285514 190302
rect 282678 189620 282684 189684
rect 282748 189682 282754 189684
rect 289721 189682 289787 189685
rect 282748 189680 289787 189682
rect 282748 189624 289726 189680
rect 289782 189624 289787 189680
rect 282748 189622 289787 189624
rect 282748 189620 282754 189622
rect 289721 189619 289787 189622
rect 283782 189484 283788 189548
rect 283852 189546 283858 189548
rect 297030 189546 297036 189548
rect 283852 189486 297036 189546
rect 283852 189484 283858 189486
rect 297030 189484 297036 189486
rect 297100 189484 297106 189548
rect 288014 189348 288020 189412
rect 288084 189410 288090 189412
rect 298686 189410 298692 189412
rect 288084 189350 298692 189410
rect 288084 189348 288090 189350
rect 298686 189348 298692 189350
rect 298756 189348 298762 189412
rect 284150 189212 284156 189276
rect 284220 189274 284226 189276
rect 296621 189274 296687 189277
rect 284220 189272 296687 189274
rect 284220 189216 296626 189272
rect 296682 189216 296687 189272
rect 284220 189214 296687 189216
rect 284220 189212 284226 189214
rect 296621 189211 296687 189214
rect 298134 189212 298140 189276
rect 298204 189274 298210 189276
rect 301446 189274 301452 189276
rect 298204 189214 301452 189274
rect 298204 189212 298210 189214
rect 301446 189212 301452 189214
rect 301516 189212 301522 189276
rect 9622 189076 9628 189140
rect 9692 189138 9698 189140
rect 9765 189138 9831 189141
rect 285673 189138 285739 189141
rect 289854 189138 289860 189140
rect 9692 189136 9831 189138
rect 9692 189080 9770 189136
rect 9826 189080 9831 189136
rect 9692 189078 9831 189080
rect 281704 189078 281826 189138
rect 9692 189076 9698 189078
rect 9765 189075 9831 189078
rect 281766 189002 281826 189078
rect 285673 189136 289860 189138
rect 285673 189080 285678 189136
rect 285734 189080 289860 189136
rect 285673 189078 289860 189080
rect 285673 189075 285739 189078
rect 289854 189076 289860 189078
rect 289924 189138 289930 189140
rect 299422 189138 299428 189140
rect 289924 189078 299428 189138
rect 289924 189076 289930 189078
rect 299422 189076 299428 189078
rect 299492 189076 299498 189140
rect 300761 189138 300827 189141
rect 301262 189138 301268 189140
rect 300761 189136 301268 189138
rect 300761 189080 300766 189136
rect 300822 189080 301268 189136
rect 300761 189078 301268 189080
rect 300761 189075 300827 189078
rect 301262 189076 301268 189078
rect 301332 189076 301338 189140
rect 302325 189138 302391 189141
rect 302325 189136 302496 189138
rect 302325 189080 302330 189136
rect 302386 189080 302496 189136
rect 302325 189078 302496 189080
rect 302325 189075 302391 189078
rect -960 188866 480 188956
rect 281612 188942 281826 189002
rect 302650 188942 302772 189002
rect 2814 188866 2820 188868
rect -960 188806 2820 188866
rect -960 188716 480 188806
rect 2814 188804 2820 188806
rect 2884 188804 2890 188868
rect 281674 188866 281734 188942
rect 302650 188866 302710 188942
rect 281490 188806 281734 188866
rect 302588 188806 302710 188866
rect 281490 188730 281550 188806
rect 302650 188730 302710 188806
rect 281428 188670 281550 188730
rect 302588 188670 302710 188730
rect 281490 188594 281550 188670
rect 302650 188594 302710 188670
rect 281428 188534 281826 188594
rect 281766 188322 281826 188534
rect 302190 188534 302772 188594
rect 290958 188396 290964 188460
rect 291028 188458 291034 188460
rect 299606 188458 299612 188460
rect 291028 188398 299612 188458
rect 291028 188396 291034 188398
rect 299606 188396 299612 188398
rect 299676 188396 299682 188460
rect 281612 188262 281826 188322
rect 282310 188260 282316 188324
rect 282380 188322 282386 188324
rect 287053 188322 287119 188325
rect 282380 188320 287119 188322
rect 282380 188264 287058 188320
rect 287114 188264 287119 188320
rect 282380 188262 287119 188264
rect 282380 188260 282386 188262
rect 287053 188259 287119 188262
rect 289721 188322 289787 188325
rect 293166 188322 293172 188324
rect 289721 188320 293172 188322
rect 289721 188264 289726 188320
rect 289782 188264 293172 188320
rect 289721 188262 293172 188264
rect 289721 188259 289787 188262
rect 293166 188260 293172 188262
rect 293236 188322 293242 188324
rect 301078 188322 301084 188324
rect 293236 188262 301084 188322
rect 293236 188260 293242 188262
rect 301078 188260 301084 188262
rect 301148 188260 301154 188324
rect 302190 188322 302250 188534
rect 302325 188458 302391 188461
rect 302325 188456 302588 188458
rect 302325 188400 302330 188456
rect 302386 188400 302588 188456
rect 302325 188398 302588 188400
rect 302325 188395 302391 188398
rect 302190 188262 302588 188322
rect 293534 188186 293540 188188
rect 281704 188126 293540 188186
rect 293534 188124 293540 188126
rect 293604 188186 293610 188188
rect 293604 188126 302496 188186
rect 293604 188124 293610 188126
rect 299054 188050 299060 188052
rect 281612 187990 299060 188050
rect 299054 187988 299060 187990
rect 299124 188050 299130 188052
rect 299124 187990 302588 188050
rect 299124 187988 299130 187990
rect 292430 187914 292436 187916
rect 281612 187854 292436 187914
rect 292430 187852 292436 187854
rect 292500 187914 292506 187916
rect 292500 187854 302588 187914
rect 292500 187852 292506 187854
rect 290958 187778 290964 187780
rect 281612 187718 290964 187778
rect 290958 187716 290964 187718
rect 291028 187716 291034 187780
rect 295006 187716 295012 187780
rect 295076 187778 295082 187780
rect 299238 187778 299244 187780
rect 295076 187718 299244 187778
rect 295076 187716 295082 187718
rect 299238 187716 299244 187718
rect 299308 187716 299314 187780
rect 299606 187716 299612 187780
rect 299676 187778 299682 187780
rect 299676 187718 302588 187778
rect 299676 187716 299682 187718
rect 283281 187642 283347 187645
rect 281612 187640 283347 187642
rect 281612 187584 283286 187640
rect 283342 187584 283347 187640
rect 281612 187582 283347 187584
rect 283281 187579 283347 187582
rect 299422 187580 299428 187644
rect 299492 187642 299498 187644
rect 299492 187582 302588 187642
rect 299492 187580 299498 187582
rect 285438 187506 285444 187508
rect 281612 187446 285444 187506
rect 285438 187444 285444 187446
rect 285508 187444 285514 187508
rect 300894 187444 300900 187508
rect 300964 187506 300970 187508
rect 300964 187446 302588 187506
rect 300964 187444 300970 187446
rect 282494 187370 282500 187372
rect 281612 187310 282500 187370
rect 282494 187308 282500 187310
rect 282564 187308 282570 187372
rect 285622 187308 285628 187372
rect 285692 187370 285698 187372
rect 286961 187370 287027 187373
rect 285692 187368 287027 187370
rect 285692 187312 286966 187368
rect 287022 187312 287027 187368
rect 285692 187310 287027 187312
rect 285692 187308 285698 187310
rect 286961 187307 287027 187310
rect 300894 187308 300900 187372
rect 300964 187370 300970 187372
rect 301446 187370 301452 187372
rect 300964 187310 301452 187370
rect 300964 187308 300970 187310
rect 301446 187308 301452 187310
rect 301516 187370 301522 187372
rect 301516 187310 302588 187370
rect 301516 187308 301522 187310
rect 299974 187234 299980 187236
rect 281612 187174 299980 187234
rect 299974 187172 299980 187174
rect 300044 187234 300050 187236
rect 300044 187174 302588 187234
rect 300044 187172 300050 187174
rect 299749 187098 299815 187101
rect 281612 187096 302588 187098
rect 281612 187040 299754 187096
rect 299810 187040 302588 187096
rect 281612 187038 302588 187040
rect 299749 187035 299815 187038
rect 299238 186962 299244 186964
rect 281612 186902 299244 186962
rect 299238 186900 299244 186902
rect 299308 186962 299314 186964
rect 299308 186902 302588 186962
rect 299308 186900 299314 186902
rect 298870 186826 298876 186828
rect 281612 186766 298876 186826
rect 298870 186764 298876 186766
rect 298940 186826 298946 186828
rect 298940 186766 302588 186826
rect 298940 186764 298946 186766
rect 282310 186690 282316 186692
rect 281612 186630 282316 186690
rect 282310 186628 282316 186630
rect 282380 186628 282386 186692
rect 286358 186628 286364 186692
rect 286428 186690 286434 186692
rect 299606 186690 299612 186692
rect 286428 186630 299612 186690
rect 286428 186628 286434 186630
rect 299606 186628 299612 186630
rect 299676 186628 299682 186692
rect 301262 186628 301268 186692
rect 301332 186690 301338 186692
rect 301332 186630 302588 186690
rect 301332 186628 301338 186630
rect 288014 186554 288020 186556
rect 281612 186494 288020 186554
rect 288014 186492 288020 186494
rect 288084 186492 288090 186556
rect 298134 186492 298140 186556
rect 298204 186554 298210 186556
rect 298686 186554 298692 186556
rect 298204 186494 298692 186554
rect 298204 186492 298210 186494
rect 298686 186492 298692 186494
rect 298756 186554 298762 186556
rect 298756 186494 302588 186554
rect 298756 186492 298762 186494
rect 282821 186418 282887 186421
rect 297398 186418 297404 186420
rect 281612 186416 282887 186418
rect 281612 186360 282826 186416
rect 282882 186360 282887 186416
rect 281612 186358 282887 186360
rect 282821 186355 282887 186358
rect 284158 186358 297404 186418
rect 284158 186282 284218 186358
rect 297398 186356 297404 186358
rect 297468 186418 297474 186420
rect 297468 186358 297834 186418
rect 297468 186356 297474 186358
rect 281704 186222 284218 186282
rect 297774 186282 297834 186358
rect 297950 186356 297956 186420
rect 298020 186418 298026 186420
rect 298020 186358 302588 186418
rect 298020 186356 298026 186358
rect 297774 186222 302496 186282
rect 283782 186146 283788 186148
rect 281612 186086 283788 186146
rect 283782 186084 283788 186086
rect 283852 186084 283858 186148
rect 284017 186146 284083 186149
rect 293902 186146 293908 186148
rect 284017 186144 293908 186146
rect 284017 186088 284022 186144
rect 284078 186088 293908 186144
rect 284017 186086 293908 186088
rect 284017 186083 284083 186086
rect 293902 186084 293908 186086
rect 293972 186084 293978 186148
rect 297030 186084 297036 186148
rect 297100 186146 297106 186148
rect 297100 186086 302588 186146
rect 297100 186084 297106 186086
rect 284150 186010 284156 186012
rect 281612 185950 284156 186010
rect 284150 185948 284156 185950
rect 284220 185948 284226 186012
rect 295190 185948 295196 186012
rect 295260 186010 295266 186012
rect 296478 186010 296484 186012
rect 295260 185950 296484 186010
rect 295260 185948 295266 185950
rect 296478 185948 296484 185950
rect 296548 185948 296554 186012
rect 296621 186010 296687 186013
rect 296621 186008 302588 186010
rect 296621 185952 296626 186008
rect 296682 185952 302588 186008
rect 296621 185950 302588 185952
rect 296621 185947 296687 185950
rect 283966 185874 283972 185876
rect 281612 185814 283972 185874
rect 283966 185812 283972 185814
rect 284036 185812 284042 185876
rect 296294 185812 296300 185876
rect 296364 185874 296370 185876
rect 296364 185814 302588 185874
rect 296364 185812 296370 185814
rect 282729 185738 282795 185741
rect 281612 185736 282795 185738
rect 281612 185680 282734 185736
rect 282790 185680 282795 185736
rect 281612 185678 282795 185680
rect 282729 185675 282795 185678
rect 282862 185676 282868 185740
rect 282932 185738 282938 185740
rect 291326 185738 291332 185740
rect 282932 185678 291332 185738
rect 282932 185676 282938 185678
rect 291326 185676 291332 185678
rect 291396 185676 291402 185740
rect 292941 185738 293007 185741
rect 295006 185738 295012 185740
rect 292941 185736 295012 185738
rect 292941 185680 292946 185736
rect 293002 185680 295012 185736
rect 292941 185678 295012 185680
rect 292941 185675 293007 185678
rect 295006 185676 295012 185678
rect 295076 185676 295082 185740
rect 298001 185738 298067 185741
rect 296486 185736 298067 185738
rect 296486 185680 298006 185736
rect 298062 185680 298067 185736
rect 296486 185678 298067 185680
rect 293861 185602 293927 185605
rect 295926 185602 295932 185604
rect 281612 185542 293786 185602
rect 292941 185466 293007 185469
rect 281612 185464 293007 185466
rect 281612 185408 292946 185464
rect 293002 185408 293007 185464
rect 281612 185406 293007 185408
rect 293726 185466 293786 185542
rect 293861 185600 295932 185602
rect 293861 185544 293866 185600
rect 293922 185544 295932 185600
rect 293861 185542 295932 185544
rect 293861 185539 293927 185542
rect 295926 185540 295932 185542
rect 295996 185602 296002 185604
rect 296486 185602 296546 185678
rect 298001 185675 298067 185678
rect 299749 185740 299815 185741
rect 299749 185736 299796 185740
rect 299860 185738 299866 185740
rect 300853 185738 300919 185741
rect 299749 185680 299754 185736
rect 299749 185676 299796 185680
rect 299860 185678 299906 185738
rect 300853 185736 302588 185738
rect 300853 185680 300858 185736
rect 300914 185680 302588 185736
rect 300853 185678 302588 185680
rect 299860 185676 299866 185678
rect 299749 185675 299815 185676
rect 300853 185675 300919 185678
rect 295996 185542 296546 185602
rect 296670 185542 302588 185602
rect 295996 185540 296002 185542
rect 295558 185466 295564 185468
rect 293726 185406 295564 185466
rect 292941 185403 293007 185406
rect 295558 185404 295564 185406
rect 295628 185466 295634 185468
rect 296670 185466 296730 185542
rect 295628 185406 296730 185466
rect 295628 185404 295634 185406
rect 299422 185404 299428 185468
rect 299492 185466 299498 185468
rect 299492 185406 302588 185466
rect 299492 185404 299498 185406
rect 294822 185330 294828 185332
rect 281612 185270 294828 185330
rect 294822 185268 294828 185270
rect 294892 185330 294898 185332
rect 294892 185270 302588 185330
rect 294892 185268 294898 185270
rect 294454 185194 294460 185196
rect 281612 185134 294460 185194
rect 294454 185132 294460 185134
rect 294524 185194 294530 185196
rect 294524 185134 302588 185194
rect 294524 185132 294530 185134
rect 284017 185058 284083 185061
rect 281612 185056 284083 185058
rect 281612 185000 284022 185056
rect 284078 185000 284083 185056
rect 281612 184998 284083 185000
rect 284017 184995 284083 184998
rect 284158 184998 292682 185058
rect 284158 184922 284218 184998
rect 281612 184862 284218 184922
rect 285438 184860 285444 184924
rect 285508 184922 285514 184924
rect 286542 184922 286548 184924
rect 285508 184862 286548 184922
rect 285508 184860 285514 184862
rect 286542 184860 286548 184862
rect 286612 184860 286618 184924
rect 291142 184860 291148 184924
rect 291212 184922 291218 184924
rect 292481 184922 292547 184925
rect 291212 184920 292547 184922
rect 291212 184864 292486 184920
rect 292542 184864 292547 184920
rect 291212 184862 292547 184864
rect 292622 184922 292682 184998
rect 293902 184996 293908 185060
rect 293972 185058 293978 185060
rect 293972 184998 302588 185058
rect 293972 184996 293978 184998
rect 293718 184922 293724 184924
rect 292622 184862 293724 184922
rect 291212 184860 291218 184862
rect 292481 184859 292547 184862
rect 293718 184860 293724 184862
rect 293788 184922 293794 184924
rect 293788 184862 302588 184922
rect 293788 184860 293794 184862
rect 293217 184788 293283 184789
rect 282678 184786 282684 184788
rect 281612 184726 282684 184786
rect 282678 184724 282684 184726
rect 282748 184724 282754 184788
rect 293166 184724 293172 184788
rect 293236 184786 293283 184788
rect 293236 184784 293328 184786
rect 293278 184728 293328 184784
rect 293236 184726 293328 184728
rect 293236 184724 293283 184726
rect 301078 184724 301084 184788
rect 301148 184786 301154 184788
rect 301148 184726 302588 184786
rect 301148 184724 301154 184726
rect 293217 184723 293283 184724
rect 292982 184650 292988 184652
rect 281612 184590 292988 184650
rect 292982 184588 292988 184590
rect 293052 184650 293058 184652
rect 293052 184590 302588 184650
rect 293052 184588 293058 184590
rect 282862 184514 282868 184516
rect 281612 184454 282868 184514
rect 282862 184452 282868 184454
rect 282932 184452 282938 184516
rect 291326 184452 291332 184516
rect 291396 184514 291402 184516
rect 292614 184514 292620 184516
rect 291396 184454 292620 184514
rect 291396 184452 291402 184454
rect 292614 184452 292620 184454
rect 292684 184514 292690 184516
rect 292684 184454 302588 184514
rect 292684 184452 292690 184454
rect 282545 184378 282611 184381
rect 281612 184376 282611 184378
rect 281612 184320 282550 184376
rect 282606 184320 282611 184376
rect 281612 184318 282611 184320
rect 282545 184315 282611 184318
rect 282913 184378 282979 184381
rect 284518 184378 284524 184380
rect 282913 184376 284524 184378
rect 282913 184320 282918 184376
rect 282974 184320 284524 184376
rect 282913 184318 284524 184320
rect 282913 184315 282979 184318
rect 284518 184316 284524 184318
rect 284588 184316 284594 184380
rect 285581 184378 285647 184381
rect 292573 184378 292639 184381
rect 285581 184376 292639 184378
rect 285581 184320 285586 184376
rect 285642 184320 292578 184376
rect 292634 184320 292639 184376
rect 285581 184318 292639 184320
rect 285581 184315 285647 184318
rect 292573 184315 292639 184318
rect 300853 184378 300919 184381
rect 300853 184376 302588 184378
rect 300853 184320 300858 184376
rect 300914 184320 302588 184376
rect 300853 184318 302588 184320
rect 300853 184315 300919 184318
rect 291878 184242 291884 184244
rect 281704 184182 291884 184242
rect 291878 184180 291884 184182
rect 291948 184242 291954 184244
rect 291948 184182 302496 184242
rect 291948 184180 291954 184182
rect 291510 184106 291516 184108
rect 281704 184046 291516 184106
rect 291510 184044 291516 184046
rect 291580 184106 291586 184108
rect 291580 184046 302496 184106
rect 291580 184044 291586 184046
rect 290406 183970 290412 183972
rect 281612 183910 290412 183970
rect 290406 183908 290412 183910
rect 290476 183970 290482 183972
rect 290476 183910 302588 183970
rect 290476 183908 290482 183910
rect 290038 183834 290044 183836
rect 281612 183774 290044 183834
rect 290038 183772 290044 183774
rect 290108 183834 290114 183836
rect 290108 183774 302588 183834
rect 290108 183772 290114 183774
rect 281022 183636 281028 183700
rect 281092 183636 281098 183700
rect 284334 183636 284340 183700
rect 284404 183698 284410 183700
rect 285581 183698 285647 183701
rect 284404 183696 285647 183698
rect 284404 183640 285586 183696
rect 285642 183640 285647 183696
rect 284404 183638 285647 183640
rect 284404 183636 284410 183638
rect 285581 183635 285647 183638
rect 288206 183638 288634 183698
rect 288206 183562 288266 183638
rect 288433 183564 288499 183565
rect 288382 183562 288388 183564
rect 281612 183502 288266 183562
rect 288342 183502 288388 183562
rect 288452 183560 288499 183564
rect 288494 183504 288499 183560
rect 288382 183500 288388 183502
rect 288452 183500 288499 183504
rect 288574 183562 288634 183638
rect 292246 183636 292252 183700
rect 292316 183698 292322 183700
rect 292573 183698 292639 183701
rect 292316 183696 292639 183698
rect 292316 183640 292578 183696
rect 292634 183640 292639 183696
rect 292316 183638 292639 183640
rect 292316 183636 292322 183638
rect 292573 183635 292639 183638
rect 300301 183698 300367 183701
rect 300301 183696 302588 183698
rect 300301 183640 300306 183696
rect 300362 183640 302588 183696
rect 300301 183638 302588 183640
rect 300301 183635 300367 183638
rect 289302 183562 289308 183564
rect 288574 183502 289308 183562
rect 289302 183500 289308 183502
rect 289372 183562 289378 183564
rect 289372 183502 302588 183562
rect 289372 183500 289378 183502
rect 288433 183499 288499 183500
rect 288934 183426 288940 183428
rect 281612 183366 288940 183426
rect 288934 183364 288940 183366
rect 289004 183426 289010 183428
rect 289004 183366 302588 183426
rect 289004 183364 289010 183366
rect 288566 183290 288572 183292
rect 281612 183230 288572 183290
rect 288566 183228 288572 183230
rect 288636 183290 288642 183292
rect 288636 183230 302588 183290
rect 288636 183228 288642 183230
rect 288014 183154 288020 183156
rect 281612 183094 288020 183154
rect 288014 183092 288020 183094
rect 288084 183154 288090 183156
rect 288341 183154 288407 183157
rect 288084 183152 288407 183154
rect 288084 183096 288346 183152
rect 288402 183096 288407 183152
rect 288084 183094 288407 183096
rect 288084 183092 288090 183094
rect 288341 183091 288407 183094
rect 300853 183154 300919 183157
rect 300853 183152 302588 183154
rect 300853 183096 300858 183152
rect 300914 183096 302588 183152
rect 300853 183094 302588 183096
rect 300853 183091 300919 183094
rect 287830 183018 287836 183020
rect 281612 182958 287836 183018
rect 287830 182956 287836 182958
rect 287900 183018 287906 183020
rect 287900 182958 302588 183018
rect 287900 182956 287906 182958
rect 287462 182882 287468 182884
rect 281612 182822 287468 182882
rect 287462 182820 287468 182822
rect 287532 182882 287538 182884
rect 287532 182822 302588 182882
rect 287532 182820 287538 182822
rect 287094 182746 287100 182748
rect 281612 182686 287100 182746
rect 287094 182684 287100 182686
rect 287164 182746 287170 182748
rect 287164 182686 302588 182746
rect 287164 182684 287170 182686
rect 282913 182610 282979 182613
rect 281612 182608 282979 182610
rect 281612 182552 282918 182608
rect 282974 182552 282979 182608
rect 281612 182550 282979 182552
rect 282913 182547 282979 182550
rect 287053 182610 287119 182613
rect 288198 182610 288204 182612
rect 287053 182608 288204 182610
rect 287053 182552 287058 182608
rect 287114 182552 288204 182608
rect 287053 182550 288204 182552
rect 287053 182547 287119 182550
rect 288198 182548 288204 182550
rect 288268 182548 288274 182612
rect 301262 182548 301268 182612
rect 301332 182610 301338 182612
rect 301332 182550 302588 182610
rect 301332 182548 301338 182550
rect 286358 182474 286364 182476
rect 281612 182414 286364 182474
rect 286358 182412 286364 182414
rect 286428 182412 286434 182476
rect 299606 182412 299612 182476
rect 299676 182474 299682 182476
rect 299676 182414 302588 182474
rect 299676 182412 299682 182414
rect 285990 182338 285996 182340
rect 281612 182278 285996 182338
rect 285990 182276 285996 182278
rect 286060 182338 286066 182340
rect 286060 182278 302588 182338
rect 286060 182276 286066 182278
rect 283005 182202 283071 182205
rect 281612 182200 283071 182202
rect 281612 182144 283010 182200
rect 283066 182144 283071 182200
rect 281612 182142 283071 182144
rect 283005 182139 283071 182142
rect 302233 182202 302299 182205
rect 302233 182200 302588 182202
rect 302233 182144 302238 182200
rect 302294 182144 302588 182200
rect 302233 182142 302588 182144
rect 302233 182139 302299 182142
rect 285254 182066 285260 182068
rect 281612 182006 285260 182066
rect 285254 182004 285260 182006
rect 285324 182066 285330 182068
rect 285324 182006 302588 182066
rect 285324 182004 285330 182006
rect 284886 181930 284892 181932
rect 281612 181870 284892 181930
rect 284886 181868 284892 181870
rect 284956 181930 284962 181932
rect 284956 181870 302588 181930
rect 284956 181868 284962 181870
rect 284518 181794 284524 181796
rect 281612 181734 284524 181794
rect 284518 181732 284524 181734
rect 284588 181794 284594 181796
rect 284588 181734 302588 181794
rect 284588 181732 284594 181734
rect 283046 181658 283052 181660
rect 281612 181598 283052 181658
rect 283046 181596 283052 181598
rect 283116 181658 283122 181660
rect 283116 181598 302588 181658
rect 283116 181596 283122 181598
rect 284334 181522 284340 181524
rect 281704 181462 284340 181522
rect 284334 181460 284340 181462
rect 284404 181522 284410 181524
rect 284404 181462 302496 181522
rect 284404 181460 284410 181462
rect 283414 181386 283420 181388
rect 281612 181326 283420 181386
rect 283414 181324 283420 181326
rect 283484 181324 283490 181388
rect 300894 181324 300900 181388
rect 300964 181386 300970 181388
rect 300964 181326 302588 181386
rect 300964 181324 300970 181326
rect 283557 181250 283623 181253
rect 281612 181248 302588 181250
rect 281612 181192 283562 181248
rect 283618 181192 302588 181248
rect 281612 181190 302588 181192
rect 283557 181187 283623 181190
rect 281574 181052 281580 181116
rect 281644 181114 281650 181116
rect 282729 181114 282795 181117
rect 281644 181112 282795 181114
rect 281644 181056 282734 181112
rect 282790 181056 282795 181112
rect 281644 181054 282795 181056
rect 281644 181052 281650 181054
rect 282729 181051 282795 181054
rect 300945 181114 301011 181117
rect 300945 181112 302588 181114
rect 300945 181056 300950 181112
rect 301006 181056 302588 181112
rect 300945 181054 302588 181056
rect 300945 181051 301011 181054
rect 281809 180978 281875 180981
rect 281612 180976 281875 180978
rect 281612 180920 281814 180976
rect 281870 180920 281875 180976
rect 281612 180918 281875 180920
rect 281809 180915 281875 180918
rect 301773 180978 301839 180981
rect 301773 180976 302588 180978
rect 301773 180920 301778 180976
rect 301834 180920 302588 180976
rect 301773 180918 302588 180920
rect 301773 180915 301839 180918
rect 281942 180842 281948 180844
rect 281612 180782 281948 180842
rect 281942 180780 281948 180782
rect 282012 180842 282018 180844
rect 282361 180842 282427 180845
rect 296621 180842 296687 180845
rect 296846 180842 296852 180844
rect 282012 180840 282427 180842
rect 282012 180784 282366 180840
rect 282422 180784 282427 180840
rect 282012 180782 282427 180784
rect 296576 180840 296852 180842
rect 296576 180784 296626 180840
rect 296682 180784 296852 180840
rect 296576 180782 296852 180784
rect 282012 180780 282018 180782
rect 282361 180779 282427 180782
rect 296621 180779 296687 180782
rect 296846 180780 296852 180782
rect 296916 180780 296922 180844
rect 300853 180842 300919 180845
rect 300853 180840 302588 180842
rect 300853 180784 300858 180840
rect 300914 180784 302588 180840
rect 300853 180782 302588 180784
rect 300853 180779 300919 180782
rect 282494 180706 282500 180708
rect 281612 180646 282500 180706
rect 282494 180644 282500 180646
rect 282564 180706 282570 180708
rect 282564 180646 302588 180706
rect 282564 180644 282570 180646
rect 282862 180570 282868 180572
rect 281612 180510 282868 180570
rect 282862 180508 282868 180510
rect 282932 180570 282938 180572
rect 282932 180510 302588 180570
rect 282932 180508 282938 180510
rect 283414 180372 283420 180436
rect 283484 180434 283490 180436
rect 300894 180434 300900 180436
rect 283484 180374 300900 180434
rect 283484 180372 283490 180374
rect 300894 180372 300900 180374
rect 300964 180372 300970 180436
rect 295241 180298 295307 180301
rect 302325 180298 302391 180301
rect 295241 180296 302391 180298
rect 295241 180240 295246 180296
rect 295302 180240 302330 180296
rect 302386 180240 302391 180296
rect 295241 180238 302391 180240
rect 295241 180235 295307 180238
rect 302325 180235 302391 180238
rect 283005 180162 283071 180165
rect 285622 180162 285628 180164
rect 283005 180160 285628 180162
rect 283005 180104 283010 180160
rect 283066 180104 285628 180160
rect 283005 180102 285628 180104
rect 283005 180099 283071 180102
rect 285622 180100 285628 180102
rect 285692 180162 285698 180164
rect 292021 180162 292087 180165
rect 285692 180160 292087 180162
rect 285692 180104 292026 180160
rect 292082 180104 292087 180160
rect 285692 180102 292087 180104
rect 285692 180100 285698 180102
rect 292021 180099 292087 180102
rect 296110 180100 296116 180164
rect 296180 180162 296186 180164
rect 296478 180162 296484 180164
rect 296180 180102 296484 180162
rect 296180 180100 296186 180102
rect 296478 180100 296484 180102
rect 296548 180100 296554 180164
rect 286542 179964 286548 180028
rect 286612 180026 286618 180028
rect 302366 180026 302372 180028
rect 286612 179966 302372 180026
rect 286612 179964 286618 179966
rect 302366 179964 302372 179966
rect 302436 179964 302442 180028
rect 293534 179828 293540 179892
rect 293604 179890 293610 179892
rect 300526 179890 300532 179892
rect 293604 179830 300532 179890
rect 293604 179828 293610 179830
rect 300526 179828 300532 179830
rect 300596 179828 300602 179892
rect 289905 179484 289971 179485
rect 289854 179482 289860 179484
rect 289814 179422 289860 179482
rect 289924 179480 289971 179484
rect 289966 179424 289971 179480
rect 289854 179420 289860 179422
rect 289924 179420 289971 179424
rect 292430 179420 292436 179484
rect 292500 179482 292506 179484
rect 292500 179422 292682 179482
rect 292500 179420 292506 179422
rect 289905 179419 289971 179420
rect 251173 179346 251239 179349
rect 281809 179346 281875 179349
rect 251173 179344 281875 179346
rect 251173 179288 251178 179344
rect 251234 179288 281814 179344
rect 281870 179288 281875 179344
rect 251173 179286 281875 179288
rect 292622 179346 292682 179422
rect 299054 179420 299060 179484
rect 299124 179482 299130 179484
rect 302366 179482 302372 179484
rect 299124 179422 302372 179482
rect 299124 179420 299130 179422
rect 302366 179420 302372 179422
rect 302436 179420 302442 179484
rect 301630 179346 301636 179348
rect 292622 179286 301636 179346
rect 251173 179283 251239 179286
rect 281809 179283 281875 179286
rect 301630 179284 301636 179286
rect 301700 179284 301706 179348
rect 580574 179148 580580 179212
rect 580644 179210 580650 179212
rect 583520 179210 584960 179300
rect 580644 179150 584960 179210
rect 580644 179148 580650 179150
rect 583520 179060 584960 179150
rect 9438 178876 9444 178940
rect 9508 178938 9514 178940
rect 43294 178938 43300 178940
rect 9508 178878 43300 178938
rect 9508 178876 9514 178878
rect 43294 178876 43300 178878
rect 43364 178876 43370 178940
rect 286174 178876 286180 178940
rect 286244 178938 286250 178940
rect 292021 178938 292087 178941
rect 302233 178938 302299 178941
rect 286244 178878 291946 178938
rect 286244 178876 286250 178878
rect 7966 178740 7972 178804
rect 8036 178802 8042 178804
rect 111006 178802 111012 178804
rect 8036 178742 111012 178802
rect 8036 178740 8042 178742
rect 111006 178740 111012 178742
rect 111076 178740 111082 178804
rect 282821 178802 282887 178805
rect 287053 178802 287119 178805
rect 282821 178800 287119 178802
rect 282821 178744 282826 178800
rect 282882 178744 287058 178800
rect 287114 178744 287119 178800
rect 282821 178742 287119 178744
rect 291886 178802 291946 178878
rect 292021 178936 302299 178938
rect 292021 178880 292026 178936
rect 292082 178880 302238 178936
rect 302294 178880 302299 178936
rect 292021 178878 302299 178880
rect 292021 178875 292087 178878
rect 302233 178875 302299 178878
rect 300158 178802 300164 178804
rect 291886 178742 300164 178802
rect 282821 178739 282887 178742
rect 287053 178739 287119 178742
rect 300158 178740 300164 178742
rect 300228 178740 300234 178804
rect 300526 178740 300532 178804
rect 300596 178802 300602 178804
rect 334750 178802 334756 178804
rect 300596 178742 334756 178802
rect 300596 178740 300602 178742
rect 334750 178740 334756 178742
rect 334820 178740 334826 178804
rect 248086 178604 248092 178668
rect 248156 178666 248162 178668
rect 281574 178666 281580 178668
rect 248156 178606 281580 178666
rect 248156 178604 248162 178606
rect 281574 178604 281580 178606
rect 281644 178604 281650 178668
rect 295977 178666 296043 178669
rect 335353 178666 335419 178669
rect 295977 178664 335419 178666
rect 295977 178608 295982 178664
rect 296038 178608 335358 178664
rect 335414 178608 335419 178664
rect 295977 178606 335419 178608
rect 295977 178603 296043 178606
rect 335353 178603 335419 178606
rect 289670 178060 289676 178124
rect 289740 178122 289746 178124
rect 296161 178122 296227 178125
rect 289740 178120 296227 178122
rect 289740 178064 296166 178120
rect 296222 178064 296227 178120
rect 289740 178062 296227 178064
rect 289740 178060 289746 178062
rect 296161 178059 296227 178062
rect 281206 177924 281212 177988
rect 281276 177986 281282 177988
rect 282862 177986 282868 177988
rect 281276 177926 282868 177986
rect 281276 177924 281282 177926
rect 282862 177924 282868 177926
rect 282932 177924 282938 177988
rect 289670 177924 289676 177988
rect 289740 177986 289746 177988
rect 296110 177986 296116 177988
rect 289740 177926 296116 177986
rect 289740 177924 289746 177926
rect 296110 177924 296116 177926
rect 296180 177924 296186 177988
rect 282913 177442 282979 177445
rect 286726 177442 286732 177444
rect 282913 177440 286732 177442
rect 282913 177384 282918 177440
rect 282974 177384 286732 177440
rect 282913 177382 286732 177384
rect 282913 177379 282979 177382
rect 286726 177380 286732 177382
rect 286796 177442 286802 177444
rect 301262 177442 301268 177444
rect 286796 177382 301268 177442
rect 286796 177380 286802 177382
rect 301262 177380 301268 177382
rect 301332 177380 301338 177444
rect 286961 177306 287027 177309
rect 301446 177306 301452 177308
rect 286961 177304 301452 177306
rect 286961 177248 286966 177304
rect 287022 177248 301452 177304
rect 286961 177246 301452 177248
rect 286961 177243 287027 177246
rect 301446 177244 301452 177246
rect 301516 177244 301522 177308
rect 299054 176700 299060 176764
rect 299124 176762 299130 176764
rect 301078 176762 301084 176764
rect 299124 176702 301084 176762
rect 299124 176700 299130 176702
rect 301078 176700 301084 176702
rect 301148 176700 301154 176764
rect 280889 176082 280955 176085
rect 288433 176082 288499 176085
rect 280889 176080 288499 176082
rect -960 175796 480 176036
rect 280889 176024 280894 176080
rect 280950 176024 288438 176080
rect 288494 176024 288499 176080
rect 280889 176022 288499 176024
rect 280889 176019 280955 176022
rect 288433 176019 288499 176022
rect 282126 175884 282132 175948
rect 282196 175946 282202 175948
rect 283046 175946 283052 175948
rect 282196 175886 283052 175946
rect 282196 175884 282202 175886
rect 283046 175884 283052 175886
rect 283116 175884 283122 175948
rect 9581 175266 9647 175269
rect 10174 175266 10180 175268
rect 9581 175264 10180 175266
rect 9581 175208 9586 175264
rect 9642 175208 10180 175264
rect 9581 175206 10180 175208
rect 9581 175203 9647 175206
rect 10174 175204 10180 175206
rect 10244 175204 10250 175268
rect 292481 174586 292547 174589
rect 303102 174586 303108 174588
rect 292481 174584 303108 174586
rect 292481 174528 292486 174584
rect 292542 174528 303108 174584
rect 292481 174526 303108 174528
rect 292481 174523 292547 174526
rect 303102 174524 303108 174526
rect 303172 174524 303178 174588
rect 573633 174586 573699 174589
rect 580574 174586 580580 174588
rect 573633 174584 580580 174586
rect 573633 174528 573638 174584
rect 573694 174528 580580 174584
rect 573633 174526 580580 174528
rect 573633 174523 573699 174526
rect 580574 174524 580580 174526
rect 580644 174524 580650 174588
rect 583520 165732 584960 165972
rect -960 162890 480 162980
rect 4102 162890 4108 162892
rect -960 162830 4108 162890
rect -960 162740 480 162830
rect 4102 162828 4108 162830
rect 4172 162828 4178 162892
rect 301630 158068 301636 158132
rect 301700 158130 301706 158132
rect 307702 158130 307708 158132
rect 301700 158070 307708 158130
rect 301700 158068 301706 158070
rect 307702 158068 307708 158070
rect 307772 158068 307778 158132
rect 277158 157932 277164 157996
rect 277228 157994 277234 157996
rect 281758 157994 281764 157996
rect 277228 157934 281764 157994
rect 277228 157932 277234 157934
rect 281758 157932 281764 157934
rect 281828 157932 281834 157996
rect 296161 157994 296227 157997
rect 306373 157994 306439 157997
rect 296161 157992 306439 157994
rect 296161 157936 296166 157992
rect 296222 157936 306378 157992
rect 306434 157936 306439 157992
rect 296161 157934 306439 157936
rect 296161 157931 296227 157934
rect 306373 157931 306439 157934
rect 10174 157388 10180 157452
rect 10244 157450 10250 157452
rect 11697 157450 11763 157453
rect 10244 157448 11763 157450
rect 10244 157392 11702 157448
rect 11758 157392 11763 157448
rect 10244 157390 11763 157392
rect 10244 157388 10250 157390
rect 11697 157387 11763 157390
rect 279918 157388 279924 157452
rect 279988 157450 279994 157452
rect 282126 157450 282132 157452
rect 279988 157390 282132 157450
rect 279988 157388 279994 157390
rect 282126 157388 282132 157390
rect 282196 157388 282202 157452
rect 299054 157388 299060 157452
rect 299124 157450 299130 157452
rect 299124 157390 299674 157450
rect 299124 157388 299130 157390
rect 299614 157042 299674 157390
rect 300158 157388 300164 157452
rect 300228 157450 300234 157452
rect 303654 157450 303660 157452
rect 300228 157390 303660 157450
rect 300228 157388 300234 157390
rect 303654 157388 303660 157390
rect 303724 157388 303730 157452
rect 302734 157116 302740 157180
rect 302804 157178 302810 157180
rect 306414 157178 306420 157180
rect 302804 157118 306420 157178
rect 302804 157116 302810 157118
rect 306414 157116 306420 157118
rect 306484 157116 306490 157180
rect 299614 156982 306390 157042
rect 302601 156906 302667 156909
rect 305678 156906 305684 156908
rect 302601 156904 305684 156906
rect 302601 156848 302606 156904
rect 302662 156848 305684 156904
rect 302601 156846 305684 156848
rect 302601 156843 302667 156846
rect 305678 156844 305684 156846
rect 305748 156844 305754 156908
rect 248086 156708 248092 156772
rect 248156 156770 248162 156772
rect 264094 156770 264100 156772
rect 248156 156710 264100 156770
rect 248156 156708 248162 156710
rect 264094 156708 264100 156710
rect 264164 156708 264170 156772
rect 306330 156770 306390 156982
rect 311934 156770 311940 156772
rect 306330 156710 311940 156770
rect 311934 156708 311940 156710
rect 312004 156708 312010 156772
rect 4102 156572 4108 156636
rect 4172 156634 4178 156636
rect 272374 156634 272380 156636
rect 4172 156574 272380 156634
rect 4172 156572 4178 156574
rect 272374 156572 272380 156574
rect 272444 156572 272450 156636
rect 274398 156572 274404 156636
rect 274468 156634 274474 156636
rect 283414 156634 283420 156636
rect 274468 156574 283420 156634
rect 274468 156572 274474 156574
rect 283414 156572 283420 156574
rect 283484 156572 283490 156636
rect 285581 156634 285647 156637
rect 285581 156632 296730 156634
rect 285581 156576 285586 156632
rect 285642 156576 296730 156632
rect 285581 156574 296730 156576
rect 285581 156571 285647 156574
rect 296670 156498 296730 156574
rect 300526 156572 300532 156636
rect 300596 156634 300602 156636
rect 303838 156634 303844 156636
rect 300596 156574 303844 156634
rect 300596 156572 300602 156574
rect 303838 156572 303844 156574
rect 303908 156572 303914 156636
rect 307886 156572 307892 156636
rect 307956 156634 307962 156636
rect 578734 156634 578740 156636
rect 307956 156574 578740 156634
rect 307956 156572 307962 156574
rect 578734 156572 578740 156574
rect 578804 156572 578810 156636
rect 304993 156498 305059 156501
rect 296670 156496 305059 156498
rect 296670 156440 304998 156496
rect 305054 156440 305059 156496
rect 296670 156438 305059 156440
rect 304993 156435 305059 156438
rect 3550 155212 3556 155276
rect 3620 155274 3626 155276
rect 269614 155274 269620 155276
rect 3620 155214 269620 155274
rect 3620 155212 3626 155214
rect 269614 155212 269620 155214
rect 269684 155212 269690 155276
rect 311014 155212 311020 155276
rect 311084 155274 311090 155276
rect 580206 155274 580212 155276
rect 311084 155214 580212 155274
rect 311084 155212 311090 155214
rect 580206 155212 580212 155214
rect 580276 155212 580282 155276
rect 4654 153716 4660 153780
rect 4724 153778 4730 153780
rect 278998 153778 279004 153780
rect 4724 153718 279004 153778
rect 4724 153716 4730 153718
rect 278998 153716 279004 153718
rect 279068 153716 279074 153780
rect 309358 153716 309364 153780
rect 309428 153778 309434 153780
rect 577630 153778 577636 153780
rect 309428 153718 577636 153778
rect 309428 153716 309434 153718
rect 577630 153716 577636 153718
rect 577700 153716 577706 153780
rect 580901 152690 580967 152693
rect 583520 152690 584960 152780
rect 580901 152688 584960 152690
rect 580901 152632 580906 152688
rect 580962 152632 584960 152688
rect 580901 152630 584960 152632
rect 580901 152627 580967 152630
rect 583520 152540 584960 152630
rect 6126 152356 6132 152420
rect 6196 152418 6202 152420
rect 274582 152418 274588 152420
rect 6196 152358 274588 152418
rect 6196 152356 6202 152358
rect 274582 152356 274588 152358
rect 274652 152356 274658 152420
rect 7414 150996 7420 151060
rect 7484 151058 7490 151060
rect 277526 151058 277532 151060
rect 7484 150998 277532 151058
rect 7484 150996 7490 150998
rect 277526 150996 277532 150998
rect 277596 150996 277602 151060
rect -960 149834 480 149924
rect 2814 149834 2820 149836
rect -960 149774 2820 149834
rect -960 149684 480 149774
rect 2814 149772 2820 149774
rect 2884 149772 2890 149836
rect 3366 149636 3372 149700
rect 3436 149698 3442 149700
rect 271086 149698 271092 149700
rect 3436 149638 271092 149698
rect 3436 149636 3442 149638
rect 271086 149636 271092 149638
rect 271156 149636 271162 149700
rect 11697 148338 11763 148341
rect 262857 148338 262923 148341
rect 11697 148336 262923 148338
rect 11697 148280 11702 148336
rect 11758 148280 262862 148336
rect 262918 148280 262923 148336
rect 11697 148278 262923 148280
rect 11697 148275 11763 148278
rect 262857 148275 262923 148278
rect 580901 139362 580967 139365
rect 583520 139362 584960 139452
rect 580901 139360 584960 139362
rect 580901 139304 580906 139360
rect 580962 139304 584960 139360
rect 580901 139302 584960 139304
rect 580901 139299 580967 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 2773 136778 2839 136781
rect -960 136776 2839 136778
rect -960 136720 2778 136776
rect 2834 136720 2839 136776
rect -960 136718 2839 136720
rect -960 136628 480 136718
rect 2773 136715 2839 136718
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 580901 112842 580967 112845
rect 583520 112842 584960 112932
rect 580901 112840 584960 112842
rect 580901 112784 580906 112840
rect 580962 112784 584960 112840
rect 580901 112782 584960 112784
rect 580901 112779 580967 112782
rect 583520 112692 584960 112782
rect -960 110516 480 110756
rect 580901 99514 580967 99517
rect 583520 99514 584960 99604
rect 580901 99512 584960 99514
rect 580901 99456 580906 99512
rect 580962 99456 584960 99512
rect 580901 99454 584960 99456
rect 580901 99451 580967 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 2814 97610 2820 97612
rect -960 97550 2820 97610
rect -960 97460 480 97550
rect 2814 97548 2820 97550
rect 2884 97548 2890 97612
rect 4838 87484 4844 87548
rect 4908 87546 4914 87548
rect 276790 87546 276796 87548
rect 4908 87486 276796 87546
rect 4908 87484 4914 87486
rect 276790 87484 276796 87486
rect 276860 87484 276866 87548
rect 583520 86036 584960 86276
rect -960 84690 480 84780
rect 2814 84690 2820 84692
rect -960 84630 2820 84690
rect -960 84540 480 84630
rect 2814 84628 2820 84630
rect 2884 84628 2890 84692
rect 974 76468 980 76532
rect 1044 76530 1050 76532
rect 280286 76530 280292 76532
rect 1044 76470 280292 76530
rect 1044 76468 1050 76470
rect 280286 76468 280292 76470
rect 280356 76468 280362 76532
rect 308990 75108 308996 75172
rect 309060 75170 309066 75172
rect 577446 75170 577452 75172
rect 309060 75110 577452 75170
rect 309060 75108 309066 75110
rect 577446 75108 577452 75110
rect 577516 75108 577522 75172
rect 301814 74700 301820 74764
rect 301884 74762 301890 74764
rect 307702 74762 307708 74764
rect 301884 74702 307708 74762
rect 301884 74700 301890 74702
rect 307702 74700 307708 74702
rect 307772 74700 307778 74764
rect 300710 74564 300716 74628
rect 300780 74626 300786 74628
rect 306414 74626 306420 74628
rect 300780 74566 306420 74626
rect 300780 74564 300786 74566
rect 306414 74564 306420 74566
rect 306484 74564 306490 74628
rect 9070 73884 9076 73948
rect 9140 73946 9146 73948
rect 274214 73946 274220 73948
rect 9140 73886 274220 73946
rect 9140 73884 9146 73886
rect 274214 73884 274220 73886
rect 274284 73884 274290 73948
rect 2630 73748 2636 73812
rect 2700 73810 2706 73812
rect 278262 73810 278268 73812
rect 2700 73750 278268 73810
rect 2700 73748 2706 73750
rect 278262 73748 278268 73750
rect 278332 73748 278338 73812
rect 307150 73748 307156 73812
rect 307220 73810 307226 73812
rect 574686 73810 574692 73812
rect 307220 73750 574692 73810
rect 307220 73748 307226 73750
rect 574686 73748 574692 73750
rect 574756 73748 574762 73812
rect 580901 72994 580967 72997
rect 583520 72994 584960 73084
rect 580901 72992 584960 72994
rect 580901 72936 580906 72992
rect 580962 72936 584960 72992
rect 580901 72934 584960 72936
rect 580901 72931 580967 72934
rect 583520 72844 584960 72934
rect 304901 72450 304967 72453
rect 306373 72450 306439 72453
rect 304901 72448 306439 72450
rect 304901 72392 304906 72448
rect 304962 72392 306378 72448
rect 306434 72392 306439 72448
rect 304901 72390 306439 72392
rect 304901 72387 304967 72390
rect 306373 72387 306439 72390
rect 307518 72388 307524 72452
rect 307588 72450 307594 72452
rect 575974 72450 575980 72452
rect 307588 72390 575980 72450
rect 307588 72388 307594 72390
rect 575974 72388 575980 72390
rect 576044 72388 576050 72452
rect -960 71634 480 71724
rect 3366 71634 3372 71636
rect -960 71574 3372 71634
rect -960 71484 480 71574
rect 3366 71572 3372 71574
rect 3436 71572 3442 71636
rect 264094 71300 264100 71364
rect 264164 71362 264170 71364
rect 272558 71362 272564 71364
rect 264164 71302 272564 71362
rect 264164 71300 264170 71302
rect 272558 71300 272564 71302
rect 272628 71300 272634 71364
rect 43294 71164 43300 71228
rect 43364 71226 43370 71228
rect 276054 71226 276060 71228
rect 43364 71166 276060 71226
rect 43364 71164 43370 71166
rect 276054 71164 276060 71166
rect 276124 71164 276130 71228
rect 5390 71028 5396 71092
rect 5460 71090 5466 71092
rect 274950 71090 274956 71092
rect 5460 71030 274956 71090
rect 5460 71028 5466 71030
rect 274950 71028 274956 71030
rect 275020 71028 275026 71092
rect 277158 71028 277164 71092
rect 277228 71090 277234 71092
rect 281942 71090 281948 71092
rect 277228 71030 281948 71090
rect 277228 71028 277234 71030
rect 281942 71028 281948 71030
rect 282012 71028 282018 71092
rect 308254 71028 308260 71092
rect 308324 71090 308330 71092
rect 574870 71090 574876 71092
rect 308324 71030 574876 71090
rect 308324 71028 308330 71030
rect 574870 71028 574876 71030
rect 574940 71028 574946 71092
rect 262857 70818 262923 70821
rect 265065 70818 265131 70821
rect 262857 70816 265131 70818
rect 262857 70760 262862 70816
rect 262918 70760 265070 70816
rect 265126 70760 265131 70816
rect 262857 70758 265131 70760
rect 262857 70755 262923 70758
rect 265065 70755 265131 70758
rect 274398 69668 274404 69732
rect 274468 69730 274474 69732
rect 283414 69730 283420 69732
rect 274468 69670 283420 69730
rect 274468 69668 274474 69670
rect 283414 69668 283420 69670
rect 283484 69668 283490 69732
rect 8886 69532 8892 69596
rect 8956 69594 8962 69596
rect 278630 69594 278636 69596
rect 8956 69534 278636 69594
rect 8956 69532 8962 69534
rect 278630 69532 278636 69534
rect 278700 69532 278706 69596
rect 282821 69594 282887 69597
rect 306230 69594 306236 69596
rect 282821 69592 306236 69594
rect 282821 69536 282826 69592
rect 282882 69536 306236 69592
rect 282821 69534 306236 69536
rect 282821 69531 282887 69534
rect 306230 69532 306236 69534
rect 306300 69532 306306 69596
rect 308622 69532 308628 69596
rect 308692 69594 308698 69596
rect 578918 69594 578924 69596
rect 308692 69534 578924 69594
rect 308692 69532 308698 69534
rect 578918 69532 578924 69534
rect 578988 69532 578994 69596
rect 279918 68852 279924 68916
rect 279988 68914 279994 68916
rect 284150 68914 284156 68916
rect 279988 68854 284156 68914
rect 279988 68852 279994 68854
rect 284150 68852 284156 68854
rect 284220 68852 284226 68916
rect 293217 68914 293283 68917
rect 293350 68914 293356 68916
rect 293217 68912 293356 68914
rect 293217 68856 293222 68912
rect 293278 68856 293356 68912
rect 293217 68854 293356 68856
rect 293217 68851 293283 68854
rect 293350 68852 293356 68854
rect 293420 68852 293426 68916
rect 300853 68914 300919 68917
rect 301078 68914 301084 68916
rect 300853 68912 301084 68914
rect 300853 68856 300858 68912
rect 300914 68856 301084 68912
rect 300853 68854 301084 68856
rect 300853 68851 300919 68854
rect 301078 68852 301084 68854
rect 301148 68852 301154 68916
rect 301446 68852 301452 68916
rect 301516 68914 301522 68916
rect 304206 68914 304212 68916
rect 301516 68854 304212 68914
rect 301516 68852 301522 68854
rect 304206 68852 304212 68854
rect 304276 68852 304282 68916
rect 304993 68914 305059 68917
rect 305310 68914 305316 68916
rect 304993 68912 305316 68914
rect 304993 68856 304998 68912
rect 305054 68856 305316 68912
rect 304993 68854 305316 68856
rect 304993 68851 305059 68854
rect 305310 68852 305316 68854
rect 305380 68852 305386 68916
rect 300342 68716 300348 68780
rect 300412 68778 300418 68780
rect 303838 68778 303844 68780
rect 300412 68718 303844 68778
rect 300412 68716 300418 68718
rect 303838 68716 303844 68718
rect 303908 68716 303914 68780
rect 272558 68580 272564 68644
rect 272628 68642 272634 68644
rect 282678 68642 282684 68644
rect 272628 68582 282684 68642
rect 272628 68580 272634 68582
rect 282678 68580 282684 68582
rect 282748 68580 282754 68644
rect 298502 68580 298508 68644
rect 298572 68642 298578 68644
rect 311934 68642 311940 68644
rect 298572 68582 311940 68642
rect 298572 68580 298578 68582
rect 311934 68580 311940 68582
rect 312004 68580 312010 68644
rect 9857 68506 9923 68509
rect 279734 68506 279740 68508
rect 9857 68504 279740 68506
rect 9857 68448 9862 68504
rect 9918 68448 279740 68504
rect 9857 68446 279740 68448
rect 9857 68443 9923 68446
rect 279734 68444 279740 68446
rect 279804 68444 279810 68508
rect 304574 68444 304580 68508
rect 304644 68506 304650 68508
rect 335353 68506 335419 68509
rect 304644 68504 335419 68506
rect 304644 68448 335358 68504
rect 335414 68448 335419 68504
rect 304644 68446 335419 68448
rect 304644 68444 304650 68446
rect 335353 68443 335419 68446
rect 1894 68308 1900 68372
rect 1964 68370 1970 68372
rect 275318 68370 275324 68372
rect 1964 68310 275324 68370
rect 1964 68308 1970 68310
rect 275318 68308 275324 68310
rect 275388 68308 275394 68372
rect 302550 68308 302556 68372
rect 302620 68370 302626 68372
rect 334750 68370 334756 68372
rect 302620 68310 334756 68370
rect 302620 68308 302626 68310
rect 334750 68308 334756 68310
rect 334820 68308 334826 68372
rect 1158 68172 1164 68236
rect 1228 68234 1234 68236
rect 276422 68234 276428 68236
rect 1228 68174 276428 68234
rect 1228 68172 1234 68174
rect 276422 68172 276428 68174
rect 276492 68172 276498 68236
rect 277894 68172 277900 68236
rect 277964 68234 277970 68236
rect 303654 68234 303660 68236
rect 277964 68174 303660 68234
rect 277964 68172 277970 68174
rect 303654 68172 303660 68174
rect 303724 68172 303730 68236
rect 306782 68172 306788 68236
rect 306852 68234 306858 68236
rect 582373 68234 582439 68237
rect 306852 68232 582439 68234
rect 306852 68176 582378 68232
rect 582434 68176 582439 68232
rect 306852 68174 582439 68176
rect 306852 68172 306858 68174
rect 582373 68171 582439 68174
rect 282177 67690 282243 67693
rect 282310 67690 282316 67692
rect 282177 67688 282316 67690
rect 282177 67632 282182 67688
rect 282238 67632 282316 67688
rect 282177 67630 282316 67632
rect 282177 67627 282243 67630
rect 282310 67628 282316 67630
rect 282380 67628 282386 67692
rect 279366 67492 279372 67556
rect 279436 67554 279442 67556
rect 280797 67554 280863 67557
rect 279436 67552 280863 67554
rect 279436 67496 280802 67552
rect 280858 67496 280863 67552
rect 279436 67494 280863 67496
rect 279436 67492 279442 67494
rect 280797 67491 280863 67494
rect 283046 67492 283052 67556
rect 283116 67554 283122 67556
rect 283557 67554 283623 67557
rect 283116 67552 283623 67554
rect 283116 67496 283562 67552
rect 283618 67496 283623 67552
rect 283116 67494 283623 67496
rect 283116 67492 283122 67494
rect 283557 67491 283623 67494
rect 304901 67554 304967 67557
rect 306046 67554 306052 67556
rect 304901 67552 306052 67554
rect 304901 67496 304906 67552
rect 304962 67496 306052 67552
rect 304901 67494 306052 67496
rect 304901 67491 304967 67494
rect 306046 67492 306052 67494
rect 306116 67492 306122 67556
rect 265065 67146 265131 67149
rect 303838 67146 303844 67148
rect 265065 67144 303844 67146
rect 265065 67088 265070 67144
rect 265126 67088 303844 67144
rect 265065 67086 303844 67088
rect 265065 67083 265131 67086
rect 303838 67084 303844 67086
rect 303908 67084 303914 67148
rect 111006 66948 111012 67012
rect 111076 67010 111082 67012
rect 277158 67010 277164 67012
rect 111076 66950 277164 67010
rect 111076 66948 111082 66950
rect 277158 66948 277164 66950
rect 277228 66948 277234 67012
rect 290958 66948 290964 67012
rect 291028 67010 291034 67012
rect 301446 67010 301452 67012
rect 291028 66950 301452 67010
rect 291028 66948 291034 66950
rect 301446 66948 301452 66950
rect 301516 66948 301522 67012
rect 6678 66812 6684 66876
rect 6748 66874 6754 66876
rect 275686 66874 275692 66876
rect 6748 66814 275692 66874
rect 6748 66812 6754 66814
rect 275686 66812 275692 66814
rect 275756 66812 275762 66876
rect 290457 66874 290523 66877
rect 304942 66874 304948 66876
rect 290457 66872 304948 66874
rect 290457 66816 290462 66872
rect 290518 66816 304948 66872
rect 290457 66814 304948 66816
rect 290457 66811 290523 66814
rect 304942 66812 304948 66814
rect 305012 66812 305018 66876
rect 580901 59666 580967 59669
rect 583520 59666 584960 59756
rect 580901 59664 584960 59666
rect 580901 59608 580906 59664
rect 580962 59608 584960 59664
rect 580901 59606 584960 59608
rect 580901 59603 580967 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 2814 58578 2820 58580
rect -960 58518 2820 58578
rect -960 58428 480 58518
rect 2814 58516 2820 58518
rect 2884 58516 2890 58580
rect 583520 46188 584960 46428
rect -960 45522 480 45612
rect 2773 45522 2839 45525
rect -960 45520 2839 45522
rect -960 45464 2778 45520
rect 2834 45464 2839 45520
rect -960 45462 2839 45464
rect -960 45372 480 45462
rect 2773 45459 2839 45462
rect 2773 44298 2839 44301
rect 3417 44298 3483 44301
rect 2773 44296 3483 44298
rect 2773 44240 2778 44296
rect 2834 44240 3422 44296
rect 3478 44240 3483 44296
rect 2773 44238 3483 44240
rect 2773 44235 2839 44238
rect 3417 44235 3483 44238
rect 580901 33146 580967 33149
rect 583520 33146 584960 33236
rect 580901 33144 584960 33146
rect 580901 33088 580906 33144
rect 580962 33088 584960 33144
rect 580901 33086 584960 33088
rect 580901 33083 580967 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 3417 24170 3483 24173
rect 273253 24170 273319 24173
rect 3417 24168 273319 24170
rect 3417 24112 3422 24168
rect 3478 24112 273258 24168
rect 273314 24112 273319 24168
rect 3417 24110 273319 24112
rect 3417 24107 3483 24110
rect 273253 24107 273319 24110
rect 3366 22612 3372 22676
rect 3436 22674 3442 22676
rect 273294 22674 273300 22676
rect 3436 22614 273300 22674
rect 3436 22612 3442 22614
rect 273294 22612 273300 22614
rect 273364 22612 273370 22676
rect 269614 21932 269620 21996
rect 269684 21994 269690 21996
rect 276238 21994 276244 21996
rect 269684 21934 276244 21994
rect 269684 21932 269690 21934
rect 276238 21932 276244 21934
rect 276308 21932 276314 21996
rect 306414 21932 306420 21996
rect 306484 21994 306490 21996
rect 576158 21994 576164 21996
rect 306484 21934 576164 21994
rect 306484 21932 306490 21934
rect 576158 21932 576164 21934
rect 576228 21932 576234 21996
rect 8150 21796 8156 21860
rect 8220 21858 8226 21860
rect 275502 21858 275508 21860
rect 8220 21798 275508 21858
rect 8220 21796 8226 21798
rect 275502 21796 275508 21798
rect 275572 21796 275578 21860
rect 6310 21660 6316 21724
rect 6380 21722 6386 21724
rect 276606 21722 276612 21724
rect 6380 21662 276612 21722
rect 6380 21660 6386 21662
rect 276606 21660 276612 21662
rect 276676 21660 276682 21724
rect 2814 20572 2820 20636
rect 2884 20634 2890 20636
rect 2884 20574 6930 20634
rect 2884 20572 2890 20574
rect 6870 20498 6930 20574
rect 273294 20572 273300 20636
rect 273364 20634 273370 20636
rect 278262 20634 278268 20636
rect 273364 20574 278268 20634
rect 273364 20572 273370 20574
rect 278262 20572 278268 20574
rect 278332 20572 278338 20636
rect 306598 20572 306604 20636
rect 306668 20634 306674 20636
rect 311014 20634 311020 20636
rect 306668 20574 311020 20634
rect 306668 20572 306674 20574
rect 311014 20572 311020 20574
rect 311084 20572 311090 20636
rect 277894 20498 277900 20500
rect 6870 20438 277900 20498
rect 277894 20436 277900 20438
rect 277964 20498 277970 20500
rect 573357 20498 573423 20501
rect 277964 20496 573423 20498
rect 277964 20440 573362 20496
rect 573418 20440 573423 20496
rect 277964 20438 573423 20440
rect 277964 20436 277970 20438
rect 573357 20435 573423 20438
rect 2078 20300 2084 20364
rect 2148 20362 2154 20364
rect 277158 20362 277164 20364
rect 2148 20302 277164 20362
rect 2148 20300 2154 20302
rect 277158 20300 277164 20302
rect 277228 20300 277234 20364
rect 273253 20226 273319 20229
rect 277526 20226 277532 20228
rect 273253 20224 277532 20226
rect 273253 20168 273258 20224
rect 273314 20168 277532 20224
rect 273253 20166 277532 20168
rect 273253 20163 273319 20166
rect 277526 20164 277532 20166
rect 277596 20226 277602 20228
rect 278681 20226 278747 20229
rect 277596 20224 278747 20226
rect 277596 20168 278686 20224
rect 278742 20168 278747 20224
rect 277596 20166 278747 20168
rect 277596 20164 277602 20166
rect 278681 20163 278747 20166
rect 54 20028 60 20092
rect 124 20090 130 20092
rect 275318 20090 275324 20092
rect 124 20030 275324 20090
rect 124 20028 130 20030
rect 275318 20028 275324 20030
rect 275388 20028 275394 20092
rect 580901 19818 580967 19821
rect 583520 19818 584960 19908
rect 576810 19816 584960 19818
rect 576810 19760 580906 19816
rect 580962 19760 584960 19816
rect 576810 19758 584960 19760
rect 2773 19548 2839 19549
rect 2773 19546 2820 19548
rect 2638 19544 2820 19546
rect -960 19410 480 19500
rect 2638 19488 2778 19544
rect 2638 19486 2820 19488
rect 2638 19410 2698 19486
rect 2773 19484 2820 19486
rect 2884 19484 2890 19548
rect 277301 19546 277367 19549
rect 277301 19544 277410 19546
rect 277301 19488 277306 19544
rect 277362 19488 277410 19544
rect 2773 19483 2839 19484
rect 277301 19483 277410 19488
rect -960 19350 2698 19410
rect -960 19260 480 19350
rect 7598 19212 7604 19276
rect 7668 19274 7674 19276
rect 276422 19274 276428 19276
rect 7668 19214 276428 19274
rect 7668 19212 7674 19214
rect 276422 19212 276428 19214
rect 276492 19212 276498 19276
rect 277350 19274 277410 19483
rect 278681 19410 278747 19413
rect 576810 19410 576870 19758
rect 580901 19755 580967 19758
rect 583520 19668 584960 19758
rect 278681 19408 279250 19410
rect 278681 19352 278686 19408
rect 278742 19352 279250 19408
rect 278681 19350 279250 19352
rect 278681 19347 278747 19350
rect 278998 19274 279004 19276
rect 277350 19214 279004 19274
rect 278998 19212 279004 19214
rect 279068 19212 279074 19276
rect 279190 19274 279250 19350
rect 572670 19350 576870 19410
rect 572670 19274 572730 19350
rect 279190 19214 572730 19274
rect 272374 19076 272380 19140
rect 272444 19138 272450 19140
rect 278630 19138 278636 19140
rect 272444 19078 278636 19138
rect 272444 19076 272450 19078
rect 278630 19076 278636 19078
rect 278700 19076 278706 19140
rect 271086 18940 271092 19004
rect 271156 19002 271162 19004
rect 277301 19002 277367 19005
rect 271156 19000 277367 19002
rect 271156 18944 277306 19000
rect 277362 18944 277367 19000
rect 271156 18942 277367 18944
rect 271156 18940 271162 18942
rect 277301 18939 277367 18942
rect -960 6490 480 6580
rect 2773 6490 2839 6493
rect -960 6488 2839 6490
rect -960 6432 2778 6488
rect 2834 6432 2839 6488
rect 583520 6476 584960 6716
rect -960 6430 2839 6432
rect -960 6340 480 6430
rect 2773 6427 2839 6430
rect 579797 3498 579863 3501
rect 580758 3498 580764 3500
rect 579797 3496 580764 3498
rect 579797 3440 579802 3496
rect 579858 3440 580764 3496
rect 579797 3438 580764 3440
rect 579797 3435 579863 3438
rect 580758 3436 580764 3438
rect 580828 3436 580834 3500
<< via3 >>
rect 284340 699756 284404 699820
rect 9812 684252 9876 684316
rect 3372 671196 3436 671260
rect 574692 670652 574756 670716
rect 291148 658140 291212 658204
rect 8892 632028 8956 632092
rect 4660 619108 4724 619172
rect 575980 617476 576044 617540
rect 288388 606052 288452 606116
rect 7420 579940 7484 580004
rect 282132 566884 282196 566948
rect 578740 564300 578804 564364
rect 17908 553828 17972 553892
rect 2820 527852 2884 527916
rect 4844 514796 4908 514860
rect 574876 511260 574940 511324
rect 12388 501740 12452 501804
rect 1900 475628 1964 475692
rect 13860 462572 13924 462636
rect 578924 458084 578988 458148
rect 11100 449516 11164 449580
rect 9076 423540 9140 423604
rect 6132 410484 6196 410548
rect 577452 404908 577516 404972
rect 15148 397428 15212 397492
rect 60 371588 124 371652
rect 9812 358396 9876 358460
rect 577636 351868 577700 351932
rect 3556 345340 3620 345404
rect 7604 319228 7668 319292
rect 3372 306988 3436 307052
rect 16620 306988 16684 307052
rect 3740 306172 3804 306236
rect 580212 298692 580276 298756
rect 2084 293116 2148 293180
rect 3372 267140 3436 267204
rect 3740 256668 3804 256732
rect 6316 256668 6380 256732
rect 3004 254220 3068 254284
rect 576164 245516 576228 245580
rect 1164 242796 1228 242860
rect 2820 242796 2884 242860
rect 580580 232324 580644 232388
rect 580764 218996 580828 219060
rect 285628 214508 285692 214572
rect 10180 213828 10244 213892
rect 12388 213828 12452 213892
rect 9444 213692 9508 213756
rect 11100 213692 11164 213756
rect 6684 213556 6748 213620
rect 13860 213556 13924 213620
rect 5396 213420 5460 213484
rect 15148 213420 15212 213484
rect 2636 213284 2700 213348
rect 17908 213284 17972 213348
rect 980 213148 1044 213212
rect 16620 213148 16684 213212
rect 288204 210292 288268 210356
rect 3004 201860 3068 201924
rect 8156 196012 8220 196076
rect 9812 196012 9876 196076
rect 7972 194516 8036 194580
rect 10180 194516 10244 194580
rect 289676 192476 289740 192540
rect 580580 192476 580644 192540
rect 282868 192204 282932 192268
rect 298140 192204 298204 192268
rect 284524 192068 284588 192132
rect 281028 191932 281092 191996
rect 295196 191932 295260 191996
rect 297956 191796 298020 191860
rect 282132 191524 282196 191588
rect 286180 191524 286244 191588
rect 295196 190844 295260 190908
rect 283972 190572 284036 190636
rect 296300 190572 296364 190636
rect 285444 190300 285508 190364
rect 300900 190436 300964 190500
rect 282684 189620 282748 189684
rect 283788 189484 283852 189548
rect 297036 189484 297100 189548
rect 288020 189348 288084 189412
rect 298692 189348 298756 189412
rect 284156 189212 284220 189276
rect 298140 189212 298204 189276
rect 301452 189212 301516 189276
rect 9628 189076 9692 189140
rect 289860 189076 289924 189140
rect 299428 189076 299492 189140
rect 301268 189076 301332 189140
rect 2820 188804 2884 188868
rect 290964 188396 291028 188460
rect 299612 188396 299676 188460
rect 282316 188260 282380 188324
rect 293172 188260 293236 188324
rect 301084 188260 301148 188324
rect 293540 188124 293604 188188
rect 299060 187988 299124 188052
rect 292436 187852 292500 187916
rect 290964 187716 291028 187780
rect 295012 187716 295076 187780
rect 299244 187716 299308 187780
rect 299612 187716 299676 187780
rect 299428 187580 299492 187644
rect 285444 187444 285508 187508
rect 300900 187444 300964 187508
rect 282500 187308 282564 187372
rect 285628 187308 285692 187372
rect 300900 187308 300964 187372
rect 301452 187308 301516 187372
rect 299980 187172 300044 187236
rect 299244 186900 299308 186964
rect 298876 186764 298940 186828
rect 282316 186628 282380 186692
rect 286364 186628 286428 186692
rect 299612 186628 299676 186692
rect 301268 186628 301332 186692
rect 288020 186492 288084 186556
rect 298140 186492 298204 186556
rect 298692 186492 298756 186556
rect 297404 186356 297468 186420
rect 297956 186356 298020 186420
rect 283788 186084 283852 186148
rect 293908 186084 293972 186148
rect 297036 186084 297100 186148
rect 284156 185948 284220 186012
rect 295196 185948 295260 186012
rect 296484 185948 296548 186012
rect 283972 185812 284036 185876
rect 296300 185812 296364 185876
rect 282868 185676 282932 185740
rect 291332 185676 291396 185740
rect 295012 185676 295076 185740
rect 295932 185540 295996 185604
rect 299796 185736 299860 185740
rect 299796 185680 299810 185736
rect 299810 185680 299860 185736
rect 299796 185676 299860 185680
rect 295564 185404 295628 185468
rect 299428 185404 299492 185468
rect 294828 185268 294892 185332
rect 294460 185132 294524 185196
rect 285444 184860 285508 184924
rect 286548 184860 286612 184924
rect 291148 184860 291212 184924
rect 293908 184996 293972 185060
rect 293724 184860 293788 184924
rect 282684 184724 282748 184788
rect 293172 184784 293236 184788
rect 293172 184728 293222 184784
rect 293222 184728 293236 184784
rect 293172 184724 293236 184728
rect 301084 184724 301148 184788
rect 292988 184588 293052 184652
rect 282868 184452 282932 184516
rect 291332 184452 291396 184516
rect 292620 184452 292684 184516
rect 284524 184316 284588 184380
rect 291884 184180 291948 184244
rect 291516 184044 291580 184108
rect 290412 183908 290476 183972
rect 290044 183772 290108 183836
rect 281028 183636 281092 183700
rect 284340 183636 284404 183700
rect 288388 183560 288452 183564
rect 288388 183504 288438 183560
rect 288438 183504 288452 183560
rect 288388 183500 288452 183504
rect 292252 183636 292316 183700
rect 289308 183500 289372 183564
rect 288940 183364 289004 183428
rect 288572 183228 288636 183292
rect 288020 183092 288084 183156
rect 287836 182956 287900 183020
rect 287468 182820 287532 182884
rect 287100 182684 287164 182748
rect 288204 182548 288268 182612
rect 301268 182548 301332 182612
rect 286364 182412 286428 182476
rect 299612 182412 299676 182476
rect 285996 182276 286060 182340
rect 285260 182004 285324 182068
rect 284892 181868 284956 181932
rect 284524 181732 284588 181796
rect 283052 181596 283116 181660
rect 284340 181460 284404 181524
rect 283420 181324 283484 181388
rect 300900 181324 300964 181388
rect 281580 181052 281644 181116
rect 281948 180780 282012 180844
rect 296852 180780 296916 180844
rect 282500 180644 282564 180708
rect 282868 180508 282932 180572
rect 283420 180372 283484 180436
rect 300900 180372 300964 180436
rect 285628 180100 285692 180164
rect 296116 180100 296180 180164
rect 296484 180100 296548 180164
rect 286548 179964 286612 180028
rect 302372 179964 302436 180028
rect 293540 179828 293604 179892
rect 300532 179828 300596 179892
rect 289860 179480 289924 179484
rect 289860 179424 289910 179480
rect 289910 179424 289924 179480
rect 289860 179420 289924 179424
rect 292436 179420 292500 179484
rect 299060 179420 299124 179484
rect 302372 179420 302436 179484
rect 301636 179284 301700 179348
rect 580580 179148 580644 179212
rect 9444 178876 9508 178940
rect 43300 178876 43364 178940
rect 286180 178876 286244 178940
rect 7972 178740 8036 178804
rect 111012 178740 111076 178804
rect 300164 178740 300228 178804
rect 300532 178740 300596 178804
rect 334756 178740 334820 178804
rect 248092 178604 248156 178668
rect 281580 178604 281644 178668
rect 289676 178060 289740 178124
rect 281212 177924 281276 177988
rect 282868 177924 282932 177988
rect 289676 177924 289740 177988
rect 296116 177924 296180 177988
rect 286732 177380 286796 177444
rect 301268 177380 301332 177444
rect 301452 177244 301516 177308
rect 299060 176700 299124 176764
rect 301084 176700 301148 176764
rect 282132 175884 282196 175948
rect 283052 175884 283116 175948
rect 10180 175204 10244 175268
rect 303108 174524 303172 174588
rect 580580 174524 580644 174588
rect 4108 162828 4172 162892
rect 301636 158068 301700 158132
rect 307708 158068 307772 158132
rect 277164 157932 277228 157996
rect 281764 157932 281828 157996
rect 10180 157388 10244 157452
rect 279924 157388 279988 157452
rect 282132 157388 282196 157452
rect 299060 157388 299124 157452
rect 300164 157388 300228 157452
rect 303660 157388 303724 157452
rect 302740 157116 302804 157180
rect 306420 157116 306484 157180
rect 305684 156844 305748 156908
rect 248092 156708 248156 156772
rect 264100 156708 264164 156772
rect 311940 156708 312004 156772
rect 4108 156572 4172 156636
rect 272380 156572 272444 156636
rect 274404 156572 274468 156636
rect 283420 156572 283484 156636
rect 300532 156572 300596 156636
rect 303844 156572 303908 156636
rect 307892 156572 307956 156636
rect 578740 156572 578804 156636
rect 3556 155212 3620 155276
rect 269620 155212 269684 155276
rect 311020 155212 311084 155276
rect 580212 155212 580276 155276
rect 4660 153716 4724 153780
rect 279004 153716 279068 153780
rect 309364 153716 309428 153780
rect 577636 153716 577700 153780
rect 6132 152356 6196 152420
rect 274588 152356 274652 152420
rect 7420 150996 7484 151060
rect 277532 150996 277596 151060
rect 2820 149772 2884 149836
rect 3372 149636 3436 149700
rect 271092 149636 271156 149700
rect 2820 97548 2884 97612
rect 4844 87484 4908 87548
rect 276796 87484 276860 87548
rect 2820 84628 2884 84692
rect 980 76468 1044 76532
rect 280292 76468 280356 76532
rect 308996 75108 309060 75172
rect 577452 75108 577516 75172
rect 301820 74700 301884 74764
rect 307708 74700 307772 74764
rect 300716 74564 300780 74628
rect 306420 74564 306484 74628
rect 9076 73884 9140 73948
rect 274220 73884 274284 73948
rect 2636 73748 2700 73812
rect 278268 73748 278332 73812
rect 307156 73748 307220 73812
rect 574692 73748 574756 73812
rect 307524 72388 307588 72452
rect 575980 72388 576044 72452
rect 3372 71572 3436 71636
rect 264100 71300 264164 71364
rect 272564 71300 272628 71364
rect 43300 71164 43364 71228
rect 276060 71164 276124 71228
rect 5396 71028 5460 71092
rect 274956 71028 275020 71092
rect 277164 71028 277228 71092
rect 281948 71028 282012 71092
rect 308260 71028 308324 71092
rect 574876 71028 574940 71092
rect 274404 69668 274468 69732
rect 283420 69668 283484 69732
rect 8892 69532 8956 69596
rect 278636 69532 278700 69596
rect 306236 69532 306300 69596
rect 308628 69532 308692 69596
rect 578924 69532 578988 69596
rect 279924 68852 279988 68916
rect 284156 68852 284220 68916
rect 293356 68852 293420 68916
rect 301084 68852 301148 68916
rect 301452 68852 301516 68916
rect 304212 68852 304276 68916
rect 305316 68852 305380 68916
rect 300348 68716 300412 68780
rect 303844 68716 303908 68780
rect 272564 68580 272628 68644
rect 282684 68580 282748 68644
rect 298508 68580 298572 68644
rect 311940 68580 312004 68644
rect 279740 68444 279804 68508
rect 304580 68444 304644 68508
rect 1900 68308 1964 68372
rect 275324 68308 275388 68372
rect 302556 68308 302620 68372
rect 334756 68308 334820 68372
rect 1164 68172 1228 68236
rect 276428 68172 276492 68236
rect 277900 68172 277964 68236
rect 303660 68172 303724 68236
rect 306788 68172 306852 68236
rect 282316 67628 282380 67692
rect 279372 67492 279436 67556
rect 283052 67492 283116 67556
rect 306052 67492 306116 67556
rect 303844 67084 303908 67148
rect 111012 66948 111076 67012
rect 277164 66948 277228 67012
rect 290964 66948 291028 67012
rect 301452 66948 301516 67012
rect 6684 66812 6748 66876
rect 275692 66812 275756 66876
rect 304948 66812 305012 66876
rect 2820 58516 2884 58580
rect 3372 22612 3436 22676
rect 273300 22612 273364 22676
rect 269620 21932 269684 21996
rect 276244 21932 276308 21996
rect 306420 21932 306484 21996
rect 576164 21932 576228 21996
rect 8156 21796 8220 21860
rect 275508 21796 275572 21860
rect 6316 21660 6380 21724
rect 276612 21660 276676 21724
rect 2820 20572 2884 20636
rect 273300 20572 273364 20636
rect 278268 20572 278332 20636
rect 306604 20572 306668 20636
rect 311020 20572 311084 20636
rect 277900 20436 277964 20500
rect 2084 20300 2148 20364
rect 277164 20300 277228 20364
rect 277532 20164 277596 20228
rect 60 20028 124 20092
rect 275324 20028 275388 20092
rect 2820 19544 2884 19548
rect 2820 19488 2834 19544
rect 2834 19488 2884 19544
rect 2820 19484 2884 19488
rect 7604 19212 7668 19276
rect 276428 19212 276492 19276
rect 279004 19212 279068 19276
rect 272380 19076 272444 19140
rect 278636 19076 278700 19140
rect 271092 18940 271156 19004
rect 580764 3436 580828 3500
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 -7066 -8106 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 -6106 -7146 710042
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 -5146 -6186 709082
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 -4186 -5226 708122
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 -3226 -4266 707162
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 -2266 -3306 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 694454 -2346 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 694218 -2934 694454
rect -2698 694218 -2614 694454
rect -2378 694218 -2346 694454
rect -2966 694134 -2346 694218
rect -2966 693898 -2934 694134
rect -2698 693898 -2614 694134
rect -2378 693898 -2346 694134
rect -2966 684454 -2346 693898
rect -2966 684218 -2934 684454
rect -2698 684218 -2614 684454
rect -2378 684218 -2346 684454
rect -2966 684134 -2346 684218
rect -2966 683898 -2934 684134
rect -2698 683898 -2614 684134
rect -2378 683898 -2346 684134
rect -2966 674454 -2346 683898
rect -2966 674218 -2934 674454
rect -2698 674218 -2614 674454
rect -2378 674218 -2346 674454
rect -2966 674134 -2346 674218
rect -2966 673898 -2934 674134
rect -2698 673898 -2614 674134
rect -2378 673898 -2346 674134
rect -2966 664454 -2346 673898
rect -2966 664218 -2934 664454
rect -2698 664218 -2614 664454
rect -2378 664218 -2346 664454
rect -2966 664134 -2346 664218
rect -2966 663898 -2934 664134
rect -2698 663898 -2614 664134
rect -2378 663898 -2346 664134
rect -2966 654454 -2346 663898
rect -2966 654218 -2934 654454
rect -2698 654218 -2614 654454
rect -2378 654218 -2346 654454
rect -2966 654134 -2346 654218
rect -2966 653898 -2934 654134
rect -2698 653898 -2614 654134
rect -2378 653898 -2346 654134
rect -2966 644454 -2346 653898
rect -2966 644218 -2934 644454
rect -2698 644218 -2614 644454
rect -2378 644218 -2346 644454
rect -2966 644134 -2346 644218
rect -2966 643898 -2934 644134
rect -2698 643898 -2614 644134
rect -2378 643898 -2346 644134
rect -2966 634454 -2346 643898
rect -2966 634218 -2934 634454
rect -2698 634218 -2614 634454
rect -2378 634218 -2346 634454
rect -2966 634134 -2346 634218
rect -2966 633898 -2934 634134
rect -2698 633898 -2614 634134
rect -2378 633898 -2346 634134
rect -2966 624454 -2346 633898
rect -2966 624218 -2934 624454
rect -2698 624218 -2614 624454
rect -2378 624218 -2346 624454
rect -2966 624134 -2346 624218
rect -2966 623898 -2934 624134
rect -2698 623898 -2614 624134
rect -2378 623898 -2346 624134
rect -2966 614454 -2346 623898
rect -2966 614218 -2934 614454
rect -2698 614218 -2614 614454
rect -2378 614218 -2346 614454
rect -2966 614134 -2346 614218
rect -2966 613898 -2934 614134
rect -2698 613898 -2614 614134
rect -2378 613898 -2346 614134
rect -2966 604454 -2346 613898
rect -2966 604218 -2934 604454
rect -2698 604218 -2614 604454
rect -2378 604218 -2346 604454
rect -2966 604134 -2346 604218
rect -2966 603898 -2934 604134
rect -2698 603898 -2614 604134
rect -2378 603898 -2346 604134
rect -2966 594454 -2346 603898
rect -2966 594218 -2934 594454
rect -2698 594218 -2614 594454
rect -2378 594218 -2346 594454
rect -2966 594134 -2346 594218
rect -2966 593898 -2934 594134
rect -2698 593898 -2614 594134
rect -2378 593898 -2346 594134
rect -2966 584454 -2346 593898
rect -2966 584218 -2934 584454
rect -2698 584218 -2614 584454
rect -2378 584218 -2346 584454
rect -2966 584134 -2346 584218
rect -2966 583898 -2934 584134
rect -2698 583898 -2614 584134
rect -2378 583898 -2346 584134
rect -2966 574454 -2346 583898
rect -2966 574218 -2934 574454
rect -2698 574218 -2614 574454
rect -2378 574218 -2346 574454
rect -2966 574134 -2346 574218
rect -2966 573898 -2934 574134
rect -2698 573898 -2614 574134
rect -2378 573898 -2346 574134
rect -2966 564454 -2346 573898
rect -2966 564218 -2934 564454
rect -2698 564218 -2614 564454
rect -2378 564218 -2346 564454
rect -2966 564134 -2346 564218
rect -2966 563898 -2934 564134
rect -2698 563898 -2614 564134
rect -2378 563898 -2346 564134
rect -2966 554454 -2346 563898
rect -2966 554218 -2934 554454
rect -2698 554218 -2614 554454
rect -2378 554218 -2346 554454
rect -2966 554134 -2346 554218
rect -2966 553898 -2934 554134
rect -2698 553898 -2614 554134
rect -2378 553898 -2346 554134
rect -2966 544454 -2346 553898
rect -2966 544218 -2934 544454
rect -2698 544218 -2614 544454
rect -2378 544218 -2346 544454
rect -2966 544134 -2346 544218
rect -2966 543898 -2934 544134
rect -2698 543898 -2614 544134
rect -2378 543898 -2346 544134
rect -2966 534454 -2346 543898
rect -2966 534218 -2934 534454
rect -2698 534218 -2614 534454
rect -2378 534218 -2346 534454
rect -2966 534134 -2346 534218
rect -2966 533898 -2934 534134
rect -2698 533898 -2614 534134
rect -2378 533898 -2346 534134
rect -2966 524454 -2346 533898
rect -2966 524218 -2934 524454
rect -2698 524218 -2614 524454
rect -2378 524218 -2346 524454
rect -2966 524134 -2346 524218
rect -2966 523898 -2934 524134
rect -2698 523898 -2614 524134
rect -2378 523898 -2346 524134
rect -2966 514454 -2346 523898
rect -2966 514218 -2934 514454
rect -2698 514218 -2614 514454
rect -2378 514218 -2346 514454
rect -2966 514134 -2346 514218
rect -2966 513898 -2934 514134
rect -2698 513898 -2614 514134
rect -2378 513898 -2346 514134
rect -2966 504454 -2346 513898
rect -2966 504218 -2934 504454
rect -2698 504218 -2614 504454
rect -2378 504218 -2346 504454
rect -2966 504134 -2346 504218
rect -2966 503898 -2934 504134
rect -2698 503898 -2614 504134
rect -2378 503898 -2346 504134
rect -2966 494454 -2346 503898
rect -2966 494218 -2934 494454
rect -2698 494218 -2614 494454
rect -2378 494218 -2346 494454
rect -2966 494134 -2346 494218
rect -2966 493898 -2934 494134
rect -2698 493898 -2614 494134
rect -2378 493898 -2346 494134
rect -2966 484454 -2346 493898
rect -2966 484218 -2934 484454
rect -2698 484218 -2614 484454
rect -2378 484218 -2346 484454
rect -2966 484134 -2346 484218
rect -2966 483898 -2934 484134
rect -2698 483898 -2614 484134
rect -2378 483898 -2346 484134
rect -2966 474454 -2346 483898
rect -2966 474218 -2934 474454
rect -2698 474218 -2614 474454
rect -2378 474218 -2346 474454
rect -2966 474134 -2346 474218
rect -2966 473898 -2934 474134
rect -2698 473898 -2614 474134
rect -2378 473898 -2346 474134
rect -2966 464454 -2346 473898
rect -2966 464218 -2934 464454
rect -2698 464218 -2614 464454
rect -2378 464218 -2346 464454
rect -2966 464134 -2346 464218
rect -2966 463898 -2934 464134
rect -2698 463898 -2614 464134
rect -2378 463898 -2346 464134
rect -2966 454454 -2346 463898
rect -2966 454218 -2934 454454
rect -2698 454218 -2614 454454
rect -2378 454218 -2346 454454
rect -2966 454134 -2346 454218
rect -2966 453898 -2934 454134
rect -2698 453898 -2614 454134
rect -2378 453898 -2346 454134
rect -2966 444454 -2346 453898
rect -2966 444218 -2934 444454
rect -2698 444218 -2614 444454
rect -2378 444218 -2346 444454
rect -2966 444134 -2346 444218
rect -2966 443898 -2934 444134
rect -2698 443898 -2614 444134
rect -2378 443898 -2346 444134
rect -2966 434454 -2346 443898
rect -2966 434218 -2934 434454
rect -2698 434218 -2614 434454
rect -2378 434218 -2346 434454
rect -2966 434134 -2346 434218
rect -2966 433898 -2934 434134
rect -2698 433898 -2614 434134
rect -2378 433898 -2346 434134
rect -2966 424454 -2346 433898
rect -2966 424218 -2934 424454
rect -2698 424218 -2614 424454
rect -2378 424218 -2346 424454
rect -2966 424134 -2346 424218
rect -2966 423898 -2934 424134
rect -2698 423898 -2614 424134
rect -2378 423898 -2346 424134
rect -2966 414454 -2346 423898
rect -2966 414218 -2934 414454
rect -2698 414218 -2614 414454
rect -2378 414218 -2346 414454
rect -2966 414134 -2346 414218
rect -2966 413898 -2934 414134
rect -2698 413898 -2614 414134
rect -2378 413898 -2346 414134
rect -2966 404454 -2346 413898
rect -2966 404218 -2934 404454
rect -2698 404218 -2614 404454
rect -2378 404218 -2346 404454
rect -2966 404134 -2346 404218
rect -2966 403898 -2934 404134
rect -2698 403898 -2614 404134
rect -2378 403898 -2346 404134
rect -2966 394454 -2346 403898
rect -2966 394218 -2934 394454
rect -2698 394218 -2614 394454
rect -2378 394218 -2346 394454
rect -2966 394134 -2346 394218
rect -2966 393898 -2934 394134
rect -2698 393898 -2614 394134
rect -2378 393898 -2346 394134
rect -2966 384454 -2346 393898
rect -2966 384218 -2934 384454
rect -2698 384218 -2614 384454
rect -2378 384218 -2346 384454
rect -2966 384134 -2346 384218
rect -2966 383898 -2934 384134
rect -2698 383898 -2614 384134
rect -2378 383898 -2346 384134
rect -2966 374454 -2346 383898
rect -2966 374218 -2934 374454
rect -2698 374218 -2614 374454
rect -2378 374218 -2346 374454
rect -2966 374134 -2346 374218
rect -2966 373898 -2934 374134
rect -2698 373898 -2614 374134
rect -2378 373898 -2346 374134
rect -2966 364454 -2346 373898
rect -2966 364218 -2934 364454
rect -2698 364218 -2614 364454
rect -2378 364218 -2346 364454
rect -2966 364134 -2346 364218
rect -2966 363898 -2934 364134
rect -2698 363898 -2614 364134
rect -2378 363898 -2346 364134
rect -2966 354454 -2346 363898
rect -2966 354218 -2934 354454
rect -2698 354218 -2614 354454
rect -2378 354218 -2346 354454
rect -2966 354134 -2346 354218
rect -2966 353898 -2934 354134
rect -2698 353898 -2614 354134
rect -2378 353898 -2346 354134
rect -2966 344454 -2346 353898
rect -2966 344218 -2934 344454
rect -2698 344218 -2614 344454
rect -2378 344218 -2346 344454
rect -2966 344134 -2346 344218
rect -2966 343898 -2934 344134
rect -2698 343898 -2614 344134
rect -2378 343898 -2346 344134
rect -2966 334454 -2346 343898
rect -2966 334218 -2934 334454
rect -2698 334218 -2614 334454
rect -2378 334218 -2346 334454
rect -2966 334134 -2346 334218
rect -2966 333898 -2934 334134
rect -2698 333898 -2614 334134
rect -2378 333898 -2346 334134
rect -2966 324454 -2346 333898
rect -2966 324218 -2934 324454
rect -2698 324218 -2614 324454
rect -2378 324218 -2346 324454
rect -2966 324134 -2346 324218
rect -2966 323898 -2934 324134
rect -2698 323898 -2614 324134
rect -2378 323898 -2346 324134
rect -2966 314454 -2346 323898
rect -2966 314218 -2934 314454
rect -2698 314218 -2614 314454
rect -2378 314218 -2346 314454
rect -2966 314134 -2346 314218
rect -2966 313898 -2934 314134
rect -2698 313898 -2614 314134
rect -2378 313898 -2346 314134
rect -2966 304454 -2346 313898
rect -2966 304218 -2934 304454
rect -2698 304218 -2614 304454
rect -2378 304218 -2346 304454
rect -2966 304134 -2346 304218
rect -2966 303898 -2934 304134
rect -2698 303898 -2614 304134
rect -2378 303898 -2346 304134
rect -2966 294454 -2346 303898
rect -2966 294218 -2934 294454
rect -2698 294218 -2614 294454
rect -2378 294218 -2346 294454
rect -2966 294134 -2346 294218
rect -2966 293898 -2934 294134
rect -2698 293898 -2614 294134
rect -2378 293898 -2346 294134
rect -2966 284454 -2346 293898
rect -2966 284218 -2934 284454
rect -2698 284218 -2614 284454
rect -2378 284218 -2346 284454
rect -2966 284134 -2346 284218
rect -2966 283898 -2934 284134
rect -2698 283898 -2614 284134
rect -2378 283898 -2346 284134
rect -2966 274454 -2346 283898
rect -2966 274218 -2934 274454
rect -2698 274218 -2614 274454
rect -2378 274218 -2346 274454
rect -2966 274134 -2346 274218
rect -2966 273898 -2934 274134
rect -2698 273898 -2614 274134
rect -2378 273898 -2346 274134
rect -2966 264454 -2346 273898
rect -2966 264218 -2934 264454
rect -2698 264218 -2614 264454
rect -2378 264218 -2346 264454
rect -2966 264134 -2346 264218
rect -2966 263898 -2934 264134
rect -2698 263898 -2614 264134
rect -2378 263898 -2346 264134
rect -2966 254454 -2346 263898
rect -2966 254218 -2934 254454
rect -2698 254218 -2614 254454
rect -2378 254218 -2346 254454
rect -2966 254134 -2346 254218
rect -2966 253898 -2934 254134
rect -2698 253898 -2614 254134
rect -2378 253898 -2346 254134
rect -2966 244454 -2346 253898
rect -2966 244218 -2934 244454
rect -2698 244218 -2614 244454
rect -2378 244218 -2346 244454
rect -2966 244134 -2346 244218
rect -2966 243898 -2934 244134
rect -2698 243898 -2614 244134
rect -2378 243898 -2346 244134
rect -2966 234454 -2346 243898
rect -2966 234218 -2934 234454
rect -2698 234218 -2614 234454
rect -2378 234218 -2346 234454
rect -2966 234134 -2346 234218
rect -2966 233898 -2934 234134
rect -2698 233898 -2614 234134
rect -2378 233898 -2346 234134
rect -2966 224454 -2346 233898
rect -2966 224218 -2934 224454
rect -2698 224218 -2614 224454
rect -2378 224218 -2346 224454
rect -2966 224134 -2346 224218
rect -2966 223898 -2934 224134
rect -2698 223898 -2614 224134
rect -2378 223898 -2346 224134
rect -2966 214454 -2346 223898
rect -2966 214218 -2934 214454
rect -2698 214218 -2614 214454
rect -2378 214218 -2346 214454
rect -2966 214134 -2346 214218
rect -2966 213898 -2934 214134
rect -2698 213898 -2614 214134
rect -2378 213898 -2346 214134
rect -2966 204454 -2346 213898
rect -2966 204218 -2934 204454
rect -2698 204218 -2614 204454
rect -2378 204218 -2346 204454
rect -2966 204134 -2346 204218
rect -2966 203898 -2934 204134
rect -2698 203898 -2614 204134
rect -2378 203898 -2346 204134
rect -2966 194454 -2346 203898
rect -2966 194218 -2934 194454
rect -2698 194218 -2614 194454
rect -2378 194218 -2346 194454
rect -2966 194134 -2346 194218
rect -2966 193898 -2934 194134
rect -2698 193898 -2614 194134
rect -2378 193898 -2346 194134
rect -2966 184454 -2346 193898
rect -2966 184218 -2934 184454
rect -2698 184218 -2614 184454
rect -2378 184218 -2346 184454
rect -2966 184134 -2346 184218
rect -2966 183898 -2934 184134
rect -2698 183898 -2614 184134
rect -2378 183898 -2346 184134
rect -2966 174454 -2346 183898
rect -2966 174218 -2934 174454
rect -2698 174218 -2614 174454
rect -2378 174218 -2346 174454
rect -2966 174134 -2346 174218
rect -2966 173898 -2934 174134
rect -2698 173898 -2614 174134
rect -2378 173898 -2346 174134
rect -2966 164454 -2346 173898
rect -2966 164218 -2934 164454
rect -2698 164218 -2614 164454
rect -2378 164218 -2346 164454
rect -2966 164134 -2346 164218
rect -2966 163898 -2934 164134
rect -2698 163898 -2614 164134
rect -2378 163898 -2346 164134
rect -2966 154454 -2346 163898
rect -2966 154218 -2934 154454
rect -2698 154218 -2614 154454
rect -2378 154218 -2346 154454
rect -2966 154134 -2346 154218
rect -2966 153898 -2934 154134
rect -2698 153898 -2614 154134
rect -2378 153898 -2346 154134
rect -2966 144454 -2346 153898
rect -2966 144218 -2934 144454
rect -2698 144218 -2614 144454
rect -2378 144218 -2346 144454
rect -2966 144134 -2346 144218
rect -2966 143898 -2934 144134
rect -2698 143898 -2614 144134
rect -2378 143898 -2346 144134
rect -2966 134454 -2346 143898
rect -2966 134218 -2934 134454
rect -2698 134218 -2614 134454
rect -2378 134218 -2346 134454
rect -2966 134134 -2346 134218
rect -2966 133898 -2934 134134
rect -2698 133898 -2614 134134
rect -2378 133898 -2346 134134
rect -2966 124454 -2346 133898
rect -2966 124218 -2934 124454
rect -2698 124218 -2614 124454
rect -2378 124218 -2346 124454
rect -2966 124134 -2346 124218
rect -2966 123898 -2934 124134
rect -2698 123898 -2614 124134
rect -2378 123898 -2346 124134
rect -2966 114454 -2346 123898
rect -2966 114218 -2934 114454
rect -2698 114218 -2614 114454
rect -2378 114218 -2346 114454
rect -2966 114134 -2346 114218
rect -2966 113898 -2934 114134
rect -2698 113898 -2614 114134
rect -2378 113898 -2346 114134
rect -2966 104454 -2346 113898
rect -2966 104218 -2934 104454
rect -2698 104218 -2614 104454
rect -2378 104218 -2346 104454
rect -2966 104134 -2346 104218
rect -2966 103898 -2934 104134
rect -2698 103898 -2614 104134
rect -2378 103898 -2346 104134
rect -2966 94454 -2346 103898
rect -2966 94218 -2934 94454
rect -2698 94218 -2614 94454
rect -2378 94218 -2346 94454
rect -2966 94134 -2346 94218
rect -2966 93898 -2934 94134
rect -2698 93898 -2614 94134
rect -2378 93898 -2346 94134
rect -2966 84454 -2346 93898
rect -2966 84218 -2934 84454
rect -2698 84218 -2614 84454
rect -2378 84218 -2346 84454
rect -2966 84134 -2346 84218
rect -2966 83898 -2934 84134
rect -2698 83898 -2614 84134
rect -2378 83898 -2346 84134
rect -2966 74454 -2346 83898
rect -2966 74218 -2934 74454
rect -2698 74218 -2614 74454
rect -2378 74218 -2346 74454
rect -2966 74134 -2346 74218
rect -2966 73898 -2934 74134
rect -2698 73898 -2614 74134
rect -2378 73898 -2346 74134
rect -2966 64454 -2346 73898
rect -2966 64218 -2934 64454
rect -2698 64218 -2614 64454
rect -2378 64218 -2346 64454
rect -2966 64134 -2346 64218
rect -2966 63898 -2934 64134
rect -2698 63898 -2614 64134
rect -2378 63898 -2346 64134
rect -2966 54454 -2346 63898
rect -2966 54218 -2934 54454
rect -2698 54218 -2614 54454
rect -2378 54218 -2346 54454
rect -2966 54134 -2346 54218
rect -2966 53898 -2934 54134
rect -2698 53898 -2614 54134
rect -2378 53898 -2346 54134
rect -2966 44454 -2346 53898
rect -2966 44218 -2934 44454
rect -2698 44218 -2614 44454
rect -2378 44218 -2346 44454
rect -2966 44134 -2346 44218
rect -2966 43898 -2934 44134
rect -2698 43898 -2614 44134
rect -2378 43898 -2346 44134
rect -2966 34454 -2346 43898
rect -2966 34218 -2934 34454
rect -2698 34218 -2614 34454
rect -2378 34218 -2346 34454
rect -2966 34134 -2346 34218
rect -2966 33898 -2934 34134
rect -2698 33898 -2614 34134
rect -2378 33898 -2346 34134
rect -2966 -1306 -2346 33898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 698174 -1386 704282
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 284339 699820 284405 699821
rect 284339 699756 284340 699820
rect 284404 699756 284405 699820
rect 284339 699755 284405 699756
rect -2006 697938 -1974 698174
rect -1738 697938 -1654 698174
rect -1418 697938 -1386 698174
rect -2006 697854 -1386 697938
rect -2006 697618 -1974 697854
rect -1738 697618 -1654 697854
rect -1418 697618 -1386 697854
rect -2006 688174 -1386 697618
rect -2006 687938 -1974 688174
rect -1738 687938 -1654 688174
rect -1418 687938 -1386 688174
rect -2006 687854 -1386 687938
rect -2006 687618 -1974 687854
rect -1738 687618 -1654 687854
rect -1418 687618 -1386 687854
rect -2006 678174 -1386 687618
rect 9811 684316 9877 684317
rect 9811 684252 9812 684316
rect 9876 684252 9877 684316
rect 9811 684251 9877 684252
rect -2006 677938 -1974 678174
rect -1738 677938 -1654 678174
rect -1418 677938 -1386 678174
rect -2006 677854 -1386 677938
rect -2006 677618 -1974 677854
rect -1738 677618 -1654 677854
rect -1418 677618 -1386 677854
rect -2006 668174 -1386 677618
rect 3371 671260 3437 671261
rect 3371 671196 3372 671260
rect 3436 671196 3437 671260
rect 3371 671195 3437 671196
rect -2006 667938 -1974 668174
rect -1738 667938 -1654 668174
rect -1418 667938 -1386 668174
rect -2006 667854 -1386 667938
rect -2006 667618 -1974 667854
rect -1738 667618 -1654 667854
rect -1418 667618 -1386 667854
rect -2006 658174 -1386 667618
rect -2006 657938 -1974 658174
rect -1738 657938 -1654 658174
rect -1418 657938 -1386 658174
rect -2006 657854 -1386 657938
rect -2006 657618 -1974 657854
rect -1738 657618 -1654 657854
rect -1418 657618 -1386 657854
rect -2006 648174 -1386 657618
rect -2006 647938 -1974 648174
rect -1738 647938 -1654 648174
rect -1418 647938 -1386 648174
rect -2006 647854 -1386 647938
rect -2006 647618 -1974 647854
rect -1738 647618 -1654 647854
rect -1418 647618 -1386 647854
rect -2006 638174 -1386 647618
rect -2006 637938 -1974 638174
rect -1738 637938 -1654 638174
rect -1418 637938 -1386 638174
rect -2006 637854 -1386 637938
rect -2006 637618 -1974 637854
rect -1738 637618 -1654 637854
rect -1418 637618 -1386 637854
rect -2006 628174 -1386 637618
rect -2006 627938 -1974 628174
rect -1738 627938 -1654 628174
rect -1418 627938 -1386 628174
rect -2006 627854 -1386 627938
rect -2006 627618 -1974 627854
rect -1738 627618 -1654 627854
rect -1418 627618 -1386 627854
rect -2006 618174 -1386 627618
rect -2006 617938 -1974 618174
rect -1738 617938 -1654 618174
rect -1418 617938 -1386 618174
rect -2006 617854 -1386 617938
rect -2006 617618 -1974 617854
rect -1738 617618 -1654 617854
rect -1418 617618 -1386 617854
rect -2006 608174 -1386 617618
rect -2006 607938 -1974 608174
rect -1738 607938 -1654 608174
rect -1418 607938 -1386 608174
rect -2006 607854 -1386 607938
rect -2006 607618 -1974 607854
rect -1738 607618 -1654 607854
rect -1418 607618 -1386 607854
rect -2006 598174 -1386 607618
rect -2006 597938 -1974 598174
rect -1738 597938 -1654 598174
rect -1418 597938 -1386 598174
rect -2006 597854 -1386 597938
rect -2006 597618 -1974 597854
rect -1738 597618 -1654 597854
rect -1418 597618 -1386 597854
rect -2006 588174 -1386 597618
rect -2006 587938 -1974 588174
rect -1738 587938 -1654 588174
rect -1418 587938 -1386 588174
rect -2006 587854 -1386 587938
rect -2006 587618 -1974 587854
rect -1738 587618 -1654 587854
rect -1418 587618 -1386 587854
rect -2006 578174 -1386 587618
rect -2006 577938 -1974 578174
rect -1738 577938 -1654 578174
rect -1418 577938 -1386 578174
rect -2006 577854 -1386 577938
rect -2006 577618 -1974 577854
rect -1738 577618 -1654 577854
rect -1418 577618 -1386 577854
rect -2006 568174 -1386 577618
rect -2006 567938 -1974 568174
rect -1738 567938 -1654 568174
rect -1418 567938 -1386 568174
rect -2006 567854 -1386 567938
rect -2006 567618 -1974 567854
rect -1738 567618 -1654 567854
rect -1418 567618 -1386 567854
rect -2006 558174 -1386 567618
rect -2006 557938 -1974 558174
rect -1738 557938 -1654 558174
rect -1418 557938 -1386 558174
rect -2006 557854 -1386 557938
rect -2006 557618 -1974 557854
rect -1738 557618 -1654 557854
rect -1418 557618 -1386 557854
rect -2006 548174 -1386 557618
rect -2006 547938 -1974 548174
rect -1738 547938 -1654 548174
rect -1418 547938 -1386 548174
rect -2006 547854 -1386 547938
rect -2006 547618 -1974 547854
rect -1738 547618 -1654 547854
rect -1418 547618 -1386 547854
rect -2006 538174 -1386 547618
rect -2006 537938 -1974 538174
rect -1738 537938 -1654 538174
rect -1418 537938 -1386 538174
rect -2006 537854 -1386 537938
rect -2006 537618 -1974 537854
rect -1738 537618 -1654 537854
rect -1418 537618 -1386 537854
rect -2006 528174 -1386 537618
rect -2006 527938 -1974 528174
rect -1738 527938 -1654 528174
rect -1418 527938 -1386 528174
rect -2006 527854 -1386 527938
rect -2006 527618 -1974 527854
rect -1738 527618 -1654 527854
rect -1418 527618 -1386 527854
rect 2819 527916 2885 527917
rect 2819 527852 2820 527916
rect 2884 527852 2885 527916
rect 2819 527851 2885 527852
rect -2006 518174 -1386 527618
rect -2006 517938 -1974 518174
rect -1738 517938 -1654 518174
rect -1418 517938 -1386 518174
rect -2006 517854 -1386 517938
rect -2006 517618 -1974 517854
rect -1738 517618 -1654 517854
rect -1418 517618 -1386 517854
rect -2006 508174 -1386 517618
rect -2006 507938 -1974 508174
rect -1738 507938 -1654 508174
rect -1418 507938 -1386 508174
rect -2006 507854 -1386 507938
rect -2006 507618 -1974 507854
rect -1738 507618 -1654 507854
rect -1418 507618 -1386 507854
rect -2006 498174 -1386 507618
rect -2006 497938 -1974 498174
rect -1738 497938 -1654 498174
rect -1418 497938 -1386 498174
rect -2006 497854 -1386 497938
rect -2006 497618 -1974 497854
rect -1738 497618 -1654 497854
rect -1418 497618 -1386 497854
rect -2006 488174 -1386 497618
rect -2006 487938 -1974 488174
rect -1738 487938 -1654 488174
rect -1418 487938 -1386 488174
rect -2006 487854 -1386 487938
rect -2006 487618 -1974 487854
rect -1738 487618 -1654 487854
rect -1418 487618 -1386 487854
rect -2006 478174 -1386 487618
rect -2006 477938 -1974 478174
rect -1738 477938 -1654 478174
rect -1418 477938 -1386 478174
rect -2006 477854 -1386 477938
rect -2006 477618 -1974 477854
rect -1738 477618 -1654 477854
rect -1418 477618 -1386 477854
rect -2006 468174 -1386 477618
rect 1899 475692 1965 475693
rect 1899 475628 1900 475692
rect 1964 475628 1965 475692
rect 1899 475627 1965 475628
rect -2006 467938 -1974 468174
rect -1738 467938 -1654 468174
rect -1418 467938 -1386 468174
rect -2006 467854 -1386 467938
rect -2006 467618 -1974 467854
rect -1738 467618 -1654 467854
rect -1418 467618 -1386 467854
rect -2006 458174 -1386 467618
rect -2006 457938 -1974 458174
rect -1738 457938 -1654 458174
rect -1418 457938 -1386 458174
rect -2006 457854 -1386 457938
rect -2006 457618 -1974 457854
rect -1738 457618 -1654 457854
rect -1418 457618 -1386 457854
rect -2006 448174 -1386 457618
rect -2006 447938 -1974 448174
rect -1738 447938 -1654 448174
rect -1418 447938 -1386 448174
rect -2006 447854 -1386 447938
rect -2006 447618 -1974 447854
rect -1738 447618 -1654 447854
rect -1418 447618 -1386 447854
rect -2006 438174 -1386 447618
rect -2006 437938 -1974 438174
rect -1738 437938 -1654 438174
rect -1418 437938 -1386 438174
rect -2006 437854 -1386 437938
rect -2006 437618 -1974 437854
rect -1738 437618 -1654 437854
rect -1418 437618 -1386 437854
rect -2006 428174 -1386 437618
rect -2006 427938 -1974 428174
rect -1738 427938 -1654 428174
rect -1418 427938 -1386 428174
rect -2006 427854 -1386 427938
rect -2006 427618 -1974 427854
rect -1738 427618 -1654 427854
rect -1418 427618 -1386 427854
rect -2006 418174 -1386 427618
rect -2006 417938 -1974 418174
rect -1738 417938 -1654 418174
rect -1418 417938 -1386 418174
rect -2006 417854 -1386 417938
rect -2006 417618 -1974 417854
rect -1738 417618 -1654 417854
rect -1418 417618 -1386 417854
rect -2006 408174 -1386 417618
rect -2006 407938 -1974 408174
rect -1738 407938 -1654 408174
rect -1418 407938 -1386 408174
rect -2006 407854 -1386 407938
rect -2006 407618 -1974 407854
rect -1738 407618 -1654 407854
rect -1418 407618 -1386 407854
rect -2006 398174 -1386 407618
rect -2006 397938 -1974 398174
rect -1738 397938 -1654 398174
rect -1418 397938 -1386 398174
rect -2006 397854 -1386 397938
rect -2006 397618 -1974 397854
rect -1738 397618 -1654 397854
rect -1418 397618 -1386 397854
rect -2006 388174 -1386 397618
rect -2006 387938 -1974 388174
rect -1738 387938 -1654 388174
rect -1418 387938 -1386 388174
rect -2006 387854 -1386 387938
rect -2006 387618 -1974 387854
rect -1738 387618 -1654 387854
rect -1418 387618 -1386 387854
rect -2006 378174 -1386 387618
rect -2006 377938 -1974 378174
rect -1738 377938 -1654 378174
rect -1418 377938 -1386 378174
rect -2006 377854 -1386 377938
rect -2006 377618 -1974 377854
rect -1738 377618 -1654 377854
rect -1418 377618 -1386 377854
rect -2006 368174 -1386 377618
rect 59 371652 125 371653
rect 59 371588 60 371652
rect 124 371588 125 371652
rect 59 371587 125 371588
rect -2006 367938 -1974 368174
rect -1738 367938 -1654 368174
rect -1418 367938 -1386 368174
rect -2006 367854 -1386 367938
rect -2006 367618 -1974 367854
rect -1738 367618 -1654 367854
rect -1418 367618 -1386 367854
rect -2006 358174 -1386 367618
rect -2006 357938 -1974 358174
rect -1738 357938 -1654 358174
rect -1418 357938 -1386 358174
rect -2006 357854 -1386 357938
rect -2006 357618 -1974 357854
rect -1738 357618 -1654 357854
rect -1418 357618 -1386 357854
rect -2006 348174 -1386 357618
rect -2006 347938 -1974 348174
rect -1738 347938 -1654 348174
rect -1418 347938 -1386 348174
rect -2006 347854 -1386 347938
rect -2006 347618 -1974 347854
rect -1738 347618 -1654 347854
rect -1418 347618 -1386 347854
rect -2006 338174 -1386 347618
rect -2006 337938 -1974 338174
rect -1738 337938 -1654 338174
rect -1418 337938 -1386 338174
rect -2006 337854 -1386 337938
rect -2006 337618 -1974 337854
rect -1738 337618 -1654 337854
rect -1418 337618 -1386 337854
rect -2006 328174 -1386 337618
rect -2006 327938 -1974 328174
rect -1738 327938 -1654 328174
rect -1418 327938 -1386 328174
rect -2006 327854 -1386 327938
rect -2006 327618 -1974 327854
rect -1738 327618 -1654 327854
rect -1418 327618 -1386 327854
rect -2006 318174 -1386 327618
rect -2006 317938 -1974 318174
rect -1738 317938 -1654 318174
rect -1418 317938 -1386 318174
rect -2006 317854 -1386 317938
rect -2006 317618 -1974 317854
rect -1738 317618 -1654 317854
rect -1418 317618 -1386 317854
rect -2006 308174 -1386 317618
rect -2006 307938 -1974 308174
rect -1738 307938 -1654 308174
rect -1418 307938 -1386 308174
rect -2006 307854 -1386 307938
rect -2006 307618 -1974 307854
rect -1738 307618 -1654 307854
rect -1418 307618 -1386 307854
rect -2006 298174 -1386 307618
rect -2006 297938 -1974 298174
rect -1738 297938 -1654 298174
rect -1418 297938 -1386 298174
rect -2006 297854 -1386 297938
rect -2006 297618 -1974 297854
rect -1738 297618 -1654 297854
rect -1418 297618 -1386 297854
rect -2006 288174 -1386 297618
rect -2006 287938 -1974 288174
rect -1738 287938 -1654 288174
rect -1418 287938 -1386 288174
rect -2006 287854 -1386 287938
rect -2006 287618 -1974 287854
rect -1738 287618 -1654 287854
rect -1418 287618 -1386 287854
rect -2006 278174 -1386 287618
rect -2006 277938 -1974 278174
rect -1738 277938 -1654 278174
rect -1418 277938 -1386 278174
rect -2006 277854 -1386 277938
rect -2006 277618 -1974 277854
rect -1738 277618 -1654 277854
rect -1418 277618 -1386 277854
rect -2006 268174 -1386 277618
rect -2006 267938 -1974 268174
rect -1738 267938 -1654 268174
rect -1418 267938 -1386 268174
rect -2006 267854 -1386 267938
rect -2006 267618 -1974 267854
rect -1738 267618 -1654 267854
rect -1418 267618 -1386 267854
rect -2006 258174 -1386 267618
rect -2006 257938 -1974 258174
rect -1738 257938 -1654 258174
rect -1418 257938 -1386 258174
rect -2006 257854 -1386 257938
rect -2006 257618 -1974 257854
rect -1738 257618 -1654 257854
rect -1418 257618 -1386 257854
rect -2006 248174 -1386 257618
rect -2006 247938 -1974 248174
rect -1738 247938 -1654 248174
rect -1418 247938 -1386 248174
rect -2006 247854 -1386 247938
rect -2006 247618 -1974 247854
rect -1738 247618 -1654 247854
rect -1418 247618 -1386 247854
rect -2006 238174 -1386 247618
rect -2006 237938 -1974 238174
rect -1738 237938 -1654 238174
rect -1418 237938 -1386 238174
rect -2006 237854 -1386 237938
rect -2006 237618 -1974 237854
rect -1738 237618 -1654 237854
rect -1418 237618 -1386 237854
rect -2006 228174 -1386 237618
rect -2006 227938 -1974 228174
rect -1738 227938 -1654 228174
rect -1418 227938 -1386 228174
rect -2006 227854 -1386 227938
rect -2006 227618 -1974 227854
rect -1738 227618 -1654 227854
rect -1418 227618 -1386 227854
rect -2006 218174 -1386 227618
rect -2006 217938 -1974 218174
rect -1738 217938 -1654 218174
rect -1418 217938 -1386 218174
rect -2006 217854 -1386 217938
rect -2006 217618 -1974 217854
rect -1738 217618 -1654 217854
rect -1418 217618 -1386 217854
rect -2006 208174 -1386 217618
rect -2006 207938 -1974 208174
rect -1738 207938 -1654 208174
rect -1418 207938 -1386 208174
rect -2006 207854 -1386 207938
rect -2006 207618 -1974 207854
rect -1738 207618 -1654 207854
rect -1418 207618 -1386 207854
rect -2006 198174 -1386 207618
rect -2006 197938 -1974 198174
rect -1738 197938 -1654 198174
rect -1418 197938 -1386 198174
rect -2006 197854 -1386 197938
rect -2006 197618 -1974 197854
rect -1738 197618 -1654 197854
rect -1418 197618 -1386 197854
rect -2006 188174 -1386 197618
rect -2006 187938 -1974 188174
rect -1738 187938 -1654 188174
rect -1418 187938 -1386 188174
rect -2006 187854 -1386 187938
rect -2006 187618 -1974 187854
rect -1738 187618 -1654 187854
rect -1418 187618 -1386 187854
rect -2006 178174 -1386 187618
rect -2006 177938 -1974 178174
rect -1738 177938 -1654 178174
rect -1418 177938 -1386 178174
rect -2006 177854 -1386 177938
rect -2006 177618 -1974 177854
rect -1738 177618 -1654 177854
rect -1418 177618 -1386 177854
rect -2006 168174 -1386 177618
rect -2006 167938 -1974 168174
rect -1738 167938 -1654 168174
rect -1418 167938 -1386 168174
rect -2006 167854 -1386 167938
rect -2006 167618 -1974 167854
rect -1738 167618 -1654 167854
rect -1418 167618 -1386 167854
rect -2006 158174 -1386 167618
rect -2006 157938 -1974 158174
rect -1738 157938 -1654 158174
rect -1418 157938 -1386 158174
rect -2006 157854 -1386 157938
rect -2006 157618 -1974 157854
rect -1738 157618 -1654 157854
rect -1418 157618 -1386 157854
rect -2006 148174 -1386 157618
rect -2006 147938 -1974 148174
rect -1738 147938 -1654 148174
rect -1418 147938 -1386 148174
rect -2006 147854 -1386 147938
rect -2006 147618 -1974 147854
rect -1738 147618 -1654 147854
rect -1418 147618 -1386 147854
rect -2006 138174 -1386 147618
rect -2006 137938 -1974 138174
rect -1738 137938 -1654 138174
rect -1418 137938 -1386 138174
rect -2006 137854 -1386 137938
rect -2006 137618 -1974 137854
rect -1738 137618 -1654 137854
rect -1418 137618 -1386 137854
rect -2006 128174 -1386 137618
rect -2006 127938 -1974 128174
rect -1738 127938 -1654 128174
rect -1418 127938 -1386 128174
rect -2006 127854 -1386 127938
rect -2006 127618 -1974 127854
rect -1738 127618 -1654 127854
rect -1418 127618 -1386 127854
rect -2006 118174 -1386 127618
rect -2006 117938 -1974 118174
rect -1738 117938 -1654 118174
rect -1418 117938 -1386 118174
rect -2006 117854 -1386 117938
rect -2006 117618 -1974 117854
rect -1738 117618 -1654 117854
rect -1418 117618 -1386 117854
rect -2006 108174 -1386 117618
rect -2006 107938 -1974 108174
rect -1738 107938 -1654 108174
rect -1418 107938 -1386 108174
rect -2006 107854 -1386 107938
rect -2006 107618 -1974 107854
rect -1738 107618 -1654 107854
rect -1418 107618 -1386 107854
rect -2006 98174 -1386 107618
rect -2006 97938 -1974 98174
rect -1738 97938 -1654 98174
rect -1418 97938 -1386 98174
rect -2006 97854 -1386 97938
rect -2006 97618 -1974 97854
rect -1738 97618 -1654 97854
rect -1418 97618 -1386 97854
rect -2006 88174 -1386 97618
rect -2006 87938 -1974 88174
rect -1738 87938 -1654 88174
rect -1418 87938 -1386 88174
rect -2006 87854 -1386 87938
rect -2006 87618 -1974 87854
rect -1738 87618 -1654 87854
rect -1418 87618 -1386 87854
rect -2006 78174 -1386 87618
rect -2006 77938 -1974 78174
rect -1738 77938 -1654 78174
rect -1418 77938 -1386 78174
rect -2006 77854 -1386 77938
rect -2006 77618 -1974 77854
rect -1738 77618 -1654 77854
rect -1418 77618 -1386 77854
rect -2006 68174 -1386 77618
rect -2006 67938 -1974 68174
rect -1738 67938 -1654 68174
rect -1418 67938 -1386 68174
rect -2006 67854 -1386 67938
rect -2006 67618 -1974 67854
rect -1738 67618 -1654 67854
rect -1418 67618 -1386 67854
rect -2006 58174 -1386 67618
rect -2006 57938 -1974 58174
rect -1738 57938 -1654 58174
rect -1418 57938 -1386 58174
rect -2006 57854 -1386 57938
rect -2006 57618 -1974 57854
rect -1738 57618 -1654 57854
rect -1418 57618 -1386 57854
rect -2006 48174 -1386 57618
rect -2006 47938 -1974 48174
rect -1738 47938 -1654 48174
rect -1418 47938 -1386 48174
rect -2006 47854 -1386 47938
rect -2006 47618 -1974 47854
rect -1738 47618 -1654 47854
rect -1418 47618 -1386 47854
rect -2006 38174 -1386 47618
rect -2006 37938 -1974 38174
rect -1738 37938 -1654 38174
rect -1418 37938 -1386 38174
rect -2006 37854 -1386 37938
rect -2006 37618 -1974 37854
rect -1738 37618 -1654 37854
rect -1418 37618 -1386 37854
rect -2006 -346 -1386 37618
rect 62 20093 122 371587
rect 1163 242860 1229 242861
rect 1163 242796 1164 242860
rect 1228 242796 1229 242860
rect 1163 242795 1229 242796
rect 979 213212 1045 213213
rect 979 213148 980 213212
rect 1044 213148 1045 213212
rect 979 213147 1045 213148
rect 982 76533 1042 213147
rect 979 76532 1045 76533
rect 979 76468 980 76532
rect 1044 76468 1045 76532
rect 979 76467 1045 76468
rect 1166 68237 1226 242795
rect 1902 68373 1962 475627
rect 2083 293180 2149 293181
rect 2083 293116 2084 293180
rect 2148 293116 2149 293180
rect 2083 293115 2149 293116
rect 1899 68372 1965 68373
rect 1899 68308 1900 68372
rect 1964 68308 1965 68372
rect 1899 68307 1965 68308
rect 1163 68236 1229 68237
rect 1163 68172 1164 68236
rect 1228 68172 1229 68236
rect 1163 68171 1229 68172
rect 2086 20365 2146 293115
rect 2822 242861 2882 527851
rect 3374 307053 3434 671195
rect 8891 632092 8957 632093
rect 8891 632028 8892 632092
rect 8956 632028 8957 632092
rect 8891 632027 8957 632028
rect 4659 619172 4725 619173
rect 4659 619108 4660 619172
rect 4724 619108 4725 619172
rect 4659 619107 4725 619108
rect 3555 345404 3621 345405
rect 3555 345340 3556 345404
rect 3620 345340 3621 345404
rect 3555 345339 3621 345340
rect 3371 307052 3437 307053
rect 3371 306988 3372 307052
rect 3436 306988 3437 307052
rect 3371 306987 3437 306988
rect 3371 267204 3437 267205
rect 3371 267140 3372 267204
rect 3436 267140 3437 267204
rect 3371 267139 3437 267140
rect 3003 254284 3069 254285
rect 3003 254220 3004 254284
rect 3068 254220 3069 254284
rect 3003 254219 3069 254220
rect 2819 242860 2885 242861
rect 2819 242796 2820 242860
rect 2884 242796 2885 242860
rect 2819 242795 2885 242796
rect 2635 213348 2701 213349
rect 2635 213284 2636 213348
rect 2700 213284 2701 213348
rect 2635 213283 2701 213284
rect 2638 73813 2698 213283
rect 3006 201925 3066 254219
rect 3003 201924 3069 201925
rect 3003 201860 3004 201924
rect 3068 201860 3069 201924
rect 3003 201859 3069 201860
rect 3006 200130 3066 201859
rect 2822 200070 3066 200130
rect 2822 188869 2882 200070
rect 2819 188868 2885 188869
rect 2819 188804 2820 188868
rect 2884 188804 2885 188868
rect 2819 188803 2885 188804
rect 2822 149837 2882 188803
rect 2819 149836 2885 149837
rect 2819 149772 2820 149836
rect 2884 149772 2885 149836
rect 2819 149771 2885 149772
rect 2822 97613 2882 149771
rect 3374 149701 3434 267139
rect 3558 155277 3618 345339
rect 3739 306236 3805 306237
rect 3739 306172 3740 306236
rect 3804 306172 3805 306236
rect 3739 306171 3805 306172
rect 3742 256733 3802 306171
rect 3739 256732 3805 256733
rect 3739 256668 3740 256732
rect 3804 256668 3805 256732
rect 3739 256667 3805 256668
rect 4107 162892 4173 162893
rect 4107 162828 4108 162892
rect 4172 162828 4173 162892
rect 4107 162827 4173 162828
rect 4110 156637 4170 162827
rect 4107 156636 4173 156637
rect 4107 156572 4108 156636
rect 4172 156572 4173 156636
rect 4107 156571 4173 156572
rect 3555 155276 3621 155277
rect 3555 155212 3556 155276
rect 3620 155212 3621 155276
rect 3555 155211 3621 155212
rect 4662 153781 4722 619107
rect 7419 580004 7485 580005
rect 7419 579940 7420 580004
rect 7484 579940 7485 580004
rect 7419 579939 7485 579940
rect 4843 514860 4909 514861
rect 4843 514796 4844 514860
rect 4908 514796 4909 514860
rect 4843 514795 4909 514796
rect 4659 153780 4725 153781
rect 4659 153716 4660 153780
rect 4724 153716 4725 153780
rect 4659 153715 4725 153716
rect 3371 149700 3437 149701
rect 3371 149636 3372 149700
rect 3436 149636 3437 149700
rect 3371 149635 3437 149636
rect 2819 97612 2885 97613
rect 2819 97548 2820 97612
rect 2884 97548 2885 97612
rect 2819 97547 2885 97548
rect 2822 84693 2882 97547
rect 4846 87549 4906 514795
rect 6131 410548 6197 410549
rect 6131 410484 6132 410548
rect 6196 410484 6197 410548
rect 6131 410483 6197 410484
rect 5395 213484 5461 213485
rect 5395 213420 5396 213484
rect 5460 213420 5461 213484
rect 5395 213419 5461 213420
rect 4843 87548 4909 87549
rect 4843 87484 4844 87548
rect 4908 87484 4909 87548
rect 4843 87483 4909 87484
rect 2819 84692 2885 84693
rect 2819 84628 2820 84692
rect 2884 84628 2885 84692
rect 2819 84627 2885 84628
rect 2635 73812 2701 73813
rect 2635 73748 2636 73812
rect 2700 73748 2701 73812
rect 2635 73747 2701 73748
rect 2822 58581 2882 84627
rect 3371 71636 3437 71637
rect 3371 71572 3372 71636
rect 3436 71572 3437 71636
rect 3371 71571 3437 71572
rect 2819 58580 2885 58581
rect 2819 58516 2820 58580
rect 2884 58516 2885 58580
rect 2819 58515 2885 58516
rect 2822 20637 2882 58515
rect 3374 22677 3434 71571
rect 5398 71093 5458 213419
rect 6134 152421 6194 410483
rect 6315 256732 6381 256733
rect 6315 256668 6316 256732
rect 6380 256668 6381 256732
rect 6315 256667 6381 256668
rect 6131 152420 6197 152421
rect 6131 152356 6132 152420
rect 6196 152356 6197 152420
rect 6131 152355 6197 152356
rect 5395 71092 5461 71093
rect 5395 71028 5396 71092
rect 5460 71028 5461 71092
rect 5395 71027 5461 71028
rect 3371 22676 3437 22677
rect 3371 22612 3372 22676
rect 3436 22612 3437 22676
rect 3371 22611 3437 22612
rect 6318 21725 6378 256667
rect 6683 213620 6749 213621
rect 6683 213556 6684 213620
rect 6748 213556 6749 213620
rect 6683 213555 6749 213556
rect 6686 66877 6746 213555
rect 7422 151061 7482 579939
rect 7603 319292 7669 319293
rect 7603 319228 7604 319292
rect 7668 319228 7669 319292
rect 7603 319227 7669 319228
rect 7419 151060 7485 151061
rect 7419 150996 7420 151060
rect 7484 150996 7485 151060
rect 7419 150995 7485 150996
rect 6683 66876 6749 66877
rect 6683 66812 6684 66876
rect 6748 66812 6749 66876
rect 6683 66811 6749 66812
rect 6315 21724 6381 21725
rect 6315 21660 6316 21724
rect 6380 21660 6381 21724
rect 6315 21659 6381 21660
rect 2819 20636 2885 20637
rect 2819 20572 2820 20636
rect 2884 20572 2885 20636
rect 2819 20571 2885 20572
rect 2083 20364 2149 20365
rect 2083 20300 2084 20364
rect 2148 20300 2149 20364
rect 2083 20299 2149 20300
rect 59 20092 125 20093
rect 59 20028 60 20092
rect 124 20028 125 20092
rect 59 20027 125 20028
rect 2822 19549 2882 20571
rect 2819 19548 2885 19549
rect 2819 19484 2820 19548
rect 2884 19484 2885 19548
rect 2819 19483 2885 19484
rect 7606 19277 7666 319227
rect 8155 196076 8221 196077
rect 8155 196012 8156 196076
rect 8220 196012 8221 196076
rect 8155 196011 8221 196012
rect 7971 194580 8037 194581
rect 7971 194516 7972 194580
rect 8036 194516 8037 194580
rect 7971 194515 8037 194516
rect 7974 178805 8034 194515
rect 7971 178804 8037 178805
rect 7971 178740 7972 178804
rect 8036 178740 8037 178804
rect 7971 178739 8037 178740
rect 8158 21861 8218 196011
rect 8894 69597 8954 632027
rect 9075 423604 9141 423605
rect 9075 423540 9076 423604
rect 9140 423540 9141 423604
rect 9075 423539 9141 423540
rect 9078 73949 9138 423539
rect 9814 364350 9874 684251
rect 282131 566948 282197 566949
rect 282131 566884 282132 566948
rect 282196 566884 282197 566948
rect 282131 566883 282197 566884
rect 17907 553892 17973 553893
rect 17907 553828 17908 553892
rect 17972 553828 17973 553892
rect 17907 553827 17973 553828
rect 12387 501804 12453 501805
rect 12387 501740 12388 501804
rect 12452 501740 12453 501804
rect 12387 501739 12453 501740
rect 11099 449580 11165 449581
rect 11099 449516 11100 449580
rect 11164 449516 11165 449580
rect 11099 449515 11165 449516
rect 9630 364290 9874 364350
rect 9443 213756 9509 213757
rect 9443 213692 9444 213756
rect 9508 213692 9509 213756
rect 9443 213691 9509 213692
rect 9446 178941 9506 213691
rect 9630 189141 9690 364290
rect 9811 358460 9877 358461
rect 9811 358396 9812 358460
rect 9876 358396 9877 358460
rect 9811 358395 9877 358396
rect 9814 196077 9874 358395
rect 10179 213892 10245 213893
rect 10179 213828 10180 213892
rect 10244 213828 10245 213892
rect 10179 213827 10245 213828
rect 9811 196076 9877 196077
rect 9811 196012 9812 196076
rect 9876 196012 9877 196076
rect 9811 196011 9877 196012
rect 10182 194581 10242 213827
rect 11102 213757 11162 449515
rect 12390 213893 12450 501739
rect 13859 462636 13925 462637
rect 13859 462572 13860 462636
rect 13924 462572 13925 462636
rect 13859 462571 13925 462572
rect 12387 213892 12453 213893
rect 12387 213828 12388 213892
rect 12452 213828 12453 213892
rect 12387 213827 12453 213828
rect 11099 213756 11165 213757
rect 11099 213692 11100 213756
rect 11164 213692 11165 213756
rect 11099 213691 11165 213692
rect 13862 213621 13922 462571
rect 15147 397492 15213 397493
rect 15147 397428 15148 397492
rect 15212 397428 15213 397492
rect 15147 397427 15213 397428
rect 13859 213620 13925 213621
rect 13859 213556 13860 213620
rect 13924 213556 13925 213620
rect 13859 213555 13925 213556
rect 15150 213485 15210 397427
rect 16619 307052 16685 307053
rect 16619 306988 16620 307052
rect 16684 306988 16685 307052
rect 16619 306987 16685 306988
rect 15147 213484 15213 213485
rect 15147 213420 15148 213484
rect 15212 213420 15213 213484
rect 15147 213419 15213 213420
rect 16622 213213 16682 306987
rect 17910 213349 17970 553827
rect 17907 213348 17973 213349
rect 17907 213284 17908 213348
rect 17972 213284 17973 213348
rect 17907 213283 17973 213284
rect 16619 213212 16685 213213
rect 16619 213148 16620 213212
rect 16684 213148 16685 213212
rect 16619 213147 16685 213148
rect 14065 208174 14385 208206
rect 14065 207938 14107 208174
rect 14343 207938 14385 208174
rect 14065 207854 14385 207938
rect 14065 207618 14107 207854
rect 14343 207618 14385 207854
rect 14065 207586 14385 207618
rect 21907 208174 22227 208206
rect 21907 207938 21949 208174
rect 22185 207938 22227 208174
rect 21907 207854 22227 207938
rect 21907 207618 21949 207854
rect 22185 207618 22227 207854
rect 21907 207586 22227 207618
rect 29749 208174 30069 208206
rect 29749 207938 29791 208174
rect 30027 207938 30069 208174
rect 29749 207854 30069 207938
rect 29749 207618 29791 207854
rect 30027 207618 30069 207854
rect 29749 207586 30069 207618
rect 37591 208174 37911 208206
rect 37591 207938 37633 208174
rect 37869 207938 37911 208174
rect 37591 207854 37911 207938
rect 37591 207618 37633 207854
rect 37869 207618 37911 207854
rect 37591 207586 37911 207618
rect 48197 208174 48517 208206
rect 48197 207938 48239 208174
rect 48475 207938 48517 208174
rect 48197 207854 48517 207938
rect 48197 207618 48239 207854
rect 48475 207618 48517 207854
rect 48197 207586 48517 207618
rect 56039 208174 56359 208206
rect 56039 207938 56081 208174
rect 56317 207938 56359 208174
rect 56039 207854 56359 207938
rect 56039 207618 56081 207854
rect 56317 207618 56359 207854
rect 56039 207586 56359 207618
rect 63881 208174 64201 208206
rect 63881 207938 63923 208174
rect 64159 207938 64201 208174
rect 63881 207854 64201 207938
rect 63881 207618 63923 207854
rect 64159 207618 64201 207854
rect 63881 207586 64201 207618
rect 71723 208174 72043 208206
rect 71723 207938 71765 208174
rect 72001 207938 72043 208174
rect 71723 207854 72043 207938
rect 71723 207618 71765 207854
rect 72001 207618 72043 207854
rect 71723 207586 72043 207618
rect 82329 208174 82649 208206
rect 82329 207938 82371 208174
rect 82607 207938 82649 208174
rect 82329 207854 82649 207938
rect 82329 207618 82371 207854
rect 82607 207618 82649 207854
rect 82329 207586 82649 207618
rect 90171 208174 90491 208206
rect 90171 207938 90213 208174
rect 90449 207938 90491 208174
rect 90171 207854 90491 207938
rect 90171 207618 90213 207854
rect 90449 207618 90491 207854
rect 90171 207586 90491 207618
rect 98013 208174 98333 208206
rect 98013 207938 98055 208174
rect 98291 207938 98333 208174
rect 98013 207854 98333 207938
rect 98013 207618 98055 207854
rect 98291 207618 98333 207854
rect 98013 207586 98333 207618
rect 105855 208174 106175 208206
rect 105855 207938 105897 208174
rect 106133 207938 106175 208174
rect 105855 207854 106175 207938
rect 105855 207618 105897 207854
rect 106133 207618 106175 207854
rect 105855 207586 106175 207618
rect 116461 208174 116781 208206
rect 116461 207938 116503 208174
rect 116739 207938 116781 208174
rect 116461 207854 116781 207938
rect 116461 207618 116503 207854
rect 116739 207618 116781 207854
rect 116461 207586 116781 207618
rect 124303 208174 124623 208206
rect 124303 207938 124345 208174
rect 124581 207938 124623 208174
rect 124303 207854 124623 207938
rect 124303 207618 124345 207854
rect 124581 207618 124623 207854
rect 124303 207586 124623 207618
rect 132145 208174 132465 208206
rect 132145 207938 132187 208174
rect 132423 207938 132465 208174
rect 132145 207854 132465 207938
rect 132145 207618 132187 207854
rect 132423 207618 132465 207854
rect 132145 207586 132465 207618
rect 139987 208174 140307 208206
rect 139987 207938 140029 208174
rect 140265 207938 140307 208174
rect 139987 207854 140307 207938
rect 139987 207618 140029 207854
rect 140265 207618 140307 207854
rect 139987 207586 140307 207618
rect 150593 208174 150913 208206
rect 150593 207938 150635 208174
rect 150871 207938 150913 208174
rect 150593 207854 150913 207938
rect 150593 207618 150635 207854
rect 150871 207618 150913 207854
rect 150593 207586 150913 207618
rect 158435 208174 158755 208206
rect 158435 207938 158477 208174
rect 158713 207938 158755 208174
rect 158435 207854 158755 207938
rect 158435 207618 158477 207854
rect 158713 207618 158755 207854
rect 158435 207586 158755 207618
rect 166277 208174 166597 208206
rect 166277 207938 166319 208174
rect 166555 207938 166597 208174
rect 166277 207854 166597 207938
rect 166277 207618 166319 207854
rect 166555 207618 166597 207854
rect 166277 207586 166597 207618
rect 174119 208174 174439 208206
rect 174119 207938 174161 208174
rect 174397 207938 174439 208174
rect 174119 207854 174439 207938
rect 174119 207618 174161 207854
rect 174397 207618 174439 207854
rect 174119 207586 174439 207618
rect 184725 208174 185045 208206
rect 184725 207938 184767 208174
rect 185003 207938 185045 208174
rect 184725 207854 185045 207938
rect 184725 207618 184767 207854
rect 185003 207618 185045 207854
rect 184725 207586 185045 207618
rect 192567 208174 192887 208206
rect 192567 207938 192609 208174
rect 192845 207938 192887 208174
rect 192567 207854 192887 207938
rect 192567 207618 192609 207854
rect 192845 207618 192887 207854
rect 192567 207586 192887 207618
rect 200409 208174 200729 208206
rect 200409 207938 200451 208174
rect 200687 207938 200729 208174
rect 200409 207854 200729 207938
rect 200409 207618 200451 207854
rect 200687 207618 200729 207854
rect 200409 207586 200729 207618
rect 208251 208174 208571 208206
rect 208251 207938 208293 208174
rect 208529 207938 208571 208174
rect 208251 207854 208571 207938
rect 208251 207618 208293 207854
rect 208529 207618 208571 207854
rect 208251 207586 208571 207618
rect 218857 208174 219177 208206
rect 218857 207938 218899 208174
rect 219135 207938 219177 208174
rect 218857 207854 219177 207938
rect 218857 207618 218899 207854
rect 219135 207618 219177 207854
rect 218857 207586 219177 207618
rect 226699 208174 227019 208206
rect 226699 207938 226741 208174
rect 226977 207938 227019 208174
rect 226699 207854 227019 207938
rect 226699 207618 226741 207854
rect 226977 207618 227019 207854
rect 226699 207586 227019 207618
rect 234541 208174 234861 208206
rect 234541 207938 234583 208174
rect 234819 207938 234861 208174
rect 234541 207854 234861 207938
rect 234541 207618 234583 207854
rect 234819 207618 234861 207854
rect 234541 207586 234861 207618
rect 242383 208174 242703 208206
rect 242383 207938 242425 208174
rect 242661 207938 242703 208174
rect 242383 207854 242703 207938
rect 242383 207618 242425 207854
rect 242661 207618 242703 207854
rect 242383 207586 242703 207618
rect 252989 208174 253309 208206
rect 252989 207938 253031 208174
rect 253267 207938 253309 208174
rect 252989 207854 253309 207938
rect 252989 207618 253031 207854
rect 253267 207618 253309 207854
rect 252989 207586 253309 207618
rect 260831 208174 261151 208206
rect 260831 207938 260873 208174
rect 261109 207938 261151 208174
rect 260831 207854 261151 207938
rect 260831 207618 260873 207854
rect 261109 207618 261151 207854
rect 260831 207586 261151 207618
rect 268673 208174 268993 208206
rect 268673 207938 268715 208174
rect 268951 207938 268993 208174
rect 268673 207854 268993 207938
rect 268673 207618 268715 207854
rect 268951 207618 268993 207854
rect 268673 207586 268993 207618
rect 276515 208174 276835 208206
rect 276515 207938 276557 208174
rect 276793 207938 276835 208174
rect 276515 207854 276835 207938
rect 276515 207618 276557 207854
rect 276793 207618 276835 207854
rect 276515 207586 276835 207618
rect 17986 204454 18306 204486
rect 17986 204218 18028 204454
rect 18264 204218 18306 204454
rect 17986 204134 18306 204218
rect 17986 203898 18028 204134
rect 18264 203898 18306 204134
rect 17986 203866 18306 203898
rect 25828 204454 26148 204486
rect 25828 204218 25870 204454
rect 26106 204218 26148 204454
rect 25828 204134 26148 204218
rect 25828 203898 25870 204134
rect 26106 203898 26148 204134
rect 25828 203866 26148 203898
rect 33670 204454 33990 204486
rect 33670 204218 33712 204454
rect 33948 204218 33990 204454
rect 33670 204134 33990 204218
rect 33670 203898 33712 204134
rect 33948 203898 33990 204134
rect 33670 203866 33990 203898
rect 41512 204454 41832 204486
rect 41512 204218 41554 204454
rect 41790 204218 41832 204454
rect 41512 204134 41832 204218
rect 41512 203898 41554 204134
rect 41790 203898 41832 204134
rect 41512 203866 41832 203898
rect 52118 204454 52438 204486
rect 52118 204218 52160 204454
rect 52396 204218 52438 204454
rect 52118 204134 52438 204218
rect 52118 203898 52160 204134
rect 52396 203898 52438 204134
rect 52118 203866 52438 203898
rect 59960 204454 60280 204486
rect 59960 204218 60002 204454
rect 60238 204218 60280 204454
rect 59960 204134 60280 204218
rect 59960 203898 60002 204134
rect 60238 203898 60280 204134
rect 59960 203866 60280 203898
rect 67802 204454 68122 204486
rect 67802 204218 67844 204454
rect 68080 204218 68122 204454
rect 67802 204134 68122 204218
rect 67802 203898 67844 204134
rect 68080 203898 68122 204134
rect 67802 203866 68122 203898
rect 75644 204454 75964 204486
rect 75644 204218 75686 204454
rect 75922 204218 75964 204454
rect 75644 204134 75964 204218
rect 75644 203898 75686 204134
rect 75922 203898 75964 204134
rect 75644 203866 75964 203898
rect 86250 204454 86570 204486
rect 86250 204218 86292 204454
rect 86528 204218 86570 204454
rect 86250 204134 86570 204218
rect 86250 203898 86292 204134
rect 86528 203898 86570 204134
rect 86250 203866 86570 203898
rect 94092 204454 94412 204486
rect 94092 204218 94134 204454
rect 94370 204218 94412 204454
rect 94092 204134 94412 204218
rect 94092 203898 94134 204134
rect 94370 203898 94412 204134
rect 94092 203866 94412 203898
rect 101934 204454 102254 204486
rect 101934 204218 101976 204454
rect 102212 204218 102254 204454
rect 101934 204134 102254 204218
rect 101934 203898 101976 204134
rect 102212 203898 102254 204134
rect 101934 203866 102254 203898
rect 109776 204454 110096 204486
rect 109776 204218 109818 204454
rect 110054 204218 110096 204454
rect 109776 204134 110096 204218
rect 109776 203898 109818 204134
rect 110054 203898 110096 204134
rect 109776 203866 110096 203898
rect 120382 204454 120702 204486
rect 120382 204218 120424 204454
rect 120660 204218 120702 204454
rect 120382 204134 120702 204218
rect 120382 203898 120424 204134
rect 120660 203898 120702 204134
rect 120382 203866 120702 203898
rect 128224 204454 128544 204486
rect 128224 204218 128266 204454
rect 128502 204218 128544 204454
rect 128224 204134 128544 204218
rect 128224 203898 128266 204134
rect 128502 203898 128544 204134
rect 128224 203866 128544 203898
rect 136066 204454 136386 204486
rect 136066 204218 136108 204454
rect 136344 204218 136386 204454
rect 136066 204134 136386 204218
rect 136066 203898 136108 204134
rect 136344 203898 136386 204134
rect 136066 203866 136386 203898
rect 143908 204454 144228 204486
rect 143908 204218 143950 204454
rect 144186 204218 144228 204454
rect 143908 204134 144228 204218
rect 143908 203898 143950 204134
rect 144186 203898 144228 204134
rect 143908 203866 144228 203898
rect 154514 204454 154834 204486
rect 154514 204218 154556 204454
rect 154792 204218 154834 204454
rect 154514 204134 154834 204218
rect 154514 203898 154556 204134
rect 154792 203898 154834 204134
rect 154514 203866 154834 203898
rect 162356 204454 162676 204486
rect 162356 204218 162398 204454
rect 162634 204218 162676 204454
rect 162356 204134 162676 204218
rect 162356 203898 162398 204134
rect 162634 203898 162676 204134
rect 162356 203866 162676 203898
rect 170198 204454 170518 204486
rect 170198 204218 170240 204454
rect 170476 204218 170518 204454
rect 170198 204134 170518 204218
rect 170198 203898 170240 204134
rect 170476 203898 170518 204134
rect 170198 203866 170518 203898
rect 178040 204454 178360 204486
rect 178040 204218 178082 204454
rect 178318 204218 178360 204454
rect 178040 204134 178360 204218
rect 178040 203898 178082 204134
rect 178318 203898 178360 204134
rect 178040 203866 178360 203898
rect 188646 204454 188966 204486
rect 188646 204218 188688 204454
rect 188924 204218 188966 204454
rect 188646 204134 188966 204218
rect 188646 203898 188688 204134
rect 188924 203898 188966 204134
rect 188646 203866 188966 203898
rect 196488 204454 196808 204486
rect 196488 204218 196530 204454
rect 196766 204218 196808 204454
rect 196488 204134 196808 204218
rect 196488 203898 196530 204134
rect 196766 203898 196808 204134
rect 196488 203866 196808 203898
rect 204330 204454 204650 204486
rect 204330 204218 204372 204454
rect 204608 204218 204650 204454
rect 204330 204134 204650 204218
rect 204330 203898 204372 204134
rect 204608 203898 204650 204134
rect 204330 203866 204650 203898
rect 212172 204454 212492 204486
rect 212172 204218 212214 204454
rect 212450 204218 212492 204454
rect 212172 204134 212492 204218
rect 212172 203898 212214 204134
rect 212450 203898 212492 204134
rect 212172 203866 212492 203898
rect 222778 204454 223098 204486
rect 222778 204218 222820 204454
rect 223056 204218 223098 204454
rect 222778 204134 223098 204218
rect 222778 203898 222820 204134
rect 223056 203898 223098 204134
rect 222778 203866 223098 203898
rect 230620 204454 230940 204486
rect 230620 204218 230662 204454
rect 230898 204218 230940 204454
rect 230620 204134 230940 204218
rect 230620 203898 230662 204134
rect 230898 203898 230940 204134
rect 230620 203866 230940 203898
rect 238462 204454 238782 204486
rect 238462 204218 238504 204454
rect 238740 204218 238782 204454
rect 238462 204134 238782 204218
rect 238462 203898 238504 204134
rect 238740 203898 238782 204134
rect 238462 203866 238782 203898
rect 246304 204454 246624 204486
rect 246304 204218 246346 204454
rect 246582 204218 246624 204454
rect 246304 204134 246624 204218
rect 246304 203898 246346 204134
rect 246582 203898 246624 204134
rect 246304 203866 246624 203898
rect 256910 204454 257230 204486
rect 256910 204218 256952 204454
rect 257188 204218 257230 204454
rect 256910 204134 257230 204218
rect 256910 203898 256952 204134
rect 257188 203898 257230 204134
rect 256910 203866 257230 203898
rect 264752 204454 265072 204486
rect 264752 204218 264794 204454
rect 265030 204218 265072 204454
rect 264752 204134 265072 204218
rect 264752 203898 264794 204134
rect 265030 203898 265072 204134
rect 264752 203866 265072 203898
rect 272594 204454 272914 204486
rect 272594 204218 272636 204454
rect 272872 204218 272914 204454
rect 272594 204134 272914 204218
rect 272594 203898 272636 204134
rect 272872 203898 272914 204134
rect 272594 203866 272914 203898
rect 280436 204454 280756 204486
rect 280436 204218 280478 204454
rect 280714 204218 280756 204454
rect 280436 204134 280756 204218
rect 280436 203898 280478 204134
rect 280714 203898 280756 204134
rect 280436 203866 280756 203898
rect 14065 198174 14385 198206
rect 14065 197938 14107 198174
rect 14343 197938 14385 198174
rect 14065 197854 14385 197938
rect 14065 197618 14107 197854
rect 14343 197618 14385 197854
rect 14065 197586 14385 197618
rect 21907 198174 22227 198206
rect 21907 197938 21949 198174
rect 22185 197938 22227 198174
rect 21907 197854 22227 197938
rect 21907 197618 21949 197854
rect 22185 197618 22227 197854
rect 21907 197586 22227 197618
rect 29749 198174 30069 198206
rect 29749 197938 29791 198174
rect 30027 197938 30069 198174
rect 29749 197854 30069 197938
rect 29749 197618 29791 197854
rect 30027 197618 30069 197854
rect 29749 197586 30069 197618
rect 37591 198174 37911 198206
rect 37591 197938 37633 198174
rect 37869 197938 37911 198174
rect 37591 197854 37911 197938
rect 37591 197618 37633 197854
rect 37869 197618 37911 197854
rect 37591 197586 37911 197618
rect 48197 198174 48517 198206
rect 48197 197938 48239 198174
rect 48475 197938 48517 198174
rect 48197 197854 48517 197938
rect 48197 197618 48239 197854
rect 48475 197618 48517 197854
rect 48197 197586 48517 197618
rect 56039 198174 56359 198206
rect 56039 197938 56081 198174
rect 56317 197938 56359 198174
rect 56039 197854 56359 197938
rect 56039 197618 56081 197854
rect 56317 197618 56359 197854
rect 56039 197586 56359 197618
rect 63881 198174 64201 198206
rect 63881 197938 63923 198174
rect 64159 197938 64201 198174
rect 63881 197854 64201 197938
rect 63881 197618 63923 197854
rect 64159 197618 64201 197854
rect 63881 197586 64201 197618
rect 71723 198174 72043 198206
rect 71723 197938 71765 198174
rect 72001 197938 72043 198174
rect 71723 197854 72043 197938
rect 71723 197618 71765 197854
rect 72001 197618 72043 197854
rect 71723 197586 72043 197618
rect 82329 198174 82649 198206
rect 82329 197938 82371 198174
rect 82607 197938 82649 198174
rect 82329 197854 82649 197938
rect 82329 197618 82371 197854
rect 82607 197618 82649 197854
rect 82329 197586 82649 197618
rect 90171 198174 90491 198206
rect 90171 197938 90213 198174
rect 90449 197938 90491 198174
rect 90171 197854 90491 197938
rect 90171 197618 90213 197854
rect 90449 197618 90491 197854
rect 90171 197586 90491 197618
rect 98013 198174 98333 198206
rect 98013 197938 98055 198174
rect 98291 197938 98333 198174
rect 98013 197854 98333 197938
rect 98013 197618 98055 197854
rect 98291 197618 98333 197854
rect 98013 197586 98333 197618
rect 105855 198174 106175 198206
rect 105855 197938 105897 198174
rect 106133 197938 106175 198174
rect 105855 197854 106175 197938
rect 105855 197618 105897 197854
rect 106133 197618 106175 197854
rect 105855 197586 106175 197618
rect 116461 198174 116781 198206
rect 116461 197938 116503 198174
rect 116739 197938 116781 198174
rect 116461 197854 116781 197938
rect 116461 197618 116503 197854
rect 116739 197618 116781 197854
rect 116461 197586 116781 197618
rect 124303 198174 124623 198206
rect 124303 197938 124345 198174
rect 124581 197938 124623 198174
rect 124303 197854 124623 197938
rect 124303 197618 124345 197854
rect 124581 197618 124623 197854
rect 124303 197586 124623 197618
rect 132145 198174 132465 198206
rect 132145 197938 132187 198174
rect 132423 197938 132465 198174
rect 132145 197854 132465 197938
rect 132145 197618 132187 197854
rect 132423 197618 132465 197854
rect 132145 197586 132465 197618
rect 139987 198174 140307 198206
rect 139987 197938 140029 198174
rect 140265 197938 140307 198174
rect 139987 197854 140307 197938
rect 139987 197618 140029 197854
rect 140265 197618 140307 197854
rect 139987 197586 140307 197618
rect 150593 198174 150913 198206
rect 150593 197938 150635 198174
rect 150871 197938 150913 198174
rect 150593 197854 150913 197938
rect 150593 197618 150635 197854
rect 150871 197618 150913 197854
rect 150593 197586 150913 197618
rect 158435 198174 158755 198206
rect 158435 197938 158477 198174
rect 158713 197938 158755 198174
rect 158435 197854 158755 197938
rect 158435 197618 158477 197854
rect 158713 197618 158755 197854
rect 158435 197586 158755 197618
rect 166277 198174 166597 198206
rect 166277 197938 166319 198174
rect 166555 197938 166597 198174
rect 166277 197854 166597 197938
rect 166277 197618 166319 197854
rect 166555 197618 166597 197854
rect 166277 197586 166597 197618
rect 174119 198174 174439 198206
rect 174119 197938 174161 198174
rect 174397 197938 174439 198174
rect 174119 197854 174439 197938
rect 174119 197618 174161 197854
rect 174397 197618 174439 197854
rect 174119 197586 174439 197618
rect 184725 198174 185045 198206
rect 184725 197938 184767 198174
rect 185003 197938 185045 198174
rect 184725 197854 185045 197938
rect 184725 197618 184767 197854
rect 185003 197618 185045 197854
rect 184725 197586 185045 197618
rect 192567 198174 192887 198206
rect 192567 197938 192609 198174
rect 192845 197938 192887 198174
rect 192567 197854 192887 197938
rect 192567 197618 192609 197854
rect 192845 197618 192887 197854
rect 192567 197586 192887 197618
rect 200409 198174 200729 198206
rect 200409 197938 200451 198174
rect 200687 197938 200729 198174
rect 200409 197854 200729 197938
rect 200409 197618 200451 197854
rect 200687 197618 200729 197854
rect 200409 197586 200729 197618
rect 208251 198174 208571 198206
rect 208251 197938 208293 198174
rect 208529 197938 208571 198174
rect 208251 197854 208571 197938
rect 208251 197618 208293 197854
rect 208529 197618 208571 197854
rect 208251 197586 208571 197618
rect 218857 198174 219177 198206
rect 218857 197938 218899 198174
rect 219135 197938 219177 198174
rect 218857 197854 219177 197938
rect 218857 197618 218899 197854
rect 219135 197618 219177 197854
rect 218857 197586 219177 197618
rect 226699 198174 227019 198206
rect 226699 197938 226741 198174
rect 226977 197938 227019 198174
rect 226699 197854 227019 197938
rect 226699 197618 226741 197854
rect 226977 197618 227019 197854
rect 226699 197586 227019 197618
rect 234541 198174 234861 198206
rect 234541 197938 234583 198174
rect 234819 197938 234861 198174
rect 234541 197854 234861 197938
rect 234541 197618 234583 197854
rect 234819 197618 234861 197854
rect 234541 197586 234861 197618
rect 242383 198174 242703 198206
rect 242383 197938 242425 198174
rect 242661 197938 242703 198174
rect 242383 197854 242703 197938
rect 242383 197618 242425 197854
rect 242661 197618 242703 197854
rect 242383 197586 242703 197618
rect 252989 198174 253309 198206
rect 252989 197938 253031 198174
rect 253267 197938 253309 198174
rect 252989 197854 253309 197938
rect 252989 197618 253031 197854
rect 253267 197618 253309 197854
rect 252989 197586 253309 197618
rect 260831 198174 261151 198206
rect 260831 197938 260873 198174
rect 261109 197938 261151 198174
rect 260831 197854 261151 197938
rect 260831 197618 260873 197854
rect 261109 197618 261151 197854
rect 260831 197586 261151 197618
rect 268673 198174 268993 198206
rect 268673 197938 268715 198174
rect 268951 197938 268993 198174
rect 268673 197854 268993 197938
rect 268673 197618 268715 197854
rect 268951 197618 268993 197854
rect 268673 197586 268993 197618
rect 276515 198174 276835 198206
rect 276515 197938 276557 198174
rect 276793 197938 276835 198174
rect 276515 197854 276835 197938
rect 276515 197618 276557 197854
rect 276793 197618 276835 197854
rect 276515 197586 276835 197618
rect 10179 194580 10245 194581
rect 10179 194516 10180 194580
rect 10244 194516 10245 194580
rect 10179 194515 10245 194516
rect 17986 194454 18306 194486
rect 17986 194218 18028 194454
rect 18264 194218 18306 194454
rect 17986 194134 18306 194218
rect 17986 193898 18028 194134
rect 18264 193898 18306 194134
rect 17986 193866 18306 193898
rect 25828 194454 26148 194486
rect 25828 194218 25870 194454
rect 26106 194218 26148 194454
rect 25828 194134 26148 194218
rect 25828 193898 25870 194134
rect 26106 193898 26148 194134
rect 25828 193866 26148 193898
rect 33670 194454 33990 194486
rect 33670 194218 33712 194454
rect 33948 194218 33990 194454
rect 33670 194134 33990 194218
rect 33670 193898 33712 194134
rect 33948 193898 33990 194134
rect 33670 193866 33990 193898
rect 41512 194454 41832 194486
rect 41512 194218 41554 194454
rect 41790 194218 41832 194454
rect 41512 194134 41832 194218
rect 41512 193898 41554 194134
rect 41790 193898 41832 194134
rect 41512 193866 41832 193898
rect 52118 194454 52438 194486
rect 52118 194218 52160 194454
rect 52396 194218 52438 194454
rect 52118 194134 52438 194218
rect 52118 193898 52160 194134
rect 52396 193898 52438 194134
rect 52118 193866 52438 193898
rect 59960 194454 60280 194486
rect 59960 194218 60002 194454
rect 60238 194218 60280 194454
rect 59960 194134 60280 194218
rect 59960 193898 60002 194134
rect 60238 193898 60280 194134
rect 59960 193866 60280 193898
rect 67802 194454 68122 194486
rect 67802 194218 67844 194454
rect 68080 194218 68122 194454
rect 67802 194134 68122 194218
rect 67802 193898 67844 194134
rect 68080 193898 68122 194134
rect 67802 193866 68122 193898
rect 75644 194454 75964 194486
rect 75644 194218 75686 194454
rect 75922 194218 75964 194454
rect 75644 194134 75964 194218
rect 75644 193898 75686 194134
rect 75922 193898 75964 194134
rect 75644 193866 75964 193898
rect 86250 194454 86570 194486
rect 86250 194218 86292 194454
rect 86528 194218 86570 194454
rect 86250 194134 86570 194218
rect 86250 193898 86292 194134
rect 86528 193898 86570 194134
rect 86250 193866 86570 193898
rect 94092 194454 94412 194486
rect 94092 194218 94134 194454
rect 94370 194218 94412 194454
rect 94092 194134 94412 194218
rect 94092 193898 94134 194134
rect 94370 193898 94412 194134
rect 94092 193866 94412 193898
rect 101934 194454 102254 194486
rect 101934 194218 101976 194454
rect 102212 194218 102254 194454
rect 101934 194134 102254 194218
rect 101934 193898 101976 194134
rect 102212 193898 102254 194134
rect 101934 193866 102254 193898
rect 109776 194454 110096 194486
rect 109776 194218 109818 194454
rect 110054 194218 110096 194454
rect 109776 194134 110096 194218
rect 109776 193898 109818 194134
rect 110054 193898 110096 194134
rect 109776 193866 110096 193898
rect 120382 194454 120702 194486
rect 120382 194218 120424 194454
rect 120660 194218 120702 194454
rect 120382 194134 120702 194218
rect 120382 193898 120424 194134
rect 120660 193898 120702 194134
rect 120382 193866 120702 193898
rect 128224 194454 128544 194486
rect 128224 194218 128266 194454
rect 128502 194218 128544 194454
rect 128224 194134 128544 194218
rect 128224 193898 128266 194134
rect 128502 193898 128544 194134
rect 128224 193866 128544 193898
rect 136066 194454 136386 194486
rect 136066 194218 136108 194454
rect 136344 194218 136386 194454
rect 136066 194134 136386 194218
rect 136066 193898 136108 194134
rect 136344 193898 136386 194134
rect 136066 193866 136386 193898
rect 143908 194454 144228 194486
rect 143908 194218 143950 194454
rect 144186 194218 144228 194454
rect 143908 194134 144228 194218
rect 143908 193898 143950 194134
rect 144186 193898 144228 194134
rect 143908 193866 144228 193898
rect 154514 194454 154834 194486
rect 154514 194218 154556 194454
rect 154792 194218 154834 194454
rect 154514 194134 154834 194218
rect 154514 193898 154556 194134
rect 154792 193898 154834 194134
rect 154514 193866 154834 193898
rect 162356 194454 162676 194486
rect 162356 194218 162398 194454
rect 162634 194218 162676 194454
rect 162356 194134 162676 194218
rect 162356 193898 162398 194134
rect 162634 193898 162676 194134
rect 162356 193866 162676 193898
rect 170198 194454 170518 194486
rect 170198 194218 170240 194454
rect 170476 194218 170518 194454
rect 170198 194134 170518 194218
rect 170198 193898 170240 194134
rect 170476 193898 170518 194134
rect 170198 193866 170518 193898
rect 178040 194454 178360 194486
rect 178040 194218 178082 194454
rect 178318 194218 178360 194454
rect 178040 194134 178360 194218
rect 178040 193898 178082 194134
rect 178318 193898 178360 194134
rect 178040 193866 178360 193898
rect 188646 194454 188966 194486
rect 188646 194218 188688 194454
rect 188924 194218 188966 194454
rect 188646 194134 188966 194218
rect 188646 193898 188688 194134
rect 188924 193898 188966 194134
rect 188646 193866 188966 193898
rect 196488 194454 196808 194486
rect 196488 194218 196530 194454
rect 196766 194218 196808 194454
rect 196488 194134 196808 194218
rect 196488 193898 196530 194134
rect 196766 193898 196808 194134
rect 196488 193866 196808 193898
rect 204330 194454 204650 194486
rect 204330 194218 204372 194454
rect 204608 194218 204650 194454
rect 204330 194134 204650 194218
rect 204330 193898 204372 194134
rect 204608 193898 204650 194134
rect 204330 193866 204650 193898
rect 212172 194454 212492 194486
rect 212172 194218 212214 194454
rect 212450 194218 212492 194454
rect 212172 194134 212492 194218
rect 212172 193898 212214 194134
rect 212450 193898 212492 194134
rect 212172 193866 212492 193898
rect 222778 194454 223098 194486
rect 222778 194218 222820 194454
rect 223056 194218 223098 194454
rect 222778 194134 223098 194218
rect 222778 193898 222820 194134
rect 223056 193898 223098 194134
rect 222778 193866 223098 193898
rect 230620 194454 230940 194486
rect 230620 194218 230662 194454
rect 230898 194218 230940 194454
rect 230620 194134 230940 194218
rect 230620 193898 230662 194134
rect 230898 193898 230940 194134
rect 230620 193866 230940 193898
rect 238462 194454 238782 194486
rect 238462 194218 238504 194454
rect 238740 194218 238782 194454
rect 238462 194134 238782 194218
rect 238462 193898 238504 194134
rect 238740 193898 238782 194134
rect 238462 193866 238782 193898
rect 246304 194454 246624 194486
rect 246304 194218 246346 194454
rect 246582 194218 246624 194454
rect 246304 194134 246624 194218
rect 246304 193898 246346 194134
rect 246582 193898 246624 194134
rect 246304 193866 246624 193898
rect 256910 194454 257230 194486
rect 256910 194218 256952 194454
rect 257188 194218 257230 194454
rect 256910 194134 257230 194218
rect 256910 193898 256952 194134
rect 257188 193898 257230 194134
rect 256910 193866 257230 193898
rect 264752 194454 265072 194486
rect 264752 194218 264794 194454
rect 265030 194218 265072 194454
rect 264752 194134 265072 194218
rect 264752 193898 264794 194134
rect 265030 193898 265072 194134
rect 264752 193866 265072 193898
rect 272594 194454 272914 194486
rect 272594 194218 272636 194454
rect 272872 194218 272914 194454
rect 272594 194134 272914 194218
rect 272594 193898 272636 194134
rect 272872 193898 272914 194134
rect 272594 193866 272914 193898
rect 280436 194454 280756 194486
rect 280436 194218 280478 194454
rect 280714 194218 280756 194454
rect 280436 194134 280756 194218
rect 280436 193898 280478 194134
rect 280714 193898 280756 194134
rect 280436 193866 280756 193898
rect 281027 191996 281093 191997
rect 281027 191932 281028 191996
rect 281092 191932 281093 191996
rect 281027 191931 281093 191932
rect 10734 190400 10794 191420
rect 11470 190400 11530 191080
rect 12206 190400 12266 191080
rect 12942 190400 13002 191420
rect 13678 190400 13738 191080
rect 14414 190400 14474 191080
rect 15150 190400 15210 191080
rect 15886 190400 15946 191080
rect 16622 190400 16682 191080
rect 17358 190400 17418 191080
rect 18094 190400 18154 191080
rect 18830 190400 18890 191420
rect 19566 190400 19626 191420
rect 20302 190400 20362 191080
rect 21038 190400 21098 191420
rect 21774 190400 21834 191080
rect 22510 190400 22570 191420
rect 23246 190400 23306 191080
rect 23982 190400 24042 191080
rect 24718 190400 24778 191420
rect 25454 190400 25514 191420
rect 26190 190400 26250 191080
rect 26926 190400 26986 191420
rect 27662 190400 27722 191080
rect 28398 190060 28458 191080
rect 29134 190060 29194 191080
rect 29870 190400 29930 191080
rect 30606 190400 30666 191080
rect 31342 190400 31402 191080
rect 32078 190060 32138 191080
rect 32814 190060 32874 191080
rect 33550 190060 33610 191080
rect 34286 190060 34346 191044
rect 35022 190400 35082 191044
rect 35758 190060 35818 191044
rect 36494 190060 36554 191044
rect 37230 190060 37290 191044
rect 37966 190400 38026 191044
rect 38702 190060 38762 191044
rect 39438 190060 39498 191420
rect 40174 190060 40234 191420
rect 40910 190400 40970 191080
rect 41646 190400 41706 191044
rect 44866 190770 44926 191420
rect 44774 190710 44926 190770
rect 44774 190470 44834 190710
rect 44774 190410 44926 190470
rect 44866 190400 44926 190410
rect 45602 190400 45662 191080
rect 46338 190400 46398 191080
rect 47074 190770 47134 191420
rect 47074 190710 47226 190770
rect 47166 190470 47226 190710
rect 47074 190410 47226 190470
rect 47074 190400 47134 190410
rect 47810 190400 47870 191080
rect 48546 190400 48606 191080
rect 49282 190400 49342 191080
rect 50018 190400 50078 191080
rect 50754 190400 50814 191080
rect 51490 190400 51550 191080
rect 52226 190400 52286 191080
rect 52962 190400 53022 191420
rect 53698 190400 53758 191420
rect 54434 190400 54494 191080
rect 55170 190400 55230 191420
rect 55906 190400 55966 191080
rect 56642 190400 56702 191420
rect 57378 190400 57438 191080
rect 58114 190400 58174 191080
rect 58850 190400 58910 191420
rect 59586 190400 59646 191420
rect 60322 190400 60382 191080
rect 61058 190400 61118 191420
rect 61794 190400 61854 191080
rect 62530 190400 62590 191080
rect 63266 190400 63326 191080
rect 64002 190400 64062 191080
rect 64738 190400 64798 191080
rect 65474 190400 65534 191080
rect 66210 190400 66270 191080
rect 66946 190400 67006 191080
rect 67682 190400 67742 191080
rect 68418 190400 68478 191044
rect 69154 190400 69214 191044
rect 69890 190400 69950 191044
rect 70626 190400 70686 191044
rect 71362 190400 71422 191044
rect 72098 190400 72158 191044
rect 72834 190400 72894 191044
rect 73570 190400 73630 191420
rect 74306 190400 74366 191420
rect 75042 190400 75102 191080
rect 75778 190400 75838 191044
rect 78998 190060 79058 191420
rect 79734 190400 79794 191080
rect 80470 190400 80530 191080
rect 81206 190400 81266 191420
rect 81942 190400 82002 191080
rect 82678 190060 82738 191080
rect 83414 190400 83474 191080
rect 84150 190060 84210 191080
rect 84886 190400 84946 191080
rect 85622 190400 85682 191080
rect 86358 190400 86418 191080
rect 87094 190400 87154 191420
rect 87830 190060 87890 191420
rect 88566 190400 88626 191080
rect 89302 190060 89362 191420
rect 90038 190400 90098 191080
rect 90774 190400 90834 191420
rect 91510 190400 91570 191080
rect 92246 190400 92306 191080
rect 92982 190400 93042 191420
rect 93718 190400 93778 191420
rect 94454 190400 94514 191080
rect 95190 190400 95250 191420
rect 95926 190400 95986 191080
rect 96662 190060 96722 191080
rect 97398 190400 97458 191080
rect 98134 190060 98194 191080
rect 98870 190400 98930 191080
rect 99606 190060 99666 191080
rect 100342 190060 100402 191080
rect 101078 190060 101138 191080
rect 101814 190060 101874 191080
rect 102550 190400 102610 191044
rect 103286 190060 103346 191044
rect 104022 190060 104082 191044
rect 104758 190400 104818 191044
rect 105494 190400 105554 191044
rect 106230 190060 106290 191044
rect 106966 190400 107026 191044
rect 107702 190060 107762 191420
rect 108438 190060 108498 191420
rect 109174 190060 109234 191080
rect 109910 190400 109970 191044
rect 113130 190770 113190 191420
rect 113130 190710 113282 190770
rect 113222 190470 113282 190710
rect 113130 190410 113282 190470
rect 113130 190400 113190 190410
rect 113866 190400 113926 191080
rect 114602 190400 114662 191080
rect 115338 190770 115398 191420
rect 115338 190710 115490 190770
rect 115430 190470 115490 190710
rect 115338 190410 115490 190470
rect 115338 190400 115398 190410
rect 116074 190400 116134 191080
rect 116810 190400 116870 191080
rect 117546 190400 117606 191080
rect 118282 190400 118342 191080
rect 119018 190400 119078 191080
rect 119754 190400 119814 191080
rect 120490 190400 120550 191080
rect 121226 190400 121286 191420
rect 121962 190400 122022 191420
rect 122698 190400 122758 191080
rect 123434 190400 123494 191420
rect 124170 190400 124230 191080
rect 124906 190400 124966 191420
rect 125642 190400 125702 191080
rect 126378 190400 126438 191080
rect 127114 190400 127174 191420
rect 127850 190400 127910 191420
rect 128586 190400 128646 191080
rect 129322 190400 129382 191420
rect 130058 190400 130118 191080
rect 130794 190400 130854 191080
rect 131530 190400 131590 191080
rect 132266 190400 132326 191080
rect 133002 190400 133062 191080
rect 133738 190400 133798 191080
rect 134474 190400 134534 191080
rect 135210 190400 135270 191080
rect 135946 190400 136006 191080
rect 136682 190400 136742 191044
rect 137418 190400 137478 191044
rect 138154 190400 138214 191044
rect 138890 190400 138950 191044
rect 139626 190400 139686 191044
rect 140362 190400 140422 191044
rect 141098 190400 141158 191044
rect 141834 190770 141894 191420
rect 142570 190770 142630 191420
rect 141834 190710 141986 190770
rect 141926 190470 141986 190710
rect 141834 190410 141986 190470
rect 142478 190710 142630 190770
rect 142478 190470 142538 190710
rect 142478 190410 142630 190470
rect 141834 190400 141894 190410
rect 142570 190400 142630 190410
rect 143306 190400 143366 191080
rect 144042 190400 144102 191044
rect 147262 190400 147322 191420
rect 147998 190400 148058 191080
rect 148734 190400 148794 191080
rect 149470 190400 149530 191420
rect 150206 190400 150266 191080
rect 150942 190400 151002 191080
rect 151678 190400 151738 191080
rect 152414 190400 152474 191080
rect 153150 190400 153210 191080
rect 153886 190400 153946 191080
rect 154622 190400 154682 191080
rect 155358 190400 155418 191420
rect 156094 190400 156154 191420
rect 156830 190400 156890 191080
rect 157566 190400 157626 191420
rect 158302 190400 158362 191080
rect 159038 190400 159098 191420
rect 159774 190400 159834 191080
rect 160510 190400 160570 191080
rect 161246 190400 161306 191420
rect 161982 190400 162042 191420
rect 162718 190400 162778 191080
rect 163454 190400 163514 191420
rect 164190 190400 164250 191080
rect 164926 190400 164986 191080
rect 165662 190400 165722 191080
rect 166398 190400 166458 191080
rect 167134 190400 167194 191080
rect 167870 190400 167930 191080
rect 168606 190400 168666 191080
rect 169342 190060 169402 191080
rect 170078 190060 170138 191080
rect 170814 190060 170874 191044
rect 171550 190060 171610 191044
rect 172286 190060 172346 191044
rect 173022 190400 173082 191044
rect 173758 190060 173818 191044
rect 174494 190060 174554 191044
rect 175230 190060 175290 191044
rect 175966 190060 176026 191420
rect 176702 190060 176762 191420
rect 177438 190060 177498 191080
rect 178174 190400 178234 191044
rect 181394 190770 181454 191420
rect 181394 190710 181546 190770
rect 181486 190470 181546 190710
rect 181394 190410 181546 190470
rect 181394 190400 181454 190410
rect 182130 190400 182190 191080
rect 182866 190400 182926 191080
rect 183602 190770 183662 191420
rect 183602 190710 183754 190770
rect 183694 190470 183754 190710
rect 183602 190410 183754 190470
rect 183602 190400 183662 190410
rect 184338 190400 184398 191080
rect 185074 190400 185134 191080
rect 185810 190400 185870 191080
rect 186546 190400 186606 191080
rect 187282 190400 187342 191080
rect 188018 190400 188078 191080
rect 188754 190400 188814 191080
rect 189490 190400 189550 191420
rect 190226 190400 190286 191420
rect 190962 190400 191022 191080
rect 191698 190400 191758 191420
rect 192434 190400 192494 191080
rect 193170 190400 193230 191420
rect 193906 190400 193966 191080
rect 194642 190400 194702 191080
rect 195378 190400 195438 191420
rect 196114 190400 196174 191420
rect 196850 190400 196910 191080
rect 197586 190400 197646 191420
rect 198322 190400 198382 191080
rect 199058 190400 199118 191080
rect 199794 190400 199854 191080
rect 200530 190400 200590 191080
rect 201266 190400 201326 191080
rect 202002 190400 202062 191080
rect 202738 190400 202798 191080
rect 203474 190400 203534 191080
rect 204210 190400 204270 191080
rect 204946 190400 205006 191044
rect 205682 190400 205742 191044
rect 206418 190400 206478 191044
rect 207154 190400 207214 191044
rect 207890 190400 207950 191044
rect 208626 190400 208686 191044
rect 209362 190400 209422 191044
rect 210098 190400 210158 191420
rect 210834 190400 210894 191420
rect 211570 190400 211630 191080
rect 212306 190400 212366 191044
rect 215526 190400 215586 191420
rect 216262 190400 216322 191080
rect 216998 190400 217058 191080
rect 217734 190400 217794 191420
rect 218470 190400 218530 191080
rect 219206 190400 219266 191080
rect 219942 190400 220002 191080
rect 220678 190400 220738 191080
rect 221414 190060 221474 191080
rect 222150 190400 222210 191080
rect 222886 190400 222946 191080
rect 223622 190400 223682 191420
rect 224358 190400 224418 191420
rect 225094 190400 225154 191080
rect 225830 190400 225890 191420
rect 226566 190400 226626 191080
rect 227302 190400 227362 191420
rect 228038 190400 228098 191080
rect 228774 190400 228834 191080
rect 229510 190400 229570 191420
rect 230246 190400 230306 191420
rect 230982 190400 231042 191080
rect 231718 190400 231778 191420
rect 232454 190400 232514 191080
rect 233190 190400 233250 191080
rect 233926 190060 233986 191080
rect 234662 190400 234722 191080
rect 235398 190060 235458 191080
rect 236134 190060 236194 191080
rect 236870 190060 236930 191080
rect 237606 190400 237666 191080
rect 238342 190060 238402 191080
rect 239078 190400 239138 191044
rect 239814 190060 239874 191044
rect 240550 190400 240610 191044
rect 241286 190060 241346 191044
rect 242022 190060 242082 191044
rect 242758 190400 242818 191044
rect 243494 190400 243554 191044
rect 244230 190400 244290 191420
rect 244966 190400 245026 191420
rect 245702 190060 245762 191080
rect 246438 190400 246498 191044
rect 249658 190770 249718 191420
rect 249658 190710 249810 190770
rect 249750 190470 249810 190710
rect 249658 190410 249810 190470
rect 249658 190400 249718 190410
rect 250394 190400 250454 191080
rect 251130 190400 251190 191080
rect 251866 190770 251926 191420
rect 251866 190710 252018 190770
rect 251958 190470 252018 190710
rect 251866 190410 252018 190470
rect 251866 190400 251926 190410
rect 252602 190400 252662 191080
rect 253338 190400 253398 191080
rect 254074 190400 254134 191080
rect 254810 190400 254870 191080
rect 255546 190400 255606 191080
rect 256282 190400 256342 191080
rect 257018 190400 257078 191080
rect 257754 190400 257814 191420
rect 258490 190400 258550 191420
rect 259226 190400 259286 191080
rect 259962 190400 260022 191420
rect 260698 190400 260758 191080
rect 261434 190400 261494 191420
rect 262170 190400 262230 191080
rect 262906 190400 262966 191080
rect 263642 190400 263702 191420
rect 264378 190400 264438 191420
rect 265114 190400 265174 191080
rect 265850 190400 265910 191420
rect 266586 190400 266646 191080
rect 267322 190400 267382 191080
rect 268058 190400 268118 191080
rect 268794 190400 268854 191080
rect 269530 190400 269590 191080
rect 270266 190400 270326 191080
rect 271002 190400 271062 191080
rect 271738 190400 271798 191080
rect 272474 190400 272534 191080
rect 273210 190400 273270 191044
rect 273946 190400 274006 191044
rect 274682 190400 274742 191044
rect 275418 190400 275478 191044
rect 276154 190400 276214 191044
rect 276890 190400 276950 191044
rect 277626 190400 277686 191044
rect 278362 190400 278422 191420
rect 279098 190400 279158 191420
rect 279834 190400 279894 191080
rect 280570 190400 280630 191044
rect 9627 189140 9693 189141
rect 9627 189076 9628 189140
rect 9692 189076 9693 189140
rect 9627 189075 9693 189076
rect 43942 188174 44262 188206
rect 43942 187938 43984 188174
rect 44220 187938 44262 188174
rect 43942 187854 44262 187938
rect 43942 187618 43984 187854
rect 44220 187618 44262 187854
rect 43942 187586 44262 187618
rect 111539 188174 111859 188206
rect 111539 187938 111581 188174
rect 111817 187938 111859 188174
rect 111539 187854 111859 187938
rect 111539 187618 111581 187854
rect 111817 187618 111859 187854
rect 111539 187586 111859 187618
rect 179136 188174 179456 188206
rect 179136 187938 179178 188174
rect 179414 187938 179456 188174
rect 179136 187854 179456 187938
rect 179136 187618 179178 187854
rect 179414 187618 179456 187854
rect 179136 187586 179456 187618
rect 246733 188174 247053 188206
rect 246733 187938 246775 188174
rect 247011 187938 247053 188174
rect 246733 187854 247053 187938
rect 246733 187618 246775 187854
rect 247011 187618 247053 187854
rect 246733 187586 247053 187618
rect 77740 184454 78060 184486
rect 77740 184218 77782 184454
rect 78018 184218 78060 184454
rect 77740 184134 78060 184218
rect 77740 183898 77782 184134
rect 78018 183898 78060 184134
rect 77740 183866 78060 183898
rect 145337 184454 145657 184486
rect 145337 184218 145379 184454
rect 145615 184218 145657 184454
rect 145337 184134 145657 184218
rect 145337 183898 145379 184134
rect 145615 183898 145657 184134
rect 145337 183866 145657 183898
rect 212934 184454 213254 184486
rect 212934 184218 212976 184454
rect 213212 184218 213254 184454
rect 212934 184134 213254 184218
rect 212934 183898 212976 184134
rect 213212 183898 213254 184134
rect 212934 183866 213254 183898
rect 280531 184454 280851 184486
rect 280531 184218 280573 184454
rect 280809 184218 280851 184454
rect 280531 184134 280851 184218
rect 280531 183898 280573 184134
rect 280809 183898 280851 184134
rect 280531 183866 280851 183898
rect 281030 183701 281090 191931
rect 282134 191589 282194 566883
rect 282867 192268 282933 192269
rect 282867 192204 282868 192268
rect 282932 192204 282933 192268
rect 282867 192203 282933 192204
rect 282870 192130 282930 192203
rect 282686 192070 282930 192130
rect 282131 191588 282197 191589
rect 282131 191524 282132 191588
rect 282196 191524 282197 191588
rect 282131 191523 282197 191524
rect 282686 190090 282746 192070
rect 283971 190636 284037 190637
rect 283971 190572 283972 190636
rect 284036 190572 284037 190636
rect 283971 190571 284037 190572
rect 282502 190030 282746 190090
rect 282315 188324 282381 188325
rect 282315 188260 282316 188324
rect 282380 188260 282381 188324
rect 282315 188259 282381 188260
rect 282318 186693 282378 188259
rect 282502 187373 282562 190030
rect 282683 189684 282749 189685
rect 282683 189620 282684 189684
rect 282748 189620 282749 189684
rect 282683 189619 282749 189620
rect 282499 187372 282565 187373
rect 282499 187308 282500 187372
rect 282564 187308 282565 187372
rect 282499 187307 282565 187308
rect 282315 186692 282381 186693
rect 282315 186628 282316 186692
rect 282380 186628 282381 186692
rect 282315 186627 282381 186628
rect 282686 184789 282746 189619
rect 283787 189548 283853 189549
rect 283787 189484 283788 189548
rect 283852 189484 283853 189548
rect 283787 189483 283853 189484
rect 283790 186149 283850 189483
rect 283787 186148 283853 186149
rect 283787 186084 283788 186148
rect 283852 186084 283853 186148
rect 283787 186083 283853 186084
rect 283974 185877 284034 190571
rect 284155 189276 284221 189277
rect 284155 189212 284156 189276
rect 284220 189212 284221 189276
rect 284155 189211 284221 189212
rect 284158 186013 284218 189211
rect 284155 186012 284221 186013
rect 284155 185948 284156 186012
rect 284220 185948 284221 186012
rect 284155 185947 284221 185948
rect 283971 185876 284037 185877
rect 283971 185812 283972 185876
rect 284036 185812 284037 185876
rect 283971 185811 284037 185812
rect 282867 185740 282933 185741
rect 282867 185676 282868 185740
rect 282932 185676 282933 185740
rect 282867 185675 282933 185676
rect 282683 184788 282749 184789
rect 282683 184724 282684 184788
rect 282748 184724 282749 184788
rect 282683 184723 282749 184724
rect 282870 184517 282930 185675
rect 282867 184516 282933 184517
rect 282867 184452 282868 184516
rect 282932 184452 282933 184516
rect 282867 184451 282933 184452
rect 284342 183701 284402 699755
rect 585310 698174 585930 704282
rect 585310 697938 585342 698174
rect 585578 697938 585662 698174
rect 585898 697938 585930 698174
rect 585310 697854 585930 697938
rect 585310 697618 585342 697854
rect 585578 697618 585662 697854
rect 585898 697618 585930 697854
rect 585310 688174 585930 697618
rect 585310 687938 585342 688174
rect 585578 687938 585662 688174
rect 585898 687938 585930 688174
rect 585310 687854 585930 687938
rect 585310 687618 585342 687854
rect 585578 687618 585662 687854
rect 585898 687618 585930 687854
rect 585310 678174 585930 687618
rect 585310 677938 585342 678174
rect 585578 677938 585662 678174
rect 585898 677938 585930 678174
rect 585310 677854 585930 677938
rect 585310 677618 585342 677854
rect 585578 677618 585662 677854
rect 585898 677618 585930 677854
rect 574691 670716 574757 670717
rect 574691 670652 574692 670716
rect 574756 670652 574757 670716
rect 574691 670651 574757 670652
rect 291147 658204 291213 658205
rect 291147 658140 291148 658204
rect 291212 658140 291213 658204
rect 291147 658139 291213 658140
rect 288387 606116 288453 606117
rect 288387 606052 288388 606116
rect 288452 606052 288453 606116
rect 288387 606051 288453 606052
rect 285627 214572 285693 214573
rect 285627 214508 285628 214572
rect 285692 214508 285693 214572
rect 285627 214507 285693 214508
rect 284523 192132 284589 192133
rect 284523 192068 284524 192132
rect 284588 192068 284589 192132
rect 284523 192067 284589 192068
rect 284526 184381 284586 192067
rect 285443 190364 285509 190365
rect 285443 190300 285444 190364
rect 285508 190300 285509 190364
rect 285443 190299 285509 190300
rect 285446 187509 285506 190299
rect 285443 187508 285509 187509
rect 285443 187444 285444 187508
rect 285508 187444 285509 187508
rect 285443 187443 285509 187444
rect 285446 184925 285506 187443
rect 285630 187373 285690 214507
rect 288203 210356 288269 210357
rect 288203 210292 288204 210356
rect 288268 210292 288269 210356
rect 288203 210291 288269 210292
rect 286179 191588 286245 191589
rect 286179 191524 286180 191588
rect 286244 191524 286245 191588
rect 286179 191523 286245 191524
rect 285627 187372 285693 187373
rect 285627 187308 285628 187372
rect 285692 187308 285693 187372
rect 285627 187307 285693 187308
rect 285443 184924 285509 184925
rect 285443 184860 285444 184924
rect 285508 184860 285509 184924
rect 285443 184859 285509 184860
rect 284523 184380 284589 184381
rect 284523 184316 284524 184380
rect 284588 184316 284589 184380
rect 284523 184315 284589 184316
rect 281027 183700 281093 183701
rect 281027 183636 281028 183700
rect 281092 183636 281093 183700
rect 281027 183635 281093 183636
rect 284339 183700 284405 183701
rect 284339 183636 284340 183700
rect 284404 183636 284405 183700
rect 284339 183635 284405 183636
rect 285995 182340 286061 182341
rect 285995 182276 285996 182340
rect 286060 182276 286061 182340
rect 285995 182275 286061 182276
rect 285259 182068 285325 182069
rect 285259 182004 285260 182068
rect 285324 182004 285325 182068
rect 285259 182003 285325 182004
rect 284891 181932 284957 181933
rect 284891 181868 284892 181932
rect 284956 181868 284957 181932
rect 284891 181867 284957 181868
rect 284523 181796 284589 181797
rect 284523 181732 284524 181796
rect 284588 181732 284589 181796
rect 284523 181731 284589 181732
rect 283051 181660 283117 181661
rect 283051 181596 283052 181660
rect 283116 181596 283117 181660
rect 283051 181595 283117 181596
rect 281579 181116 281645 181117
rect 281579 181052 281580 181116
rect 281644 181052 281645 181116
rect 281579 181051 281645 181052
rect 9443 178940 9509 178941
rect 9443 178876 9444 178940
rect 9508 178876 9509 178940
rect 9443 178875 9509 178876
rect 10734 178500 10794 179520
rect 11470 178840 11530 179520
rect 12206 178840 12266 179520
rect 12942 178500 13002 179520
rect 13678 178840 13738 179520
rect 14414 178840 14474 179520
rect 15150 178840 15210 179520
rect 15886 178840 15946 179520
rect 16622 178840 16682 179520
rect 17358 178840 17418 179520
rect 18094 178840 18154 179520
rect 18830 178500 18890 179520
rect 19566 178500 19626 179520
rect 20302 178840 20362 179520
rect 21038 178500 21098 179520
rect 21774 178840 21834 179520
rect 22510 178500 22570 179520
rect 23246 178840 23306 179520
rect 23982 178840 24042 179520
rect 24718 178500 24778 179520
rect 25454 178500 25514 179520
rect 26190 178840 26250 179520
rect 26926 178500 26986 179520
rect 27662 178840 27722 179520
rect 28398 178840 28458 179860
rect 29134 178840 29194 179860
rect 29870 178840 29930 179520
rect 30606 178840 30666 179520
rect 31342 178840 31402 179860
rect 32078 178840 32138 179860
rect 32814 178840 32874 179520
rect 33550 178840 33610 179860
rect 34286 178876 34346 179860
rect 35022 178876 35082 179520
rect 35758 178876 35818 179520
rect 36494 178876 36554 179520
rect 37230 178876 37290 179520
rect 37966 178876 38026 179520
rect 38702 178876 38762 179520
rect 39438 178500 39498 179520
rect 40174 178500 40234 179520
rect 40910 178840 40970 179520
rect 41646 178876 41706 179520
rect 43299 178940 43365 178941
rect 43299 178876 43300 178940
rect 43364 178876 43365 178940
rect 43299 178875 43365 178876
rect 14065 177879 14385 177936
rect 14065 177643 14107 177879
rect 14343 177643 14385 177879
rect 14065 177586 14385 177643
rect 21907 177879 22227 177936
rect 21907 177643 21949 177879
rect 22185 177643 22227 177879
rect 21907 177586 22227 177643
rect 29749 177879 30069 177936
rect 29749 177643 29791 177879
rect 30027 177643 30069 177879
rect 29749 177586 30069 177643
rect 37591 177879 37911 177936
rect 37591 177643 37633 177879
rect 37869 177643 37911 177879
rect 37591 177586 37911 177643
rect 10179 175268 10245 175269
rect 10179 175204 10180 175268
rect 10244 175204 10245 175268
rect 10179 175203 10245 175204
rect 10182 157453 10242 175203
rect 17986 174454 18306 174486
rect 17986 174218 18028 174454
rect 18264 174218 18306 174454
rect 17986 174134 18306 174218
rect 17986 173898 18028 174134
rect 18264 173898 18306 174134
rect 17986 173866 18306 173898
rect 25828 174454 26148 174486
rect 25828 174218 25870 174454
rect 26106 174218 26148 174454
rect 25828 174134 26148 174218
rect 25828 173898 25870 174134
rect 26106 173898 26148 174134
rect 25828 173866 26148 173898
rect 33670 174454 33990 174486
rect 33670 174218 33712 174454
rect 33948 174218 33990 174454
rect 33670 174134 33990 174218
rect 33670 173898 33712 174134
rect 33948 173898 33990 174134
rect 33670 173866 33990 173898
rect 41512 174454 41832 174486
rect 41512 174218 41554 174454
rect 41790 174218 41832 174454
rect 41512 174134 41832 174218
rect 41512 173898 41554 174134
rect 41790 173898 41832 174134
rect 41512 173866 41832 173898
rect 14065 168174 14385 168206
rect 14065 167938 14107 168174
rect 14343 167938 14385 168174
rect 14065 167854 14385 167938
rect 14065 167618 14107 167854
rect 14343 167618 14385 167854
rect 14065 167586 14385 167618
rect 21907 168174 22227 168206
rect 21907 167938 21949 168174
rect 22185 167938 22227 168174
rect 21907 167854 22227 167938
rect 21907 167618 21949 167854
rect 22185 167618 22227 167854
rect 21907 167586 22227 167618
rect 29749 168174 30069 168206
rect 29749 167938 29791 168174
rect 30027 167938 30069 168174
rect 29749 167854 30069 167938
rect 29749 167618 29791 167854
rect 30027 167618 30069 167854
rect 29749 167586 30069 167618
rect 37591 168174 37911 168206
rect 37591 167938 37633 168174
rect 37869 167938 37911 168174
rect 37591 167854 37911 167938
rect 37591 167618 37633 167854
rect 37869 167618 37911 167854
rect 37591 167586 37911 167618
rect 17986 164454 18306 164486
rect 17986 164218 18028 164454
rect 18264 164218 18306 164454
rect 17986 164134 18306 164218
rect 17986 163898 18028 164134
rect 18264 163898 18306 164134
rect 17986 163866 18306 163898
rect 25828 164454 26148 164486
rect 25828 164218 25870 164454
rect 26106 164218 26148 164454
rect 25828 164134 26148 164218
rect 25828 163898 25870 164134
rect 26106 163898 26148 164134
rect 25828 163866 26148 163898
rect 33670 164454 33990 164486
rect 33670 164218 33712 164454
rect 33948 164218 33990 164454
rect 33670 164134 33990 164218
rect 33670 163898 33712 164134
rect 33948 163898 33990 164134
rect 33670 163866 33990 163898
rect 41512 164454 41832 164486
rect 41512 164218 41554 164454
rect 41790 164218 41832 164454
rect 41512 164134 41832 164218
rect 41512 163898 41554 164134
rect 41790 163898 41832 164134
rect 41512 163866 41832 163898
rect 10179 157452 10245 157453
rect 10179 157388 10180 157452
rect 10244 157388 10245 157452
rect 10179 157387 10245 157388
rect 9075 73948 9141 73949
rect 9075 73884 9076 73948
rect 9140 73884 9141 73948
rect 9075 73883 9141 73884
rect 43302 71229 43362 178875
rect 44866 178500 44926 179520
rect 45602 178840 45662 179520
rect 46338 178840 46398 179520
rect 47074 178500 47134 179520
rect 47810 178840 47870 179520
rect 48546 178840 48606 179520
rect 49282 178840 49342 179520
rect 50018 178840 50078 179520
rect 50754 178840 50814 179520
rect 51490 178840 51550 179520
rect 52226 178840 52286 179520
rect 52962 178500 53022 179520
rect 53698 178500 53758 179520
rect 54434 178840 54494 179520
rect 55170 178500 55230 179520
rect 55906 178840 55966 179520
rect 56642 178500 56702 179520
rect 57378 178840 57438 179520
rect 58114 178840 58174 179520
rect 58850 178500 58910 179520
rect 59586 178500 59646 179520
rect 60322 178840 60382 179520
rect 61058 178500 61118 179520
rect 61794 178840 61854 179520
rect 62530 178840 62590 179520
rect 63266 178840 63326 179520
rect 64002 178840 64062 179520
rect 64738 178840 64798 179520
rect 65474 178840 65534 179520
rect 66210 178840 66270 179520
rect 66946 178840 67006 179520
rect 67682 178840 67742 179520
rect 68418 178876 68478 179520
rect 69154 178876 69214 179520
rect 69890 178876 69950 179520
rect 70626 178876 70686 179520
rect 71362 178876 71422 179520
rect 72098 178876 72158 179520
rect 72834 178876 72894 179520
rect 73570 178500 73630 179520
rect 74306 178500 74366 179520
rect 75042 178840 75102 179520
rect 75778 178876 75838 179520
rect 78998 178500 79058 179520
rect 79734 178840 79794 179520
rect 80470 178840 80530 179520
rect 81206 178500 81266 179520
rect 81942 178840 82002 179520
rect 82678 178840 82738 179520
rect 83414 178840 83474 179520
rect 84150 178840 84210 179520
rect 84886 178840 84946 179520
rect 85622 178840 85682 179520
rect 86358 178840 86418 179520
rect 87094 178500 87154 179520
rect 87830 178500 87890 179520
rect 88566 178840 88626 179520
rect 89302 178500 89362 179520
rect 90038 178840 90098 179520
rect 90774 178500 90834 179520
rect 91510 178840 91570 179520
rect 92246 178840 92306 179520
rect 92982 178500 93042 179520
rect 93718 178500 93778 179520
rect 94454 178840 94514 179520
rect 95190 178500 95250 179520
rect 95926 178840 95986 179520
rect 96662 178840 96722 179520
rect 97398 178840 97458 179520
rect 98134 178840 98194 179520
rect 98870 178840 98930 179520
rect 99606 178840 99666 179520
rect 100342 178840 100402 179520
rect 101078 178840 101138 179520
rect 101814 178840 101874 179520
rect 102550 178876 102610 179520
rect 103286 178876 103346 179520
rect 104022 178876 104082 179520
rect 104758 178876 104818 179520
rect 105494 178876 105554 179520
rect 106230 178876 106290 179520
rect 106966 178876 107026 179520
rect 107702 178500 107762 179520
rect 108438 178500 108498 179520
rect 109174 178840 109234 179520
rect 109910 178876 109970 179520
rect 111011 178804 111077 178805
rect 111011 178740 111012 178804
rect 111076 178740 111077 178804
rect 111011 178739 111077 178740
rect 48197 177879 48517 177936
rect 48197 177643 48239 177879
rect 48475 177643 48517 177879
rect 48197 177586 48517 177643
rect 56039 177879 56359 177936
rect 56039 177643 56081 177879
rect 56317 177643 56359 177879
rect 56039 177586 56359 177643
rect 63881 177879 64201 177936
rect 63881 177643 63923 177879
rect 64159 177643 64201 177879
rect 63881 177586 64201 177643
rect 71723 177879 72043 177936
rect 71723 177643 71765 177879
rect 72001 177643 72043 177879
rect 71723 177586 72043 177643
rect 82329 177879 82649 177936
rect 82329 177643 82371 177879
rect 82607 177643 82649 177879
rect 82329 177586 82649 177643
rect 90171 177879 90491 177936
rect 90171 177643 90213 177879
rect 90449 177643 90491 177879
rect 90171 177586 90491 177643
rect 98013 177879 98333 177936
rect 98013 177643 98055 177879
rect 98291 177643 98333 177879
rect 98013 177586 98333 177643
rect 105855 177879 106175 177936
rect 105855 177643 105897 177879
rect 106133 177643 106175 177879
rect 105855 177586 106175 177643
rect 52118 174454 52438 174486
rect 52118 174218 52160 174454
rect 52396 174218 52438 174454
rect 52118 174134 52438 174218
rect 52118 173898 52160 174134
rect 52396 173898 52438 174134
rect 52118 173866 52438 173898
rect 59960 174454 60280 174486
rect 59960 174218 60002 174454
rect 60238 174218 60280 174454
rect 59960 174134 60280 174218
rect 59960 173898 60002 174134
rect 60238 173898 60280 174134
rect 59960 173866 60280 173898
rect 67802 174454 68122 174486
rect 67802 174218 67844 174454
rect 68080 174218 68122 174454
rect 67802 174134 68122 174218
rect 67802 173898 67844 174134
rect 68080 173898 68122 174134
rect 67802 173866 68122 173898
rect 75644 174454 75964 174486
rect 75644 174218 75686 174454
rect 75922 174218 75964 174454
rect 75644 174134 75964 174218
rect 75644 173898 75686 174134
rect 75922 173898 75964 174134
rect 75644 173866 75964 173898
rect 86250 174454 86570 174486
rect 86250 174218 86292 174454
rect 86528 174218 86570 174454
rect 86250 174134 86570 174218
rect 86250 173898 86292 174134
rect 86528 173898 86570 174134
rect 86250 173866 86570 173898
rect 94092 174454 94412 174486
rect 94092 174218 94134 174454
rect 94370 174218 94412 174454
rect 94092 174134 94412 174218
rect 94092 173898 94134 174134
rect 94370 173898 94412 174134
rect 94092 173866 94412 173898
rect 101934 174454 102254 174486
rect 101934 174218 101976 174454
rect 102212 174218 102254 174454
rect 101934 174134 102254 174218
rect 101934 173898 101976 174134
rect 102212 173898 102254 174134
rect 101934 173866 102254 173898
rect 109776 174454 110096 174486
rect 109776 174218 109818 174454
rect 110054 174218 110096 174454
rect 109776 174134 110096 174218
rect 109776 173898 109818 174134
rect 110054 173898 110096 174134
rect 109776 173866 110096 173898
rect 48197 168174 48517 168206
rect 48197 167938 48239 168174
rect 48475 167938 48517 168174
rect 48197 167854 48517 167938
rect 48197 167618 48239 167854
rect 48475 167618 48517 167854
rect 48197 167586 48517 167618
rect 56039 168174 56359 168206
rect 56039 167938 56081 168174
rect 56317 167938 56359 168174
rect 56039 167854 56359 167938
rect 56039 167618 56081 167854
rect 56317 167618 56359 167854
rect 56039 167586 56359 167618
rect 63881 168174 64201 168206
rect 63881 167938 63923 168174
rect 64159 167938 64201 168174
rect 63881 167854 64201 167938
rect 63881 167618 63923 167854
rect 64159 167618 64201 167854
rect 63881 167586 64201 167618
rect 71723 168174 72043 168206
rect 71723 167938 71765 168174
rect 72001 167938 72043 168174
rect 71723 167854 72043 167938
rect 71723 167618 71765 167854
rect 72001 167618 72043 167854
rect 71723 167586 72043 167618
rect 82329 168174 82649 168206
rect 82329 167938 82371 168174
rect 82607 167938 82649 168174
rect 82329 167854 82649 167938
rect 82329 167618 82371 167854
rect 82607 167618 82649 167854
rect 82329 167586 82649 167618
rect 90171 168174 90491 168206
rect 90171 167938 90213 168174
rect 90449 167938 90491 168174
rect 90171 167854 90491 167938
rect 90171 167618 90213 167854
rect 90449 167618 90491 167854
rect 90171 167586 90491 167618
rect 98013 168174 98333 168206
rect 98013 167938 98055 168174
rect 98291 167938 98333 168174
rect 98013 167854 98333 167938
rect 98013 167618 98055 167854
rect 98291 167618 98333 167854
rect 98013 167586 98333 167618
rect 105855 168174 106175 168206
rect 105855 167938 105897 168174
rect 106133 167938 106175 168174
rect 105855 167854 106175 167938
rect 105855 167618 105897 167854
rect 106133 167618 106175 167854
rect 105855 167586 106175 167618
rect 52118 164454 52438 164486
rect 52118 164218 52160 164454
rect 52396 164218 52438 164454
rect 52118 164134 52438 164218
rect 52118 163898 52160 164134
rect 52396 163898 52438 164134
rect 52118 163866 52438 163898
rect 59960 164454 60280 164486
rect 59960 164218 60002 164454
rect 60238 164218 60280 164454
rect 59960 164134 60280 164218
rect 59960 163898 60002 164134
rect 60238 163898 60280 164134
rect 59960 163866 60280 163898
rect 67802 164454 68122 164486
rect 67802 164218 67844 164454
rect 68080 164218 68122 164454
rect 67802 164134 68122 164218
rect 67802 163898 67844 164134
rect 68080 163898 68122 164134
rect 67802 163866 68122 163898
rect 75644 164454 75964 164486
rect 75644 164218 75686 164454
rect 75922 164218 75964 164454
rect 75644 164134 75964 164218
rect 75644 163898 75686 164134
rect 75922 163898 75964 164134
rect 75644 163866 75964 163898
rect 86250 164454 86570 164486
rect 86250 164218 86292 164454
rect 86528 164218 86570 164454
rect 86250 164134 86570 164218
rect 86250 163898 86292 164134
rect 86528 163898 86570 164134
rect 86250 163866 86570 163898
rect 94092 164454 94412 164486
rect 94092 164218 94134 164454
rect 94370 164218 94412 164454
rect 94092 164134 94412 164218
rect 94092 163898 94134 164134
rect 94370 163898 94412 164134
rect 94092 163866 94412 163898
rect 101934 164454 102254 164486
rect 101934 164218 101976 164454
rect 102212 164218 102254 164454
rect 101934 164134 102254 164218
rect 101934 163898 101976 164134
rect 102212 163898 102254 164134
rect 101934 163866 102254 163898
rect 109776 164454 110096 164486
rect 109776 164218 109818 164454
rect 110054 164218 110096 164454
rect 109776 164134 110096 164218
rect 109776 163898 109818 164134
rect 110054 163898 110096 164134
rect 109776 163866 110096 163898
rect 43299 71228 43365 71229
rect 43299 71164 43300 71228
rect 43364 71164 43365 71228
rect 43299 71163 43365 71164
rect 8891 69596 8957 69597
rect 8891 69532 8892 69596
rect 8956 69532 8957 69596
rect 8891 69531 8957 69532
rect 111014 67013 111074 178739
rect 113130 178500 113190 179520
rect 113866 178840 113926 179520
rect 114602 178840 114662 179520
rect 115338 178500 115398 179520
rect 116074 178840 116134 179520
rect 116810 178840 116870 179520
rect 117546 178840 117606 179520
rect 118282 178840 118342 179520
rect 119018 178840 119078 179520
rect 119754 178840 119814 179520
rect 120490 178840 120550 179520
rect 121226 178500 121286 179520
rect 121962 178500 122022 179520
rect 122698 178840 122758 179520
rect 123434 178500 123494 179520
rect 124170 178840 124230 179520
rect 124906 178500 124966 179520
rect 125642 178840 125702 179520
rect 126378 178840 126438 179520
rect 127114 178500 127174 179520
rect 127850 178500 127910 179520
rect 128586 178840 128646 179520
rect 129322 178500 129382 179520
rect 130058 178840 130118 179520
rect 130794 178840 130854 179520
rect 131530 178840 131590 179520
rect 132266 178840 132326 179520
rect 133002 178840 133062 179520
rect 133738 178840 133798 179520
rect 134474 178840 134534 179520
rect 135210 178840 135270 179520
rect 135946 178840 136006 179520
rect 136682 178876 136742 179520
rect 137418 178876 137478 179520
rect 138154 178876 138214 179520
rect 138890 178876 138950 179520
rect 139626 178876 139686 179520
rect 140362 178876 140422 179520
rect 141098 178876 141158 179520
rect 141834 178500 141894 179520
rect 142570 178500 142630 179520
rect 143306 178840 143366 179520
rect 144042 178876 144102 179520
rect 147262 178500 147322 179520
rect 147998 178840 148058 179520
rect 148734 178840 148794 179520
rect 149470 178500 149530 179520
rect 150206 178840 150266 179520
rect 150942 178840 151002 179520
rect 151678 178840 151738 179520
rect 152414 178840 152474 179520
rect 153150 178840 153210 179520
rect 153886 178840 153946 179520
rect 154622 178840 154682 179520
rect 155358 178500 155418 179520
rect 156094 178500 156154 179520
rect 156830 178840 156890 179520
rect 157566 178500 157626 179520
rect 158302 178840 158362 179520
rect 159038 178500 159098 179520
rect 159774 178840 159834 179520
rect 160510 178840 160570 179520
rect 161246 178500 161306 179520
rect 161982 178500 162042 179520
rect 162718 178840 162778 179520
rect 163454 178500 163514 179520
rect 164190 178840 164250 179520
rect 164926 178840 164986 179520
rect 165662 178840 165722 179520
rect 166398 178840 166458 179860
rect 167134 178840 167194 179520
rect 167870 178840 167930 179520
rect 168606 178840 168666 179860
rect 169342 178840 169402 179520
rect 170078 178840 170138 179520
rect 170814 178876 170874 179520
rect 171550 178876 171610 179520
rect 172286 178876 172346 179520
rect 173022 178876 173082 179520
rect 173758 178876 173818 179520
rect 174494 178876 174554 179520
rect 175230 178876 175290 179520
rect 175966 178500 176026 179520
rect 176702 178500 176762 179520
rect 177438 178840 177498 179520
rect 178174 178876 178234 179520
rect 181394 178500 181454 179520
rect 182130 178840 182190 179520
rect 182866 178840 182926 179520
rect 183602 178500 183662 179520
rect 184338 178840 184398 179520
rect 185074 178840 185134 179520
rect 185810 178840 185870 179520
rect 186546 178840 186606 179520
rect 187282 178840 187342 179520
rect 188018 178840 188078 179520
rect 188754 178840 188814 179520
rect 189490 178500 189550 179520
rect 190226 178500 190286 179520
rect 190962 178840 191022 179520
rect 191698 178500 191758 179520
rect 192434 178840 192494 179520
rect 193170 178500 193230 179520
rect 193906 178840 193966 179520
rect 194642 178840 194702 179520
rect 195378 178500 195438 179520
rect 196114 178500 196174 179520
rect 196850 178840 196910 179520
rect 197586 178500 197646 179520
rect 198322 178840 198382 179520
rect 199058 178840 199118 179520
rect 199794 178840 199854 179520
rect 200530 178840 200590 179520
rect 201266 178840 201326 179520
rect 202002 178840 202062 179520
rect 202738 178840 202798 179520
rect 203474 178840 203534 179520
rect 204210 178840 204270 179520
rect 204946 178876 205006 179520
rect 205682 178876 205742 179520
rect 206418 178876 206478 179520
rect 207154 178876 207214 179520
rect 207890 178876 207950 179520
rect 208626 178876 208686 179520
rect 209362 178876 209422 179520
rect 210098 178500 210158 179520
rect 210834 178500 210894 179520
rect 211570 178840 211630 179520
rect 212306 178876 212366 179520
rect 215526 178500 215586 179520
rect 216262 178840 216322 179520
rect 216998 178840 217058 179520
rect 217734 178500 217794 179520
rect 218470 178840 218530 179520
rect 219206 178840 219266 179520
rect 219942 178840 220002 179520
rect 220678 178840 220738 179520
rect 221414 178840 221474 179520
rect 222150 178840 222210 179520
rect 222886 178840 222946 179520
rect 223622 178500 223682 179520
rect 224358 178500 224418 179520
rect 225094 178840 225154 179520
rect 225830 178500 225890 179520
rect 226566 178840 226626 179520
rect 227302 178500 227362 179520
rect 228038 178840 228098 179520
rect 228774 178840 228834 179520
rect 229510 178500 229570 179520
rect 230246 178500 230306 179520
rect 230982 178840 231042 179520
rect 231718 178500 231778 179520
rect 232454 178840 232514 179860
rect 233190 178840 233250 179520
rect 233926 178840 233986 179860
rect 234662 178840 234722 179520
rect 235398 178840 235458 179860
rect 236134 178840 236194 179520
rect 236870 178840 236930 179520
rect 237606 178840 237666 179520
rect 238342 178840 238402 179520
rect 239078 178876 239138 179520
rect 239814 178876 239874 179520
rect 240550 178876 240610 179520
rect 241286 178876 241346 179520
rect 242022 178876 242082 179520
rect 242758 178876 242818 179520
rect 243494 178876 243554 179520
rect 244230 178500 244290 179520
rect 244966 178500 245026 179860
rect 245702 178840 245762 179520
rect 246438 178876 246498 179520
rect 248091 178668 248157 178669
rect 248091 178604 248092 178668
rect 248156 178604 248157 178668
rect 248091 178603 248157 178604
rect 116461 177879 116781 177936
rect 116461 177643 116503 177879
rect 116739 177643 116781 177879
rect 116461 177586 116781 177643
rect 124303 177879 124623 177936
rect 124303 177643 124345 177879
rect 124581 177643 124623 177879
rect 124303 177586 124623 177643
rect 132145 177879 132465 177936
rect 132145 177643 132187 177879
rect 132423 177643 132465 177879
rect 132145 177586 132465 177643
rect 139987 177879 140307 177936
rect 139987 177643 140029 177879
rect 140265 177643 140307 177879
rect 139987 177586 140307 177643
rect 150593 177879 150913 177936
rect 150593 177643 150635 177879
rect 150871 177643 150913 177879
rect 150593 177586 150913 177643
rect 158435 177879 158755 177936
rect 158435 177643 158477 177879
rect 158713 177643 158755 177879
rect 158435 177586 158755 177643
rect 166277 177879 166597 177936
rect 166277 177643 166319 177879
rect 166555 177643 166597 177879
rect 166277 177586 166597 177643
rect 174119 177879 174439 177936
rect 174119 177643 174161 177879
rect 174397 177643 174439 177879
rect 174119 177586 174439 177643
rect 184725 177879 185045 177936
rect 184725 177643 184767 177879
rect 185003 177643 185045 177879
rect 184725 177586 185045 177643
rect 192567 177879 192887 177936
rect 192567 177643 192609 177879
rect 192845 177643 192887 177879
rect 192567 177586 192887 177643
rect 200409 177879 200729 177936
rect 200409 177643 200451 177879
rect 200687 177643 200729 177879
rect 200409 177586 200729 177643
rect 208251 177879 208571 177936
rect 208251 177643 208293 177879
rect 208529 177643 208571 177879
rect 208251 177586 208571 177643
rect 218857 177879 219177 177936
rect 218857 177643 218899 177879
rect 219135 177643 219177 177879
rect 218857 177586 219177 177643
rect 226699 177879 227019 177936
rect 226699 177643 226741 177879
rect 226977 177643 227019 177879
rect 226699 177586 227019 177643
rect 234541 177879 234861 177936
rect 234541 177643 234583 177879
rect 234819 177643 234861 177879
rect 234541 177586 234861 177643
rect 242383 177879 242703 177936
rect 242383 177643 242425 177879
rect 242661 177643 242703 177879
rect 242383 177586 242703 177643
rect 120382 174454 120702 174486
rect 120382 174218 120424 174454
rect 120660 174218 120702 174454
rect 120382 174134 120702 174218
rect 120382 173898 120424 174134
rect 120660 173898 120702 174134
rect 120382 173866 120702 173898
rect 128224 174454 128544 174486
rect 128224 174218 128266 174454
rect 128502 174218 128544 174454
rect 128224 174134 128544 174218
rect 128224 173898 128266 174134
rect 128502 173898 128544 174134
rect 128224 173866 128544 173898
rect 136066 174454 136386 174486
rect 136066 174218 136108 174454
rect 136344 174218 136386 174454
rect 136066 174134 136386 174218
rect 136066 173898 136108 174134
rect 136344 173898 136386 174134
rect 136066 173866 136386 173898
rect 143908 174454 144228 174486
rect 143908 174218 143950 174454
rect 144186 174218 144228 174454
rect 143908 174134 144228 174218
rect 143908 173898 143950 174134
rect 144186 173898 144228 174134
rect 143908 173866 144228 173898
rect 154514 174454 154834 174486
rect 154514 174218 154556 174454
rect 154792 174218 154834 174454
rect 154514 174134 154834 174218
rect 154514 173898 154556 174134
rect 154792 173898 154834 174134
rect 154514 173866 154834 173898
rect 162356 174454 162676 174486
rect 162356 174218 162398 174454
rect 162634 174218 162676 174454
rect 162356 174134 162676 174218
rect 162356 173898 162398 174134
rect 162634 173898 162676 174134
rect 162356 173866 162676 173898
rect 170198 174454 170518 174486
rect 170198 174218 170240 174454
rect 170476 174218 170518 174454
rect 170198 174134 170518 174218
rect 170198 173898 170240 174134
rect 170476 173898 170518 174134
rect 170198 173866 170518 173898
rect 178040 174454 178360 174486
rect 178040 174218 178082 174454
rect 178318 174218 178360 174454
rect 178040 174134 178360 174218
rect 178040 173898 178082 174134
rect 178318 173898 178360 174134
rect 178040 173866 178360 173898
rect 188646 174454 188966 174486
rect 188646 174218 188688 174454
rect 188924 174218 188966 174454
rect 188646 174134 188966 174218
rect 188646 173898 188688 174134
rect 188924 173898 188966 174134
rect 188646 173866 188966 173898
rect 196488 174454 196808 174486
rect 196488 174218 196530 174454
rect 196766 174218 196808 174454
rect 196488 174134 196808 174218
rect 196488 173898 196530 174134
rect 196766 173898 196808 174134
rect 196488 173866 196808 173898
rect 204330 174454 204650 174486
rect 204330 174218 204372 174454
rect 204608 174218 204650 174454
rect 204330 174134 204650 174218
rect 204330 173898 204372 174134
rect 204608 173898 204650 174134
rect 204330 173866 204650 173898
rect 212172 174454 212492 174486
rect 212172 174218 212214 174454
rect 212450 174218 212492 174454
rect 212172 174134 212492 174218
rect 212172 173898 212214 174134
rect 212450 173898 212492 174134
rect 212172 173866 212492 173898
rect 222778 174454 223098 174486
rect 222778 174218 222820 174454
rect 223056 174218 223098 174454
rect 222778 174134 223098 174218
rect 222778 173898 222820 174134
rect 223056 173898 223098 174134
rect 222778 173866 223098 173898
rect 230620 174454 230940 174486
rect 230620 174218 230662 174454
rect 230898 174218 230940 174454
rect 230620 174134 230940 174218
rect 230620 173898 230662 174134
rect 230898 173898 230940 174134
rect 230620 173866 230940 173898
rect 238462 174454 238782 174486
rect 238462 174218 238504 174454
rect 238740 174218 238782 174454
rect 238462 174134 238782 174218
rect 238462 173898 238504 174134
rect 238740 173898 238782 174134
rect 238462 173866 238782 173898
rect 246304 174454 246624 174486
rect 246304 174218 246346 174454
rect 246582 174218 246624 174454
rect 246304 174134 246624 174218
rect 246304 173898 246346 174134
rect 246582 173898 246624 174134
rect 246304 173866 246624 173898
rect 116461 168174 116781 168206
rect 116461 167938 116503 168174
rect 116739 167938 116781 168174
rect 116461 167854 116781 167938
rect 116461 167618 116503 167854
rect 116739 167618 116781 167854
rect 116461 167586 116781 167618
rect 124303 168174 124623 168206
rect 124303 167938 124345 168174
rect 124581 167938 124623 168174
rect 124303 167854 124623 167938
rect 124303 167618 124345 167854
rect 124581 167618 124623 167854
rect 124303 167586 124623 167618
rect 132145 168174 132465 168206
rect 132145 167938 132187 168174
rect 132423 167938 132465 168174
rect 132145 167854 132465 167938
rect 132145 167618 132187 167854
rect 132423 167618 132465 167854
rect 132145 167586 132465 167618
rect 139987 168174 140307 168206
rect 139987 167938 140029 168174
rect 140265 167938 140307 168174
rect 139987 167854 140307 167938
rect 139987 167618 140029 167854
rect 140265 167618 140307 167854
rect 139987 167586 140307 167618
rect 150593 168174 150913 168206
rect 150593 167938 150635 168174
rect 150871 167938 150913 168174
rect 150593 167854 150913 167938
rect 150593 167618 150635 167854
rect 150871 167618 150913 167854
rect 150593 167586 150913 167618
rect 158435 168174 158755 168206
rect 158435 167938 158477 168174
rect 158713 167938 158755 168174
rect 158435 167854 158755 167938
rect 158435 167618 158477 167854
rect 158713 167618 158755 167854
rect 158435 167586 158755 167618
rect 166277 168174 166597 168206
rect 166277 167938 166319 168174
rect 166555 167938 166597 168174
rect 166277 167854 166597 167938
rect 166277 167618 166319 167854
rect 166555 167618 166597 167854
rect 166277 167586 166597 167618
rect 174119 168174 174439 168206
rect 174119 167938 174161 168174
rect 174397 167938 174439 168174
rect 174119 167854 174439 167938
rect 174119 167618 174161 167854
rect 174397 167618 174439 167854
rect 174119 167586 174439 167618
rect 184725 168174 185045 168206
rect 184725 167938 184767 168174
rect 185003 167938 185045 168174
rect 184725 167854 185045 167938
rect 184725 167618 184767 167854
rect 185003 167618 185045 167854
rect 184725 167586 185045 167618
rect 192567 168174 192887 168206
rect 192567 167938 192609 168174
rect 192845 167938 192887 168174
rect 192567 167854 192887 167938
rect 192567 167618 192609 167854
rect 192845 167618 192887 167854
rect 192567 167586 192887 167618
rect 200409 168174 200729 168206
rect 200409 167938 200451 168174
rect 200687 167938 200729 168174
rect 200409 167854 200729 167938
rect 200409 167618 200451 167854
rect 200687 167618 200729 167854
rect 200409 167586 200729 167618
rect 208251 168174 208571 168206
rect 208251 167938 208293 168174
rect 208529 167938 208571 168174
rect 208251 167854 208571 167938
rect 208251 167618 208293 167854
rect 208529 167618 208571 167854
rect 208251 167586 208571 167618
rect 218857 168174 219177 168206
rect 218857 167938 218899 168174
rect 219135 167938 219177 168174
rect 218857 167854 219177 167938
rect 218857 167618 218899 167854
rect 219135 167618 219177 167854
rect 218857 167586 219177 167618
rect 226699 168174 227019 168206
rect 226699 167938 226741 168174
rect 226977 167938 227019 168174
rect 226699 167854 227019 167938
rect 226699 167618 226741 167854
rect 226977 167618 227019 167854
rect 226699 167586 227019 167618
rect 234541 168174 234861 168206
rect 234541 167938 234583 168174
rect 234819 167938 234861 168174
rect 234541 167854 234861 167938
rect 234541 167618 234583 167854
rect 234819 167618 234861 167854
rect 234541 167586 234861 167618
rect 242383 168174 242703 168206
rect 242383 167938 242425 168174
rect 242661 167938 242703 168174
rect 242383 167854 242703 167938
rect 242383 167618 242425 167854
rect 242661 167618 242703 167854
rect 242383 167586 242703 167618
rect 120382 164454 120702 164486
rect 120382 164218 120424 164454
rect 120660 164218 120702 164454
rect 120382 164134 120702 164218
rect 120382 163898 120424 164134
rect 120660 163898 120702 164134
rect 120382 163866 120702 163898
rect 128224 164454 128544 164486
rect 128224 164218 128266 164454
rect 128502 164218 128544 164454
rect 128224 164134 128544 164218
rect 128224 163898 128266 164134
rect 128502 163898 128544 164134
rect 128224 163866 128544 163898
rect 136066 164454 136386 164486
rect 136066 164218 136108 164454
rect 136344 164218 136386 164454
rect 136066 164134 136386 164218
rect 136066 163898 136108 164134
rect 136344 163898 136386 164134
rect 136066 163866 136386 163898
rect 143908 164454 144228 164486
rect 143908 164218 143950 164454
rect 144186 164218 144228 164454
rect 143908 164134 144228 164218
rect 143908 163898 143950 164134
rect 144186 163898 144228 164134
rect 143908 163866 144228 163898
rect 154514 164454 154834 164486
rect 154514 164218 154556 164454
rect 154792 164218 154834 164454
rect 154514 164134 154834 164218
rect 154514 163898 154556 164134
rect 154792 163898 154834 164134
rect 154514 163866 154834 163898
rect 162356 164454 162676 164486
rect 162356 164218 162398 164454
rect 162634 164218 162676 164454
rect 162356 164134 162676 164218
rect 162356 163898 162398 164134
rect 162634 163898 162676 164134
rect 162356 163866 162676 163898
rect 170198 164454 170518 164486
rect 170198 164218 170240 164454
rect 170476 164218 170518 164454
rect 170198 164134 170518 164218
rect 170198 163898 170240 164134
rect 170476 163898 170518 164134
rect 170198 163866 170518 163898
rect 178040 164454 178360 164486
rect 178040 164218 178082 164454
rect 178318 164218 178360 164454
rect 178040 164134 178360 164218
rect 178040 163898 178082 164134
rect 178318 163898 178360 164134
rect 178040 163866 178360 163898
rect 188646 164454 188966 164486
rect 188646 164218 188688 164454
rect 188924 164218 188966 164454
rect 188646 164134 188966 164218
rect 188646 163898 188688 164134
rect 188924 163898 188966 164134
rect 188646 163866 188966 163898
rect 196488 164454 196808 164486
rect 196488 164218 196530 164454
rect 196766 164218 196808 164454
rect 196488 164134 196808 164218
rect 196488 163898 196530 164134
rect 196766 163898 196808 164134
rect 196488 163866 196808 163898
rect 204330 164454 204650 164486
rect 204330 164218 204372 164454
rect 204608 164218 204650 164454
rect 204330 164134 204650 164218
rect 204330 163898 204372 164134
rect 204608 163898 204650 164134
rect 204330 163866 204650 163898
rect 212172 164454 212492 164486
rect 212172 164218 212214 164454
rect 212450 164218 212492 164454
rect 212172 164134 212492 164218
rect 212172 163898 212214 164134
rect 212450 163898 212492 164134
rect 212172 163866 212492 163898
rect 222778 164454 223098 164486
rect 222778 164218 222820 164454
rect 223056 164218 223098 164454
rect 222778 164134 223098 164218
rect 222778 163898 222820 164134
rect 223056 163898 223098 164134
rect 222778 163866 223098 163898
rect 230620 164454 230940 164486
rect 230620 164218 230662 164454
rect 230898 164218 230940 164454
rect 230620 164134 230940 164218
rect 230620 163898 230662 164134
rect 230898 163898 230940 164134
rect 230620 163866 230940 163898
rect 238462 164454 238782 164486
rect 238462 164218 238504 164454
rect 238740 164218 238782 164454
rect 238462 164134 238782 164218
rect 238462 163898 238504 164134
rect 238740 163898 238782 164134
rect 238462 163866 238782 163898
rect 246304 164454 246624 164486
rect 246304 164218 246346 164454
rect 246582 164218 246624 164454
rect 246304 164134 246624 164218
rect 246304 163898 246346 164134
rect 246582 163898 246624 164134
rect 246304 163866 246624 163898
rect 248094 156773 248154 178603
rect 249658 178500 249718 179520
rect 250394 178840 250454 179520
rect 251130 178840 251190 179520
rect 251866 178500 251926 179520
rect 252602 178840 252662 179520
rect 253338 178840 253398 179520
rect 254074 178840 254134 179520
rect 254810 178840 254870 179520
rect 255546 178840 255606 179520
rect 256282 178840 256342 179520
rect 257018 178840 257078 179520
rect 257754 178500 257814 179520
rect 258490 178500 258550 179520
rect 259226 178840 259286 179520
rect 259962 178500 260022 179520
rect 260698 178840 260758 179520
rect 261434 178500 261494 179520
rect 262170 178840 262230 179520
rect 262906 178840 262966 179520
rect 263642 178500 263702 179520
rect 264378 178500 264438 179520
rect 265114 178840 265174 179520
rect 265850 178500 265910 179520
rect 266586 178840 266646 179520
rect 267322 178840 267382 179520
rect 268058 178840 268118 179520
rect 268794 178840 268854 179520
rect 269530 178840 269590 179520
rect 270266 178840 270326 179520
rect 271002 178840 271062 179520
rect 271738 178840 271798 179520
rect 272474 178840 272534 179520
rect 273210 178876 273270 179520
rect 273946 178876 274006 179520
rect 274682 178876 274742 179520
rect 275418 178876 275478 179520
rect 276154 178876 276214 179520
rect 276890 178876 276950 179520
rect 277626 178876 277686 179520
rect 278362 178500 278422 179520
rect 279098 178500 279158 179520
rect 279834 178840 279894 179520
rect 280570 178876 280630 179520
rect 281582 178669 281642 181051
rect 281947 180844 282013 180845
rect 281947 180780 281948 180844
rect 282012 180780 282013 180844
rect 281947 180779 282013 180780
rect 281579 178668 281645 178669
rect 281579 178604 281580 178668
rect 281644 178604 281645 178668
rect 281579 178603 281645 178604
rect 281211 177988 281277 177989
rect 252989 177879 253309 177936
rect 252989 177643 253031 177879
rect 253267 177643 253309 177879
rect 252989 177586 253309 177643
rect 260831 177879 261151 177936
rect 260831 177643 260873 177879
rect 261109 177643 261151 177879
rect 260831 177586 261151 177643
rect 268673 177879 268993 177936
rect 268673 177643 268715 177879
rect 268951 177643 268993 177879
rect 268673 177586 268993 177643
rect 276515 177879 276835 177936
rect 281211 177924 281212 177988
rect 281276 177924 281277 177988
rect 281211 177923 281277 177924
rect 276515 177643 276557 177879
rect 276793 177643 276835 177879
rect 276515 177586 276835 177643
rect 256910 174454 257230 174486
rect 256910 174218 256952 174454
rect 257188 174218 257230 174454
rect 256910 174134 257230 174218
rect 256910 173898 256952 174134
rect 257188 173898 257230 174134
rect 256910 173866 257230 173898
rect 264752 174454 265072 174486
rect 264752 174218 264794 174454
rect 265030 174218 265072 174454
rect 264752 174134 265072 174218
rect 264752 173898 264794 174134
rect 265030 173898 265072 174134
rect 264752 173866 265072 173898
rect 272594 174454 272914 174486
rect 272594 174218 272636 174454
rect 272872 174218 272914 174454
rect 272594 174134 272914 174218
rect 272594 173898 272636 174134
rect 272872 173898 272914 174134
rect 272594 173866 272914 173898
rect 280436 174454 280756 174486
rect 280436 174218 280478 174454
rect 280714 174218 280756 174454
rect 280436 174134 280756 174218
rect 280436 173898 280478 174134
rect 280714 173898 280756 174134
rect 280436 173866 280756 173898
rect 252989 168174 253309 168206
rect 252989 167938 253031 168174
rect 253267 167938 253309 168174
rect 252989 167854 253309 167938
rect 252989 167618 253031 167854
rect 253267 167618 253309 167854
rect 252989 167586 253309 167618
rect 260831 168174 261151 168206
rect 260831 167938 260873 168174
rect 261109 167938 261151 168174
rect 260831 167854 261151 167938
rect 260831 167618 260873 167854
rect 261109 167618 261151 167854
rect 260831 167586 261151 167618
rect 268673 168174 268993 168206
rect 268673 167938 268715 168174
rect 268951 167938 268993 168174
rect 268673 167854 268993 167938
rect 268673 167618 268715 167854
rect 268951 167618 268993 167854
rect 268673 167586 268993 167618
rect 276515 168174 276835 168206
rect 276515 167938 276557 168174
rect 276793 167938 276835 168174
rect 276515 167854 276835 167938
rect 276515 167618 276557 167854
rect 276793 167618 276835 167854
rect 276515 167586 276835 167618
rect 256910 164454 257230 164486
rect 256910 164218 256952 164454
rect 257188 164218 257230 164454
rect 256910 164134 257230 164218
rect 256910 163898 256952 164134
rect 257188 163898 257230 164134
rect 256910 163866 257230 163898
rect 264752 164454 265072 164486
rect 264752 164218 264794 164454
rect 265030 164218 265072 164454
rect 264752 164134 265072 164218
rect 264752 163898 264794 164134
rect 265030 163898 265072 164134
rect 264752 163866 265072 163898
rect 272594 164454 272914 164486
rect 272594 164218 272636 164454
rect 272872 164218 272914 164454
rect 272594 164134 272914 164218
rect 272594 163898 272636 164134
rect 272872 163898 272914 164134
rect 272594 163866 272914 163898
rect 280436 164454 280756 164486
rect 280436 164218 280478 164454
rect 280714 164218 280756 164454
rect 280436 164134 280756 164218
rect 280436 163898 280478 164134
rect 280714 163898 280756 164134
rect 280436 163866 280756 163898
rect 277163 157996 277229 157997
rect 277163 157932 277164 157996
rect 277228 157932 277229 157996
rect 277163 157931 277229 157932
rect 248091 156772 248157 156773
rect 248091 156708 248092 156772
rect 248156 156708 248157 156772
rect 248091 156707 248157 156708
rect 264099 156772 264165 156773
rect 264099 156708 264100 156772
rect 264164 156708 264165 156772
rect 264099 156707 264165 156708
rect 264102 71365 264162 156707
rect 272379 156636 272445 156637
rect 272379 156572 272380 156636
rect 272444 156572 272445 156636
rect 272379 156571 272445 156572
rect 274403 156636 274469 156637
rect 274403 156572 274404 156636
rect 274468 156572 274469 156636
rect 274403 156571 274469 156572
rect 269619 155276 269685 155277
rect 269619 155212 269620 155276
rect 269684 155212 269685 155276
rect 269619 155211 269685 155212
rect 264099 71364 264165 71365
rect 264099 71300 264100 71364
rect 264164 71300 264165 71364
rect 264099 71299 264165 71300
rect 111011 67012 111077 67013
rect 111011 66948 111012 67012
rect 111076 66948 111077 67012
rect 111011 66947 111077 66948
rect 269622 21997 269682 155211
rect 271091 149700 271157 149701
rect 271091 149636 271092 149700
rect 271156 149636 271157 149700
rect 271091 149635 271157 149636
rect 269619 21996 269685 21997
rect 269619 21932 269620 21996
rect 269684 21932 269685 21996
rect 269619 21931 269685 21932
rect 8155 21860 8221 21861
rect 8155 21796 8156 21860
rect 8220 21796 8221 21860
rect 8155 21795 8221 21796
rect 7603 19276 7669 19277
rect 7603 19212 7604 19276
rect 7668 19212 7669 19276
rect 7603 19211 7669 19212
rect 271094 19005 271154 149635
rect 272382 19141 272442 156571
rect 274219 73948 274285 73949
rect 274219 73884 274220 73948
rect 274284 73884 274285 73948
rect 274219 73883 274285 73884
rect 272563 71364 272629 71365
rect 272563 71300 272564 71364
rect 272628 71300 272629 71364
rect 272563 71299 272629 71300
rect 272566 68645 272626 71299
rect 272563 68644 272629 68645
rect 272563 68580 272564 68644
rect 272628 68580 272629 68644
rect 272563 68579 272629 68580
rect 274222 65620 274282 73883
rect 274406 69733 274466 156571
rect 274587 152420 274653 152421
rect 274587 152356 274588 152420
rect 274652 152356 274653 152420
rect 274587 152355 274653 152356
rect 274403 69732 274469 69733
rect 274403 69668 274404 69732
rect 274468 69668 274469 69732
rect 274403 69667 274469 69668
rect 274590 65620 274650 152355
rect 276795 87548 276861 87549
rect 276795 87484 276796 87548
rect 276860 87484 276861 87548
rect 276795 87483 276861 87484
rect 276059 71228 276125 71229
rect 276059 71164 276060 71228
rect 276124 71164 276125 71228
rect 276059 71163 276125 71164
rect 274955 71092 275021 71093
rect 274955 71028 274956 71092
rect 275020 71028 275021 71092
rect 274955 71027 275021 71028
rect 274958 65620 275018 71027
rect 275323 68372 275389 68373
rect 275323 68308 275324 68372
rect 275388 68308 275389 68372
rect 275323 68307 275389 68308
rect 275326 65620 275386 68307
rect 275691 66876 275757 66877
rect 275691 66812 275692 66876
rect 275756 66812 275757 66876
rect 275691 66811 275757 66812
rect 275694 65620 275754 66811
rect 276062 65620 276122 71163
rect 276427 68236 276493 68237
rect 276427 68172 276428 68236
rect 276492 68172 276493 68236
rect 276427 68171 276493 68172
rect 276430 65620 276490 68171
rect 276798 65620 276858 87483
rect 277166 71093 277226 157931
rect 279923 157452 279989 157453
rect 279923 157388 279924 157452
rect 279988 157388 279989 157452
rect 279923 157387 279989 157388
rect 279003 153780 279069 153781
rect 279003 153716 279004 153780
rect 279068 153716 279069 153780
rect 279003 153715 279069 153716
rect 277531 151060 277597 151061
rect 277531 150996 277532 151060
rect 277596 150996 277597 151060
rect 277531 150995 277597 150996
rect 277163 71092 277229 71093
rect 277163 71028 277164 71092
rect 277228 71028 277229 71092
rect 277163 71027 277229 71028
rect 277163 67012 277229 67013
rect 277163 66948 277164 67012
rect 277228 66948 277229 67012
rect 277163 66947 277229 66948
rect 277166 65620 277226 66947
rect 277534 65620 277594 150995
rect 278267 73812 278333 73813
rect 278267 73748 278268 73812
rect 278332 73748 278333 73812
rect 278267 73747 278333 73748
rect 277899 68236 277965 68237
rect 277899 68172 277900 68236
rect 277964 68172 277965 68236
rect 277899 68171 277965 68172
rect 277902 65620 277962 68171
rect 278270 65620 278330 73747
rect 278635 69596 278701 69597
rect 278635 69532 278636 69596
rect 278700 69532 278701 69596
rect 278635 69531 278701 69532
rect 278638 65620 278698 69531
rect 279006 65620 279066 153715
rect 279926 68917 279986 157387
rect 280291 76532 280357 76533
rect 280291 76468 280292 76532
rect 280356 76468 280357 76532
rect 280291 76467 280357 76468
rect 280294 74550 280354 76467
rect 280110 74490 280354 74550
rect 279923 68916 279989 68917
rect 279923 68852 279924 68916
rect 279988 68852 279989 68916
rect 279923 68851 279989 68852
rect 279739 68508 279805 68509
rect 279739 68444 279740 68508
rect 279804 68444 279805 68508
rect 279739 68443 279805 68444
rect 279371 67556 279437 67557
rect 279371 67492 279372 67556
rect 279436 67492 279437 67556
rect 279371 67491 279437 67492
rect 279374 65620 279434 67491
rect 279742 65620 279802 68443
rect 280110 65620 280170 74490
rect 281214 65724 281274 177923
rect 281950 161490 282010 180779
rect 282499 180708 282565 180709
rect 282499 180644 282500 180708
rect 282564 180644 282565 180708
rect 282499 180643 282565 180644
rect 282131 175948 282197 175949
rect 282131 175884 282132 175948
rect 282196 175884 282197 175948
rect 282131 175883 282197 175884
rect 281766 161430 282010 161490
rect 281766 157997 281826 161430
rect 281763 157996 281829 157997
rect 281763 157932 281764 157996
rect 281828 157932 281829 157996
rect 281763 157931 281829 157932
rect 282134 157453 282194 175883
rect 282131 157452 282197 157453
rect 282131 157388 282132 157452
rect 282196 157388 282197 157452
rect 282131 157387 282197 157388
rect 282502 74550 282562 180643
rect 282867 180572 282933 180573
rect 282867 180508 282868 180572
rect 282932 180508 282933 180572
rect 282867 180507 282933 180508
rect 282870 177989 282930 180507
rect 282867 177988 282933 177989
rect 282867 177924 282868 177988
rect 282932 177924 282933 177988
rect 282867 177923 282933 177924
rect 283054 175949 283114 181595
rect 284339 181524 284405 181525
rect 284339 181460 284340 181524
rect 284404 181460 284405 181524
rect 284339 181459 284405 181460
rect 283419 181388 283485 181389
rect 283419 181324 283420 181388
rect 283484 181324 283485 181388
rect 283419 181323 283485 181324
rect 283422 180437 283482 181323
rect 283419 180436 283485 180437
rect 283419 180372 283420 180436
rect 283484 180372 283485 180436
rect 283419 180371 283485 180372
rect 283051 175948 283117 175949
rect 283051 175884 283052 175948
rect 283116 175884 283117 175948
rect 283051 175883 283117 175884
rect 283422 156637 283482 180371
rect 284342 177170 284402 181459
rect 283790 177110 284402 177170
rect 283419 156636 283485 156637
rect 283419 156572 283420 156636
rect 283484 156572 283485 156636
rect 283419 156571 283485 156572
rect 281766 74490 282562 74550
rect 281766 65650 281826 74490
rect 281947 71092 282013 71093
rect 281947 71028 281948 71092
rect 282012 71028 282013 71092
rect 281947 71027 282013 71028
rect 281612 65590 281826 65650
rect 281950 65620 282010 71027
rect 283419 69732 283485 69733
rect 283419 69668 283420 69732
rect 283484 69668 283485 69732
rect 283419 69667 283485 69668
rect 282683 68644 282749 68645
rect 282683 68580 282684 68644
rect 282748 68580 282749 68644
rect 282683 68579 282749 68580
rect 282315 67692 282381 67693
rect 282315 67628 282316 67692
rect 282380 67628 282381 67692
rect 282315 67627 282381 67628
rect 282318 65620 282378 67627
rect 282686 65620 282746 68579
rect 283051 67556 283117 67557
rect 283051 67492 283052 67556
rect 283116 67492 283117 67556
rect 283051 67491 283117 67492
rect 283054 65620 283114 67491
rect 283422 65620 283482 69667
rect 283790 65620 283850 177110
rect 284155 68916 284221 68917
rect 284155 68852 284156 68916
rect 284220 68852 284221 68916
rect 284155 68851 284221 68852
rect 284158 65620 284218 68851
rect 284526 65620 284586 181731
rect 284894 65620 284954 181867
rect 285262 65620 285322 182003
rect 285627 180164 285693 180165
rect 285627 180100 285628 180164
rect 285692 180100 285693 180164
rect 285627 180099 285693 180100
rect 285630 65620 285690 180099
rect 285998 65620 286058 182275
rect 286182 178941 286242 191523
rect 288019 189412 288085 189413
rect 288019 189348 288020 189412
rect 288084 189348 288085 189412
rect 288019 189347 288085 189348
rect 286363 186692 286429 186693
rect 286363 186628 286364 186692
rect 286428 186628 286429 186692
rect 286363 186627 286429 186628
rect 286366 182477 286426 186627
rect 288022 186557 288082 189347
rect 288019 186556 288085 186557
rect 288019 186492 288020 186556
rect 288084 186492 288085 186556
rect 288019 186491 288085 186492
rect 286547 184924 286613 184925
rect 286547 184860 286548 184924
rect 286612 184860 286613 184924
rect 286547 184859 286613 184860
rect 286363 182476 286429 182477
rect 286363 182412 286364 182476
rect 286428 182412 286429 182476
rect 286363 182411 286429 182412
rect 286179 178940 286245 178941
rect 286179 178876 286180 178940
rect 286244 178876 286245 178940
rect 286179 178875 286245 178876
rect 286366 65620 286426 182411
rect 286550 180029 286610 184859
rect 288019 183156 288085 183157
rect 288019 183092 288020 183156
rect 288084 183092 288085 183156
rect 288019 183091 288085 183092
rect 287835 183020 287901 183021
rect 287835 182956 287836 183020
rect 287900 182956 287901 183020
rect 287835 182955 287901 182956
rect 287467 182884 287533 182885
rect 287467 182820 287468 182884
rect 287532 182820 287533 182884
rect 287467 182819 287533 182820
rect 287099 182748 287165 182749
rect 287099 182684 287100 182748
rect 287164 182684 287165 182748
rect 287099 182683 287165 182684
rect 286547 180028 286613 180029
rect 286547 179964 286548 180028
rect 286612 179964 286613 180028
rect 286547 179963 286613 179964
rect 286731 177444 286797 177445
rect 286731 177380 286732 177444
rect 286796 177380 286797 177444
rect 286731 177379 286797 177380
rect 286734 65620 286794 177379
rect 287102 65620 287162 182683
rect 287470 65620 287530 182819
rect 287838 65620 287898 182955
rect 288022 65650 288082 183091
rect 288206 182613 288266 210291
rect 288390 183565 288450 606051
rect 289675 192540 289741 192541
rect 289675 192476 289676 192540
rect 289740 192476 289741 192540
rect 289675 192475 289741 192476
rect 288387 183564 288453 183565
rect 288387 183500 288388 183564
rect 288452 183500 288453 183564
rect 288387 183499 288453 183500
rect 289307 183564 289373 183565
rect 289307 183500 289308 183564
rect 289372 183500 289373 183564
rect 289307 183499 289373 183500
rect 288939 183428 289005 183429
rect 288939 183364 288940 183428
rect 289004 183364 289005 183428
rect 288939 183363 289005 183364
rect 288571 183292 288637 183293
rect 288571 183228 288572 183292
rect 288636 183228 288637 183292
rect 288571 183227 288637 183228
rect 288203 182612 288269 182613
rect 288203 182548 288204 182612
rect 288268 182548 288269 182612
rect 288203 182547 288269 182548
rect 288022 65590 288236 65650
rect 288574 65620 288634 183227
rect 288942 65620 289002 183363
rect 289310 65620 289370 183499
rect 289678 178125 289738 192475
rect 289859 189140 289925 189141
rect 289859 189076 289860 189140
rect 289924 189076 289925 189140
rect 289859 189075 289925 189076
rect 289862 179485 289922 189075
rect 290963 188460 291029 188461
rect 290963 188396 290964 188460
rect 291028 188396 291029 188460
rect 290963 188395 291029 188396
rect 290966 187781 291026 188395
rect 290963 187780 291029 187781
rect 290963 187716 290964 187780
rect 291028 187716 291029 187780
rect 290963 187715 291029 187716
rect 290411 183972 290477 183973
rect 290411 183908 290412 183972
rect 290476 183908 290477 183972
rect 290411 183907 290477 183908
rect 290043 183836 290109 183837
rect 290043 183772 290044 183836
rect 290108 183772 290109 183836
rect 290043 183771 290109 183772
rect 289859 179484 289925 179485
rect 289859 179420 289860 179484
rect 289924 179420 289925 179484
rect 289859 179419 289925 179420
rect 289675 178124 289741 178125
rect 289675 178060 289676 178124
rect 289740 178060 289741 178124
rect 289675 178059 289741 178060
rect 289675 177988 289741 177989
rect 289675 177924 289676 177988
rect 289740 177924 289741 177988
rect 289675 177923 289741 177924
rect 289678 65670 289738 177923
rect 290046 65620 290106 183771
rect 290414 65724 290474 183907
rect 290966 67013 291026 187715
rect 291150 184925 291210 658139
rect 307365 208174 307685 208206
rect 307365 207938 307407 208174
rect 307643 207938 307685 208174
rect 307365 207854 307685 207938
rect 307365 207618 307407 207854
rect 307643 207618 307685 207854
rect 307365 207586 307685 207618
rect 315207 208174 315527 208206
rect 315207 207938 315249 208174
rect 315485 207938 315527 208174
rect 315207 207854 315527 207938
rect 315207 207618 315249 207854
rect 315485 207618 315527 207854
rect 315207 207586 315527 207618
rect 323049 208174 323369 208206
rect 323049 207938 323091 208174
rect 323327 207938 323369 208174
rect 323049 207854 323369 207938
rect 323049 207618 323091 207854
rect 323327 207618 323369 207854
rect 323049 207586 323369 207618
rect 330891 208174 331211 208206
rect 330891 207938 330933 208174
rect 331169 207938 331211 208174
rect 330891 207854 331211 207938
rect 330891 207618 330933 207854
rect 331169 207618 331211 207854
rect 330891 207586 331211 207618
rect 341497 208174 341817 208206
rect 341497 207938 341539 208174
rect 341775 207938 341817 208174
rect 341497 207854 341817 207938
rect 341497 207618 341539 207854
rect 341775 207618 341817 207854
rect 341497 207586 341817 207618
rect 349339 208174 349659 208206
rect 349339 207938 349381 208174
rect 349617 207938 349659 208174
rect 349339 207854 349659 207938
rect 349339 207618 349381 207854
rect 349617 207618 349659 207854
rect 349339 207586 349659 207618
rect 357181 208174 357501 208206
rect 357181 207938 357223 208174
rect 357459 207938 357501 208174
rect 357181 207854 357501 207938
rect 357181 207618 357223 207854
rect 357459 207618 357501 207854
rect 357181 207586 357501 207618
rect 365023 208174 365343 208206
rect 365023 207938 365065 208174
rect 365301 207938 365343 208174
rect 365023 207854 365343 207938
rect 365023 207618 365065 207854
rect 365301 207618 365343 207854
rect 365023 207586 365343 207618
rect 375629 208174 375949 208206
rect 375629 207938 375671 208174
rect 375907 207938 375949 208174
rect 375629 207854 375949 207938
rect 375629 207618 375671 207854
rect 375907 207618 375949 207854
rect 375629 207586 375949 207618
rect 383471 208174 383791 208206
rect 383471 207938 383513 208174
rect 383749 207938 383791 208174
rect 383471 207854 383791 207938
rect 383471 207618 383513 207854
rect 383749 207618 383791 207854
rect 383471 207586 383791 207618
rect 391313 208174 391633 208206
rect 391313 207938 391355 208174
rect 391591 207938 391633 208174
rect 391313 207854 391633 207938
rect 391313 207618 391355 207854
rect 391591 207618 391633 207854
rect 391313 207586 391633 207618
rect 399155 208174 399475 208206
rect 399155 207938 399197 208174
rect 399433 207938 399475 208174
rect 399155 207854 399475 207938
rect 399155 207618 399197 207854
rect 399433 207618 399475 207854
rect 399155 207586 399475 207618
rect 409761 208174 410081 208206
rect 409761 207938 409803 208174
rect 410039 207938 410081 208174
rect 409761 207854 410081 207938
rect 409761 207618 409803 207854
rect 410039 207618 410081 207854
rect 409761 207586 410081 207618
rect 417603 208174 417923 208206
rect 417603 207938 417645 208174
rect 417881 207938 417923 208174
rect 417603 207854 417923 207938
rect 417603 207618 417645 207854
rect 417881 207618 417923 207854
rect 417603 207586 417923 207618
rect 425445 208174 425765 208206
rect 425445 207938 425487 208174
rect 425723 207938 425765 208174
rect 425445 207854 425765 207938
rect 425445 207618 425487 207854
rect 425723 207618 425765 207854
rect 425445 207586 425765 207618
rect 433287 208174 433607 208206
rect 433287 207938 433329 208174
rect 433565 207938 433607 208174
rect 433287 207854 433607 207938
rect 433287 207618 433329 207854
rect 433565 207618 433607 207854
rect 433287 207586 433607 207618
rect 443893 208174 444213 208206
rect 443893 207938 443935 208174
rect 444171 207938 444213 208174
rect 443893 207854 444213 207938
rect 443893 207618 443935 207854
rect 444171 207618 444213 207854
rect 443893 207586 444213 207618
rect 451735 208174 452055 208206
rect 451735 207938 451777 208174
rect 452013 207938 452055 208174
rect 451735 207854 452055 207938
rect 451735 207618 451777 207854
rect 452013 207618 452055 207854
rect 451735 207586 452055 207618
rect 459577 208174 459897 208206
rect 459577 207938 459619 208174
rect 459855 207938 459897 208174
rect 459577 207854 459897 207938
rect 459577 207618 459619 207854
rect 459855 207618 459897 207854
rect 459577 207586 459897 207618
rect 467419 208174 467739 208206
rect 467419 207938 467461 208174
rect 467697 207938 467739 208174
rect 467419 207854 467739 207938
rect 467419 207618 467461 207854
rect 467697 207618 467739 207854
rect 467419 207586 467739 207618
rect 478025 208174 478345 208206
rect 478025 207938 478067 208174
rect 478303 207938 478345 208174
rect 478025 207854 478345 207938
rect 478025 207618 478067 207854
rect 478303 207618 478345 207854
rect 478025 207586 478345 207618
rect 485867 208174 486187 208206
rect 485867 207938 485909 208174
rect 486145 207938 486187 208174
rect 485867 207854 486187 207938
rect 485867 207618 485909 207854
rect 486145 207618 486187 207854
rect 485867 207586 486187 207618
rect 493709 208174 494029 208206
rect 493709 207938 493751 208174
rect 493987 207938 494029 208174
rect 493709 207854 494029 207938
rect 493709 207618 493751 207854
rect 493987 207618 494029 207854
rect 493709 207586 494029 207618
rect 501551 208174 501871 208206
rect 501551 207938 501593 208174
rect 501829 207938 501871 208174
rect 501551 207854 501871 207938
rect 501551 207618 501593 207854
rect 501829 207618 501871 207854
rect 501551 207586 501871 207618
rect 512157 208174 512477 208206
rect 512157 207938 512199 208174
rect 512435 207938 512477 208174
rect 512157 207854 512477 207938
rect 512157 207618 512199 207854
rect 512435 207618 512477 207854
rect 512157 207586 512477 207618
rect 519999 208174 520319 208206
rect 519999 207938 520041 208174
rect 520277 207938 520319 208174
rect 519999 207854 520319 207938
rect 519999 207618 520041 207854
rect 520277 207618 520319 207854
rect 519999 207586 520319 207618
rect 527841 208174 528161 208206
rect 527841 207938 527883 208174
rect 528119 207938 528161 208174
rect 527841 207854 528161 207938
rect 527841 207618 527883 207854
rect 528119 207618 528161 207854
rect 527841 207586 528161 207618
rect 535683 208174 536003 208206
rect 535683 207938 535725 208174
rect 535961 207938 536003 208174
rect 535683 207854 536003 207938
rect 535683 207618 535725 207854
rect 535961 207618 536003 207854
rect 535683 207586 536003 207618
rect 546289 208174 546609 208206
rect 546289 207938 546331 208174
rect 546567 207938 546609 208174
rect 546289 207854 546609 207938
rect 546289 207618 546331 207854
rect 546567 207618 546609 207854
rect 546289 207586 546609 207618
rect 554131 208174 554451 208206
rect 554131 207938 554173 208174
rect 554409 207938 554451 208174
rect 554131 207854 554451 207938
rect 554131 207618 554173 207854
rect 554409 207618 554451 207854
rect 554131 207586 554451 207618
rect 561973 208174 562293 208206
rect 561973 207938 562015 208174
rect 562251 207938 562293 208174
rect 561973 207854 562293 207938
rect 561973 207618 562015 207854
rect 562251 207618 562293 207854
rect 561973 207586 562293 207618
rect 569815 208174 570135 208206
rect 569815 207938 569857 208174
rect 570093 207938 570135 208174
rect 569815 207854 570135 207938
rect 569815 207618 569857 207854
rect 570093 207618 570135 207854
rect 569815 207586 570135 207618
rect 303444 204454 303764 204486
rect 303444 204218 303486 204454
rect 303722 204218 303764 204454
rect 303444 204134 303764 204218
rect 303444 203898 303486 204134
rect 303722 203898 303764 204134
rect 303444 203866 303764 203898
rect 311286 204454 311606 204486
rect 311286 204218 311328 204454
rect 311564 204218 311606 204454
rect 311286 204134 311606 204218
rect 311286 203898 311328 204134
rect 311564 203898 311606 204134
rect 311286 203866 311606 203898
rect 319128 204454 319448 204486
rect 319128 204218 319170 204454
rect 319406 204218 319448 204454
rect 319128 204134 319448 204218
rect 319128 203898 319170 204134
rect 319406 203898 319448 204134
rect 319128 203866 319448 203898
rect 326970 204454 327290 204486
rect 326970 204218 327012 204454
rect 327248 204218 327290 204454
rect 326970 204134 327290 204218
rect 326970 203898 327012 204134
rect 327248 203898 327290 204134
rect 326970 203866 327290 203898
rect 337576 204454 337896 204486
rect 337576 204218 337618 204454
rect 337854 204218 337896 204454
rect 337576 204134 337896 204218
rect 337576 203898 337618 204134
rect 337854 203898 337896 204134
rect 337576 203866 337896 203898
rect 345418 204454 345738 204486
rect 345418 204218 345460 204454
rect 345696 204218 345738 204454
rect 345418 204134 345738 204218
rect 345418 203898 345460 204134
rect 345696 203898 345738 204134
rect 345418 203866 345738 203898
rect 353260 204454 353580 204486
rect 353260 204218 353302 204454
rect 353538 204218 353580 204454
rect 353260 204134 353580 204218
rect 353260 203898 353302 204134
rect 353538 203898 353580 204134
rect 353260 203866 353580 203898
rect 361102 204454 361422 204486
rect 361102 204218 361144 204454
rect 361380 204218 361422 204454
rect 361102 204134 361422 204218
rect 361102 203898 361144 204134
rect 361380 203898 361422 204134
rect 361102 203866 361422 203898
rect 371708 204454 372028 204486
rect 371708 204218 371750 204454
rect 371986 204218 372028 204454
rect 371708 204134 372028 204218
rect 371708 203898 371750 204134
rect 371986 203898 372028 204134
rect 371708 203866 372028 203898
rect 379550 204454 379870 204486
rect 379550 204218 379592 204454
rect 379828 204218 379870 204454
rect 379550 204134 379870 204218
rect 379550 203898 379592 204134
rect 379828 203898 379870 204134
rect 379550 203866 379870 203898
rect 387392 204454 387712 204486
rect 387392 204218 387434 204454
rect 387670 204218 387712 204454
rect 387392 204134 387712 204218
rect 387392 203898 387434 204134
rect 387670 203898 387712 204134
rect 387392 203866 387712 203898
rect 395234 204454 395554 204486
rect 395234 204218 395276 204454
rect 395512 204218 395554 204454
rect 395234 204134 395554 204218
rect 395234 203898 395276 204134
rect 395512 203898 395554 204134
rect 395234 203866 395554 203898
rect 405840 204454 406160 204486
rect 405840 204218 405882 204454
rect 406118 204218 406160 204454
rect 405840 204134 406160 204218
rect 405840 203898 405882 204134
rect 406118 203898 406160 204134
rect 405840 203866 406160 203898
rect 413682 204454 414002 204486
rect 413682 204218 413724 204454
rect 413960 204218 414002 204454
rect 413682 204134 414002 204218
rect 413682 203898 413724 204134
rect 413960 203898 414002 204134
rect 413682 203866 414002 203898
rect 421524 204454 421844 204486
rect 421524 204218 421566 204454
rect 421802 204218 421844 204454
rect 421524 204134 421844 204218
rect 421524 203898 421566 204134
rect 421802 203898 421844 204134
rect 421524 203866 421844 203898
rect 429366 204454 429686 204486
rect 429366 204218 429408 204454
rect 429644 204218 429686 204454
rect 429366 204134 429686 204218
rect 429366 203898 429408 204134
rect 429644 203898 429686 204134
rect 429366 203866 429686 203898
rect 439972 204454 440292 204486
rect 439972 204218 440014 204454
rect 440250 204218 440292 204454
rect 439972 204134 440292 204218
rect 439972 203898 440014 204134
rect 440250 203898 440292 204134
rect 439972 203866 440292 203898
rect 447814 204454 448134 204486
rect 447814 204218 447856 204454
rect 448092 204218 448134 204454
rect 447814 204134 448134 204218
rect 447814 203898 447856 204134
rect 448092 203898 448134 204134
rect 447814 203866 448134 203898
rect 455656 204454 455976 204486
rect 455656 204218 455698 204454
rect 455934 204218 455976 204454
rect 455656 204134 455976 204218
rect 455656 203898 455698 204134
rect 455934 203898 455976 204134
rect 455656 203866 455976 203898
rect 463498 204454 463818 204486
rect 463498 204218 463540 204454
rect 463776 204218 463818 204454
rect 463498 204134 463818 204218
rect 463498 203898 463540 204134
rect 463776 203898 463818 204134
rect 463498 203866 463818 203898
rect 474104 204454 474424 204486
rect 474104 204218 474146 204454
rect 474382 204218 474424 204454
rect 474104 204134 474424 204218
rect 474104 203898 474146 204134
rect 474382 203898 474424 204134
rect 474104 203866 474424 203898
rect 481946 204454 482266 204486
rect 481946 204218 481988 204454
rect 482224 204218 482266 204454
rect 481946 204134 482266 204218
rect 481946 203898 481988 204134
rect 482224 203898 482266 204134
rect 481946 203866 482266 203898
rect 489788 204454 490108 204486
rect 489788 204218 489830 204454
rect 490066 204218 490108 204454
rect 489788 204134 490108 204218
rect 489788 203898 489830 204134
rect 490066 203898 490108 204134
rect 489788 203866 490108 203898
rect 497630 204454 497950 204486
rect 497630 204218 497672 204454
rect 497908 204218 497950 204454
rect 497630 204134 497950 204218
rect 497630 203898 497672 204134
rect 497908 203898 497950 204134
rect 497630 203866 497950 203898
rect 508236 204454 508556 204486
rect 508236 204218 508278 204454
rect 508514 204218 508556 204454
rect 508236 204134 508556 204218
rect 508236 203898 508278 204134
rect 508514 203898 508556 204134
rect 508236 203866 508556 203898
rect 516078 204454 516398 204486
rect 516078 204218 516120 204454
rect 516356 204218 516398 204454
rect 516078 204134 516398 204218
rect 516078 203898 516120 204134
rect 516356 203898 516398 204134
rect 516078 203866 516398 203898
rect 523920 204454 524240 204486
rect 523920 204218 523962 204454
rect 524198 204218 524240 204454
rect 523920 204134 524240 204218
rect 523920 203898 523962 204134
rect 524198 203898 524240 204134
rect 523920 203866 524240 203898
rect 531762 204454 532082 204486
rect 531762 204218 531804 204454
rect 532040 204218 532082 204454
rect 531762 204134 532082 204218
rect 531762 203898 531804 204134
rect 532040 203898 532082 204134
rect 531762 203866 532082 203898
rect 542368 204454 542688 204486
rect 542368 204218 542410 204454
rect 542646 204218 542688 204454
rect 542368 204134 542688 204218
rect 542368 203898 542410 204134
rect 542646 203898 542688 204134
rect 542368 203866 542688 203898
rect 550210 204454 550530 204486
rect 550210 204218 550252 204454
rect 550488 204218 550530 204454
rect 550210 204134 550530 204218
rect 550210 203898 550252 204134
rect 550488 203898 550530 204134
rect 550210 203866 550530 203898
rect 558052 204454 558372 204486
rect 558052 204218 558094 204454
rect 558330 204218 558372 204454
rect 558052 204134 558372 204218
rect 558052 203898 558094 204134
rect 558330 203898 558372 204134
rect 558052 203866 558372 203898
rect 565894 204454 566214 204486
rect 565894 204218 565936 204454
rect 566172 204218 566214 204454
rect 565894 204134 566214 204218
rect 565894 203898 565936 204134
rect 566172 203898 566214 204134
rect 565894 203866 566214 203898
rect 307365 198174 307685 198206
rect 307365 197938 307407 198174
rect 307643 197938 307685 198174
rect 307365 197854 307685 197938
rect 307365 197618 307407 197854
rect 307643 197618 307685 197854
rect 307365 197586 307685 197618
rect 315207 198174 315527 198206
rect 315207 197938 315249 198174
rect 315485 197938 315527 198174
rect 315207 197854 315527 197938
rect 315207 197618 315249 197854
rect 315485 197618 315527 197854
rect 315207 197586 315527 197618
rect 323049 198174 323369 198206
rect 323049 197938 323091 198174
rect 323327 197938 323369 198174
rect 323049 197854 323369 197938
rect 323049 197618 323091 197854
rect 323327 197618 323369 197854
rect 323049 197586 323369 197618
rect 330891 198174 331211 198206
rect 330891 197938 330933 198174
rect 331169 197938 331211 198174
rect 330891 197854 331211 197938
rect 330891 197618 330933 197854
rect 331169 197618 331211 197854
rect 330891 197586 331211 197618
rect 341497 198174 341817 198206
rect 341497 197938 341539 198174
rect 341775 197938 341817 198174
rect 341497 197854 341817 197938
rect 341497 197618 341539 197854
rect 341775 197618 341817 197854
rect 341497 197586 341817 197618
rect 349339 198174 349659 198206
rect 349339 197938 349381 198174
rect 349617 197938 349659 198174
rect 349339 197854 349659 197938
rect 349339 197618 349381 197854
rect 349617 197618 349659 197854
rect 349339 197586 349659 197618
rect 357181 198174 357501 198206
rect 357181 197938 357223 198174
rect 357459 197938 357501 198174
rect 357181 197854 357501 197938
rect 357181 197618 357223 197854
rect 357459 197618 357501 197854
rect 357181 197586 357501 197618
rect 365023 198174 365343 198206
rect 365023 197938 365065 198174
rect 365301 197938 365343 198174
rect 365023 197854 365343 197938
rect 365023 197618 365065 197854
rect 365301 197618 365343 197854
rect 365023 197586 365343 197618
rect 375629 198174 375949 198206
rect 375629 197938 375671 198174
rect 375907 197938 375949 198174
rect 375629 197854 375949 197938
rect 375629 197618 375671 197854
rect 375907 197618 375949 197854
rect 375629 197586 375949 197618
rect 383471 198174 383791 198206
rect 383471 197938 383513 198174
rect 383749 197938 383791 198174
rect 383471 197854 383791 197938
rect 383471 197618 383513 197854
rect 383749 197618 383791 197854
rect 383471 197586 383791 197618
rect 391313 198174 391633 198206
rect 391313 197938 391355 198174
rect 391591 197938 391633 198174
rect 391313 197854 391633 197938
rect 391313 197618 391355 197854
rect 391591 197618 391633 197854
rect 391313 197586 391633 197618
rect 399155 198174 399475 198206
rect 399155 197938 399197 198174
rect 399433 197938 399475 198174
rect 399155 197854 399475 197938
rect 399155 197618 399197 197854
rect 399433 197618 399475 197854
rect 399155 197586 399475 197618
rect 409761 198174 410081 198206
rect 409761 197938 409803 198174
rect 410039 197938 410081 198174
rect 409761 197854 410081 197938
rect 409761 197618 409803 197854
rect 410039 197618 410081 197854
rect 409761 197586 410081 197618
rect 417603 198174 417923 198206
rect 417603 197938 417645 198174
rect 417881 197938 417923 198174
rect 417603 197854 417923 197938
rect 417603 197618 417645 197854
rect 417881 197618 417923 197854
rect 417603 197586 417923 197618
rect 425445 198174 425765 198206
rect 425445 197938 425487 198174
rect 425723 197938 425765 198174
rect 425445 197854 425765 197938
rect 425445 197618 425487 197854
rect 425723 197618 425765 197854
rect 425445 197586 425765 197618
rect 433287 198174 433607 198206
rect 433287 197938 433329 198174
rect 433565 197938 433607 198174
rect 433287 197854 433607 197938
rect 433287 197618 433329 197854
rect 433565 197618 433607 197854
rect 433287 197586 433607 197618
rect 443893 198174 444213 198206
rect 443893 197938 443935 198174
rect 444171 197938 444213 198174
rect 443893 197854 444213 197938
rect 443893 197618 443935 197854
rect 444171 197618 444213 197854
rect 443893 197586 444213 197618
rect 451735 198174 452055 198206
rect 451735 197938 451777 198174
rect 452013 197938 452055 198174
rect 451735 197854 452055 197938
rect 451735 197618 451777 197854
rect 452013 197618 452055 197854
rect 451735 197586 452055 197618
rect 459577 198174 459897 198206
rect 459577 197938 459619 198174
rect 459855 197938 459897 198174
rect 459577 197854 459897 197938
rect 459577 197618 459619 197854
rect 459855 197618 459897 197854
rect 459577 197586 459897 197618
rect 467419 198174 467739 198206
rect 467419 197938 467461 198174
rect 467697 197938 467739 198174
rect 467419 197854 467739 197938
rect 467419 197618 467461 197854
rect 467697 197618 467739 197854
rect 467419 197586 467739 197618
rect 478025 198174 478345 198206
rect 478025 197938 478067 198174
rect 478303 197938 478345 198174
rect 478025 197854 478345 197938
rect 478025 197618 478067 197854
rect 478303 197618 478345 197854
rect 478025 197586 478345 197618
rect 485867 198174 486187 198206
rect 485867 197938 485909 198174
rect 486145 197938 486187 198174
rect 485867 197854 486187 197938
rect 485867 197618 485909 197854
rect 486145 197618 486187 197854
rect 485867 197586 486187 197618
rect 493709 198174 494029 198206
rect 493709 197938 493751 198174
rect 493987 197938 494029 198174
rect 493709 197854 494029 197938
rect 493709 197618 493751 197854
rect 493987 197618 494029 197854
rect 493709 197586 494029 197618
rect 501551 198174 501871 198206
rect 501551 197938 501593 198174
rect 501829 197938 501871 198174
rect 501551 197854 501871 197938
rect 501551 197618 501593 197854
rect 501829 197618 501871 197854
rect 501551 197586 501871 197618
rect 512157 198174 512477 198206
rect 512157 197938 512199 198174
rect 512435 197938 512477 198174
rect 512157 197854 512477 197938
rect 512157 197618 512199 197854
rect 512435 197618 512477 197854
rect 512157 197586 512477 197618
rect 519999 198174 520319 198206
rect 519999 197938 520041 198174
rect 520277 197938 520319 198174
rect 519999 197854 520319 197938
rect 519999 197618 520041 197854
rect 520277 197618 520319 197854
rect 519999 197586 520319 197618
rect 527841 198174 528161 198206
rect 527841 197938 527883 198174
rect 528119 197938 528161 198174
rect 527841 197854 528161 197938
rect 527841 197618 527883 197854
rect 528119 197618 528161 197854
rect 527841 197586 528161 197618
rect 535683 198174 536003 198206
rect 535683 197938 535725 198174
rect 535961 197938 536003 198174
rect 535683 197854 536003 197938
rect 535683 197618 535725 197854
rect 535961 197618 536003 197854
rect 535683 197586 536003 197618
rect 546289 198174 546609 198206
rect 546289 197938 546331 198174
rect 546567 197938 546609 198174
rect 546289 197854 546609 197938
rect 546289 197618 546331 197854
rect 546567 197618 546609 197854
rect 546289 197586 546609 197618
rect 554131 198174 554451 198206
rect 554131 197938 554173 198174
rect 554409 197938 554451 198174
rect 554131 197854 554451 197938
rect 554131 197618 554173 197854
rect 554409 197618 554451 197854
rect 554131 197586 554451 197618
rect 561973 198174 562293 198206
rect 561973 197938 562015 198174
rect 562251 197938 562293 198174
rect 561973 197854 562293 197938
rect 561973 197618 562015 197854
rect 562251 197618 562293 197854
rect 561973 197586 562293 197618
rect 569815 198174 570135 198206
rect 569815 197938 569857 198174
rect 570093 197938 570135 198174
rect 569815 197854 570135 197938
rect 569815 197618 569857 197854
rect 570093 197618 570135 197854
rect 569815 197586 570135 197618
rect 303444 194454 303764 194486
rect 303444 194218 303486 194454
rect 303722 194218 303764 194454
rect 303444 194134 303764 194218
rect 303444 193898 303486 194134
rect 303722 193898 303764 194134
rect 303444 193866 303764 193898
rect 311286 194454 311606 194486
rect 311286 194218 311328 194454
rect 311564 194218 311606 194454
rect 311286 194134 311606 194218
rect 311286 193898 311328 194134
rect 311564 193898 311606 194134
rect 311286 193866 311606 193898
rect 319128 194454 319448 194486
rect 319128 194218 319170 194454
rect 319406 194218 319448 194454
rect 319128 194134 319448 194218
rect 319128 193898 319170 194134
rect 319406 193898 319448 194134
rect 319128 193866 319448 193898
rect 326970 194454 327290 194486
rect 326970 194218 327012 194454
rect 327248 194218 327290 194454
rect 326970 194134 327290 194218
rect 326970 193898 327012 194134
rect 327248 193898 327290 194134
rect 326970 193866 327290 193898
rect 337576 194454 337896 194486
rect 337576 194218 337618 194454
rect 337854 194218 337896 194454
rect 337576 194134 337896 194218
rect 337576 193898 337618 194134
rect 337854 193898 337896 194134
rect 337576 193866 337896 193898
rect 345418 194454 345738 194486
rect 345418 194218 345460 194454
rect 345696 194218 345738 194454
rect 345418 194134 345738 194218
rect 345418 193898 345460 194134
rect 345696 193898 345738 194134
rect 345418 193866 345738 193898
rect 353260 194454 353580 194486
rect 353260 194218 353302 194454
rect 353538 194218 353580 194454
rect 353260 194134 353580 194218
rect 353260 193898 353302 194134
rect 353538 193898 353580 194134
rect 353260 193866 353580 193898
rect 361102 194454 361422 194486
rect 361102 194218 361144 194454
rect 361380 194218 361422 194454
rect 361102 194134 361422 194218
rect 361102 193898 361144 194134
rect 361380 193898 361422 194134
rect 361102 193866 361422 193898
rect 371708 194454 372028 194486
rect 371708 194218 371750 194454
rect 371986 194218 372028 194454
rect 371708 194134 372028 194218
rect 371708 193898 371750 194134
rect 371986 193898 372028 194134
rect 371708 193866 372028 193898
rect 379550 194454 379870 194486
rect 379550 194218 379592 194454
rect 379828 194218 379870 194454
rect 379550 194134 379870 194218
rect 379550 193898 379592 194134
rect 379828 193898 379870 194134
rect 379550 193866 379870 193898
rect 387392 194454 387712 194486
rect 387392 194218 387434 194454
rect 387670 194218 387712 194454
rect 387392 194134 387712 194218
rect 387392 193898 387434 194134
rect 387670 193898 387712 194134
rect 387392 193866 387712 193898
rect 395234 194454 395554 194486
rect 395234 194218 395276 194454
rect 395512 194218 395554 194454
rect 395234 194134 395554 194218
rect 395234 193898 395276 194134
rect 395512 193898 395554 194134
rect 395234 193866 395554 193898
rect 405840 194454 406160 194486
rect 405840 194218 405882 194454
rect 406118 194218 406160 194454
rect 405840 194134 406160 194218
rect 405840 193898 405882 194134
rect 406118 193898 406160 194134
rect 405840 193866 406160 193898
rect 413682 194454 414002 194486
rect 413682 194218 413724 194454
rect 413960 194218 414002 194454
rect 413682 194134 414002 194218
rect 413682 193898 413724 194134
rect 413960 193898 414002 194134
rect 413682 193866 414002 193898
rect 421524 194454 421844 194486
rect 421524 194218 421566 194454
rect 421802 194218 421844 194454
rect 421524 194134 421844 194218
rect 421524 193898 421566 194134
rect 421802 193898 421844 194134
rect 421524 193866 421844 193898
rect 429366 194454 429686 194486
rect 429366 194218 429408 194454
rect 429644 194218 429686 194454
rect 429366 194134 429686 194218
rect 429366 193898 429408 194134
rect 429644 193898 429686 194134
rect 429366 193866 429686 193898
rect 439972 194454 440292 194486
rect 439972 194218 440014 194454
rect 440250 194218 440292 194454
rect 439972 194134 440292 194218
rect 439972 193898 440014 194134
rect 440250 193898 440292 194134
rect 439972 193866 440292 193898
rect 447814 194454 448134 194486
rect 447814 194218 447856 194454
rect 448092 194218 448134 194454
rect 447814 194134 448134 194218
rect 447814 193898 447856 194134
rect 448092 193898 448134 194134
rect 447814 193866 448134 193898
rect 455656 194454 455976 194486
rect 455656 194218 455698 194454
rect 455934 194218 455976 194454
rect 455656 194134 455976 194218
rect 455656 193898 455698 194134
rect 455934 193898 455976 194134
rect 455656 193866 455976 193898
rect 463498 194454 463818 194486
rect 463498 194218 463540 194454
rect 463776 194218 463818 194454
rect 463498 194134 463818 194218
rect 463498 193898 463540 194134
rect 463776 193898 463818 194134
rect 463498 193866 463818 193898
rect 474104 194454 474424 194486
rect 474104 194218 474146 194454
rect 474382 194218 474424 194454
rect 474104 194134 474424 194218
rect 474104 193898 474146 194134
rect 474382 193898 474424 194134
rect 474104 193866 474424 193898
rect 481946 194454 482266 194486
rect 481946 194218 481988 194454
rect 482224 194218 482266 194454
rect 481946 194134 482266 194218
rect 481946 193898 481988 194134
rect 482224 193898 482266 194134
rect 481946 193866 482266 193898
rect 489788 194454 490108 194486
rect 489788 194218 489830 194454
rect 490066 194218 490108 194454
rect 489788 194134 490108 194218
rect 489788 193898 489830 194134
rect 490066 193898 490108 194134
rect 489788 193866 490108 193898
rect 497630 194454 497950 194486
rect 497630 194218 497672 194454
rect 497908 194218 497950 194454
rect 497630 194134 497950 194218
rect 497630 193898 497672 194134
rect 497908 193898 497950 194134
rect 497630 193866 497950 193898
rect 508236 194454 508556 194486
rect 508236 194218 508278 194454
rect 508514 194218 508556 194454
rect 508236 194134 508556 194218
rect 508236 193898 508278 194134
rect 508514 193898 508556 194134
rect 508236 193866 508556 193898
rect 516078 194454 516398 194486
rect 516078 194218 516120 194454
rect 516356 194218 516398 194454
rect 516078 194134 516398 194218
rect 516078 193898 516120 194134
rect 516356 193898 516398 194134
rect 516078 193866 516398 193898
rect 523920 194454 524240 194486
rect 523920 194218 523962 194454
rect 524198 194218 524240 194454
rect 523920 194134 524240 194218
rect 523920 193898 523962 194134
rect 524198 193898 524240 194134
rect 523920 193866 524240 193898
rect 531762 194454 532082 194486
rect 531762 194218 531804 194454
rect 532040 194218 532082 194454
rect 531762 194134 532082 194218
rect 531762 193898 531804 194134
rect 532040 193898 532082 194134
rect 531762 193866 532082 193898
rect 542368 194454 542688 194486
rect 542368 194218 542410 194454
rect 542646 194218 542688 194454
rect 542368 194134 542688 194218
rect 542368 193898 542410 194134
rect 542646 193898 542688 194134
rect 542368 193866 542688 193898
rect 550210 194454 550530 194486
rect 550210 194218 550252 194454
rect 550488 194218 550530 194454
rect 550210 194134 550530 194218
rect 550210 193898 550252 194134
rect 550488 193898 550530 194134
rect 550210 193866 550530 193898
rect 558052 194454 558372 194486
rect 558052 194218 558094 194454
rect 558330 194218 558372 194454
rect 558052 194134 558372 194218
rect 558052 193898 558094 194134
rect 558330 193898 558372 194134
rect 558052 193866 558372 193898
rect 565894 194454 566214 194486
rect 565894 194218 565936 194454
rect 566172 194218 566214 194454
rect 565894 194134 566214 194218
rect 565894 193898 565936 194134
rect 566172 193898 566214 194134
rect 565894 193866 566214 193898
rect 298139 192268 298205 192269
rect 298139 192204 298140 192268
rect 298204 192204 298205 192268
rect 298139 192203 298205 192204
rect 295195 191996 295261 191997
rect 295195 191932 295196 191996
rect 295260 191932 295261 191996
rect 295195 191931 295261 191932
rect 295198 190909 295258 191931
rect 297955 191860 298021 191861
rect 297955 191796 297956 191860
rect 298020 191796 298021 191860
rect 297955 191795 298021 191796
rect 295195 190908 295261 190909
rect 295195 190844 295196 190908
rect 295260 190844 295261 190908
rect 295195 190843 295261 190844
rect 293171 188324 293237 188325
rect 293171 188260 293172 188324
rect 293236 188260 293237 188324
rect 293171 188259 293237 188260
rect 292435 187916 292501 187917
rect 292435 187852 292436 187916
rect 292500 187852 292501 187916
rect 292435 187851 292501 187852
rect 291331 185740 291397 185741
rect 291331 185676 291332 185740
rect 291396 185676 291397 185740
rect 291331 185675 291397 185676
rect 291147 184924 291213 184925
rect 291147 184860 291148 184924
rect 291212 184860 291213 184924
rect 291147 184859 291213 184860
rect 291334 184517 291394 185675
rect 291331 184516 291397 184517
rect 291331 184452 291332 184516
rect 291396 184452 291397 184516
rect 291331 184451 291397 184452
rect 291883 184244 291949 184245
rect 291883 184180 291884 184244
rect 291948 184180 291949 184244
rect 291883 184179 291949 184180
rect 291515 184108 291581 184109
rect 291515 184044 291516 184108
rect 291580 184044 291581 184108
rect 291515 184043 291581 184044
rect 290963 67012 291029 67013
rect 290963 66948 290964 67012
rect 291028 66948 291029 67012
rect 290963 66947 291029 66948
rect 291518 65620 291578 184043
rect 291886 65620 291946 184179
rect 292251 183700 292317 183701
rect 292251 183636 292252 183700
rect 292316 183636 292317 183700
rect 292251 183635 292317 183636
rect 292254 65620 292314 183635
rect 292438 179485 292498 187851
rect 293174 184789 293234 188259
rect 293539 188188 293605 188189
rect 293539 188124 293540 188188
rect 293604 188124 293605 188188
rect 293539 188123 293605 188124
rect 293171 184788 293237 184789
rect 293171 184724 293172 184788
rect 293236 184724 293237 184788
rect 293171 184723 293237 184724
rect 292987 184652 293053 184653
rect 292987 184588 292988 184652
rect 293052 184588 293053 184652
rect 292987 184587 293053 184588
rect 292619 184516 292685 184517
rect 292619 184452 292620 184516
rect 292684 184452 292685 184516
rect 292619 184451 292685 184452
rect 292435 179484 292501 179485
rect 292435 179420 292436 179484
rect 292500 179420 292501 179484
rect 292435 179419 292501 179420
rect 292622 65620 292682 184451
rect 292990 65620 293050 184587
rect 293542 179893 293602 188123
rect 295011 187780 295077 187781
rect 295011 187716 295012 187780
rect 295076 187716 295077 187780
rect 295011 187715 295077 187716
rect 293907 186148 293973 186149
rect 293907 186084 293908 186148
rect 293972 186084 293973 186148
rect 293907 186083 293973 186084
rect 293910 185061 293970 186083
rect 295014 185741 295074 187715
rect 295198 186013 295258 190843
rect 296299 190636 296365 190637
rect 296299 190572 296300 190636
rect 296364 190572 296365 190636
rect 296299 190571 296365 190572
rect 295195 186012 295261 186013
rect 295195 185948 295196 186012
rect 295260 185948 295261 186012
rect 295195 185947 295261 185948
rect 296302 185877 296362 190571
rect 297035 189548 297101 189549
rect 297035 189484 297036 189548
rect 297100 189484 297101 189548
rect 297035 189483 297101 189484
rect 297038 186149 297098 189483
rect 297958 186421 298018 191795
rect 298142 189277 298202 192203
rect 300899 190500 300965 190501
rect 300899 190436 300900 190500
rect 300964 190436 300965 190500
rect 300899 190435 300965 190436
rect 298691 189412 298757 189413
rect 298691 189348 298692 189412
rect 298756 189348 298757 189412
rect 298691 189347 298757 189348
rect 298139 189276 298205 189277
rect 298139 189212 298140 189276
rect 298204 189212 298205 189276
rect 298139 189211 298205 189212
rect 298694 186557 298754 189347
rect 299427 189140 299493 189141
rect 299427 189076 299428 189140
rect 299492 189076 299493 189140
rect 299427 189075 299493 189076
rect 299059 188052 299125 188053
rect 299059 187988 299060 188052
rect 299124 187988 299125 188052
rect 299059 187987 299125 187988
rect 298875 186828 298941 186829
rect 298875 186764 298876 186828
rect 298940 186764 298941 186828
rect 298875 186763 298941 186764
rect 298139 186556 298205 186557
rect 298139 186492 298140 186556
rect 298204 186492 298205 186556
rect 298139 186491 298205 186492
rect 298691 186556 298757 186557
rect 298691 186492 298692 186556
rect 298756 186492 298757 186556
rect 298691 186491 298757 186492
rect 297403 186420 297469 186421
rect 297403 186356 297404 186420
rect 297468 186356 297469 186420
rect 297403 186355 297469 186356
rect 297955 186420 298021 186421
rect 297955 186356 297956 186420
rect 298020 186356 298021 186420
rect 297955 186355 298021 186356
rect 297035 186148 297101 186149
rect 297035 186084 297036 186148
rect 297100 186084 297101 186148
rect 297035 186083 297101 186084
rect 296483 186012 296549 186013
rect 296483 185948 296484 186012
rect 296548 185948 296549 186012
rect 296483 185947 296549 185948
rect 296299 185876 296365 185877
rect 296299 185812 296300 185876
rect 296364 185812 296365 185876
rect 296299 185811 296365 185812
rect 295011 185740 295077 185741
rect 295011 185676 295012 185740
rect 295076 185676 295077 185740
rect 295011 185675 295077 185676
rect 294827 185332 294893 185333
rect 294827 185268 294828 185332
rect 294892 185268 294893 185332
rect 294827 185267 294893 185268
rect 294459 185196 294525 185197
rect 294459 185132 294460 185196
rect 294524 185132 294525 185196
rect 294459 185131 294525 185132
rect 293907 185060 293973 185061
rect 293907 184996 293908 185060
rect 293972 184996 293973 185060
rect 293907 184995 293973 184996
rect 293723 184924 293789 184925
rect 293723 184860 293724 184924
rect 293788 184860 293789 184924
rect 293723 184859 293789 184860
rect 293539 179892 293605 179893
rect 293539 179828 293540 179892
rect 293604 179828 293605 179892
rect 293539 179827 293605 179828
rect 293355 68916 293421 68917
rect 293355 68852 293356 68916
rect 293420 68852 293421 68916
rect 293355 68851 293421 68852
rect 293358 65620 293418 68851
rect 293726 65620 293786 184859
rect 293910 180810 293970 184995
rect 293910 180750 294154 180810
rect 294094 65620 294154 180750
rect 294462 65620 294522 185131
rect 294830 65620 294890 185267
rect 295014 180810 295074 185675
rect 295931 185604 295997 185605
rect 295931 185540 295932 185604
rect 295996 185540 295997 185604
rect 295931 185539 295997 185540
rect 295563 185468 295629 185469
rect 295563 185404 295564 185468
rect 295628 185404 295629 185468
rect 295563 185403 295629 185404
rect 295014 180750 295258 180810
rect 295198 65620 295258 180750
rect 295566 65620 295626 185403
rect 295934 65620 295994 185539
rect 296115 180164 296181 180165
rect 296115 180100 296116 180164
rect 296180 180100 296181 180164
rect 296115 180099 296181 180100
rect 296118 177989 296178 180099
rect 296115 177988 296181 177989
rect 296115 177924 296116 177988
rect 296180 177924 296181 177988
rect 296115 177923 296181 177924
rect 296302 65620 296362 185811
rect 296486 180165 296546 185947
rect 296851 180844 296917 180845
rect 296851 180780 296852 180844
rect 296916 180780 296917 180844
rect 296851 180779 296917 180780
rect 296483 180164 296549 180165
rect 296483 180100 296484 180164
rect 296548 180100 296549 180164
rect 296483 180099 296549 180100
rect 296854 179890 296914 180779
rect 296486 179830 296914 179890
rect 296486 66330 296546 179830
rect 296486 66270 296730 66330
rect 296670 65620 296730 66270
rect 297038 65620 297098 186083
rect 297406 65620 297466 186355
rect 297958 180810 298018 186355
rect 297774 180750 298018 180810
rect 297774 65620 297834 180750
rect 298142 65620 298202 186491
rect 298507 68644 298573 68645
rect 298507 68580 298508 68644
rect 298572 68580 298573 68644
rect 298507 68579 298573 68580
rect 298510 65620 298570 68579
rect 298878 65620 298938 186763
rect 299062 179485 299122 187987
rect 299243 187780 299309 187781
rect 299243 187716 299244 187780
rect 299308 187716 299309 187780
rect 299243 187715 299309 187716
rect 299246 187370 299306 187715
rect 299430 187645 299490 189075
rect 299611 188460 299677 188461
rect 299611 188396 299612 188460
rect 299676 188396 299677 188460
rect 299611 188395 299677 188396
rect 299614 187781 299674 188395
rect 299611 187780 299677 187781
rect 299611 187716 299612 187780
rect 299676 187716 299677 187780
rect 299611 187715 299677 187716
rect 299427 187644 299493 187645
rect 299427 187580 299428 187644
rect 299492 187580 299493 187644
rect 299427 187579 299493 187580
rect 300902 187509 300962 190435
rect 303570 190400 303630 191044
rect 304306 190400 304366 191080
rect 305042 190400 305102 191420
rect 305778 190400 305838 191420
rect 306514 190400 306574 191044
rect 307250 190400 307310 191044
rect 307986 190400 308046 191044
rect 308722 190400 308782 191044
rect 309458 190400 309518 191044
rect 310194 190400 310254 191044
rect 310930 190400 310990 191044
rect 311666 190400 311726 191080
rect 312402 190400 312462 191080
rect 313138 190400 313198 191080
rect 313874 190400 313934 191080
rect 314610 190400 314670 191080
rect 315346 190400 315406 191080
rect 316082 190400 316142 191080
rect 316818 190400 316878 191080
rect 317554 190400 317614 191080
rect 318290 190400 318350 191420
rect 319026 190400 319086 191080
rect 319762 190400 319822 191420
rect 320498 190400 320558 191420
rect 321234 190400 321294 191080
rect 321970 190400 322030 191080
rect 322706 190400 322766 191420
rect 323442 190400 323502 191080
rect 324178 190400 324238 191420
rect 324914 190400 324974 191080
rect 325650 190400 325710 191420
rect 326386 190400 326446 191420
rect 327122 190400 327182 191080
rect 327858 190400 327918 191080
rect 328594 190400 328654 191080
rect 329330 190400 329390 191080
rect 330066 190400 330126 191080
rect 330802 190400 330862 191080
rect 331538 190400 331598 191080
rect 332274 190770 332334 191420
rect 332274 190710 332426 190770
rect 332366 190470 332426 190710
rect 332274 190410 332426 190470
rect 332274 190400 332334 190410
rect 333010 190400 333070 191080
rect 333746 190400 333806 191080
rect 334482 190770 334542 191420
rect 334482 190710 334634 190770
rect 334574 190470 334634 190710
rect 334482 190410 334634 190470
rect 334482 190400 334542 190410
rect 337702 190400 337762 191044
rect 338438 190060 338498 191080
rect 339174 190400 339234 191420
rect 339910 190400 339970 191420
rect 340646 190400 340706 191044
rect 341382 190400 341442 191044
rect 342118 190060 342178 191044
rect 342854 190060 342914 191044
rect 343590 190400 343650 191044
rect 344326 190060 344386 191044
rect 345062 190400 345122 191044
rect 345798 190060 345858 191080
rect 346534 190400 346594 191080
rect 347270 190060 347330 191080
rect 348006 190060 348066 191080
rect 348742 190060 348802 191080
rect 349478 190400 349538 191080
rect 350214 190060 350274 191080
rect 350950 190400 351010 191080
rect 351686 190400 351746 191080
rect 352422 190400 352482 191420
rect 353158 190400 353218 191080
rect 353894 190400 353954 191420
rect 354660 191390 354874 191450
rect 354814 190470 354874 191390
rect 354630 190410 354874 190470
rect 354630 190400 354690 190410
rect 355366 190400 355426 191080
rect 356102 190400 356162 191080
rect 356838 190400 356898 191420
rect 357574 190400 357634 191080
rect 358310 190400 358370 191420
rect 359046 190400 359106 191080
rect 359782 190400 359842 191420
rect 360518 190400 360578 191420
rect 361254 190400 361314 191080
rect 361990 190400 362050 191080
rect 362726 190060 362786 191080
rect 363462 190400 363522 191080
rect 364198 190400 364258 191080
rect 364934 190400 364994 191080
rect 365670 190400 365730 191080
rect 366406 190400 366466 191420
rect 367142 190400 367202 191080
rect 367878 190400 367938 191080
rect 368614 190400 368674 191420
rect 371834 190400 371894 191044
rect 372570 190400 372630 191080
rect 373306 190770 373366 191420
rect 373214 190710 373366 190770
rect 374042 190770 374102 191420
rect 374042 190710 374194 190770
rect 373214 190470 373274 190710
rect 374134 190470 374194 190710
rect 373214 190410 373366 190470
rect 373306 190400 373366 190410
rect 374042 190410 374194 190470
rect 374042 190400 374102 190410
rect 374778 190400 374838 191044
rect 375514 190400 375574 191044
rect 376250 190400 376310 191044
rect 376986 190400 377046 191044
rect 377722 190400 377782 191044
rect 378458 190400 378518 191044
rect 379194 190400 379254 191044
rect 379930 190400 379990 191080
rect 380666 190400 380726 191080
rect 381402 190400 381462 191080
rect 382138 190400 382198 191080
rect 382874 190400 382934 191080
rect 383610 190400 383670 191080
rect 384346 190400 384406 191080
rect 385082 190400 385142 191080
rect 385818 190400 385878 191080
rect 386554 190400 386614 191420
rect 387290 190400 387350 191080
rect 388026 190400 388086 191420
rect 388762 190400 388822 191420
rect 389498 190400 389558 191080
rect 390234 190400 390294 191080
rect 390970 190400 391030 191420
rect 391706 190400 391766 191080
rect 392442 190400 392502 191420
rect 393178 190400 393238 191080
rect 393914 190400 393974 191420
rect 394650 190400 394710 191420
rect 395386 190400 395446 191080
rect 396122 190400 396182 191080
rect 396858 190400 396918 191080
rect 397594 190400 397654 191080
rect 398330 190400 398390 191080
rect 399066 190400 399126 191080
rect 399802 190400 399862 191080
rect 400538 190400 400598 191420
rect 401274 190400 401334 191080
rect 402010 190400 402070 191080
rect 402746 190400 402806 191420
rect 405966 190400 406026 191044
rect 406702 190060 406762 191080
rect 407438 190060 407498 191420
rect 408174 190060 408234 191420
rect 408910 190060 408970 191044
rect 409646 190060 409706 191044
rect 410382 190060 410442 191044
rect 411118 190400 411178 191044
rect 411854 190060 411914 191044
rect 412590 190060 412650 191044
rect 413326 190060 413386 191044
rect 414062 190060 414122 191080
rect 414798 190060 414858 191080
rect 415534 190400 415594 191080
rect 416270 190400 416330 191080
rect 417006 190400 417066 191080
rect 417742 190400 417802 191080
rect 418478 190400 418538 191080
rect 419214 190400 419274 191080
rect 419950 190400 420010 191080
rect 420686 190400 420746 191420
rect 421422 190400 421482 191080
rect 422158 190400 422218 191420
rect 422894 190400 422954 191420
rect 423630 190400 423690 191080
rect 424366 190400 424426 191080
rect 425102 190400 425162 191420
rect 425838 190400 425898 191080
rect 426574 190400 426634 191420
rect 427310 190400 427370 191080
rect 428046 190400 428106 191420
rect 428782 190400 428842 191420
rect 429518 190400 429578 191080
rect 430254 190400 430314 191080
rect 430990 190400 431050 191080
rect 431726 190400 431786 191080
rect 432462 190400 432522 191080
rect 433198 190400 433258 191080
rect 433934 190400 433994 191080
rect 434670 190400 434730 191420
rect 435406 190400 435466 191080
rect 436142 190400 436202 191080
rect 436878 190400 436938 191420
rect 440098 190400 440158 191044
rect 440834 190400 440894 191080
rect 441570 190770 441630 191420
rect 442306 190770 442366 191420
rect 441570 190710 441722 190770
rect 442306 190710 442458 190770
rect 441662 190470 441722 190710
rect 442398 190470 442458 190710
rect 441570 190410 441722 190470
rect 442306 190410 442458 190470
rect 441570 190400 441630 190410
rect 442306 190400 442366 190410
rect 443042 190400 443102 191044
rect 443778 190400 443838 191044
rect 444514 190400 444574 191044
rect 445250 190400 445310 191044
rect 445986 190400 446046 191044
rect 446722 190400 446782 191044
rect 447458 190400 447518 191044
rect 448194 190400 448254 191080
rect 448930 190400 448990 191080
rect 449666 190400 449726 191080
rect 450402 190400 450462 191080
rect 451138 190400 451198 191080
rect 451874 190400 451934 191080
rect 452610 190400 452670 191080
rect 453346 190400 453406 191080
rect 454082 190400 454142 191080
rect 454818 190400 454878 191420
rect 455554 190400 455614 191080
rect 456290 190400 456350 191420
rect 457026 190400 457086 191420
rect 457762 190400 457822 191080
rect 458498 190400 458558 191080
rect 459234 190400 459294 191420
rect 459970 190400 460030 191080
rect 460706 190400 460766 191420
rect 461442 190400 461502 191080
rect 462178 190400 462238 191420
rect 462914 190400 462974 191420
rect 463650 190400 463710 191080
rect 464386 190400 464446 191080
rect 465122 190400 465182 191080
rect 465858 190400 465918 191080
rect 466594 190400 466654 191080
rect 467330 190400 467390 191080
rect 468066 190400 468126 191080
rect 468802 190770 468862 191420
rect 468802 190710 468954 190770
rect 468894 190470 468954 190710
rect 468802 190410 468954 190470
rect 468802 190400 468862 190410
rect 469538 190400 469598 191080
rect 470274 190400 470334 191080
rect 471010 190770 471070 191420
rect 470918 190710 471070 190770
rect 470918 190470 470978 190710
rect 470918 190410 471070 190470
rect 471010 190400 471070 190410
rect 474230 190400 474290 191044
rect 474966 190060 475026 191080
rect 475702 190060 475762 191420
rect 476438 190060 476498 191420
rect 477174 190400 477234 191044
rect 477910 190060 477970 191044
rect 478646 190400 478706 191044
rect 479382 190400 479442 191044
rect 480118 190060 480178 191044
rect 480854 190060 480914 191044
rect 481590 190400 481650 191044
rect 482326 190060 482386 191080
rect 483062 190060 483122 191080
rect 483798 190060 483858 191080
rect 484534 190060 484594 191080
rect 485270 190400 485330 191080
rect 486006 190060 486066 191080
rect 486742 190400 486802 191080
rect 487478 190060 487538 191080
rect 488214 190400 488274 191080
rect 488950 190400 489010 191420
rect 489686 190400 489746 191080
rect 490422 190400 490482 191420
rect 491158 190400 491218 191420
rect 491894 190400 491954 191080
rect 492630 190400 492690 191080
rect 493366 190400 493426 191420
rect 494102 190400 494162 191080
rect 494838 190060 494898 191420
rect 495574 190400 495634 191080
rect 496310 190060 496370 191420
rect 497046 190400 497106 191420
rect 497782 190400 497842 191080
rect 498518 190400 498578 191080
rect 499254 190400 499314 191080
rect 499990 190060 500050 191080
rect 500726 190400 500786 191080
rect 501462 190060 501522 191080
rect 502198 190400 502258 191080
rect 502934 190400 502994 191420
rect 503670 190400 503730 191080
rect 504406 190400 504466 191080
rect 505142 190060 505202 191420
rect 508362 190400 508422 191044
rect 509098 190400 509158 191080
rect 509834 190400 509894 191420
rect 510570 190400 510630 191420
rect 511306 190400 511366 191044
rect 512042 190400 512102 191044
rect 512778 190400 512838 191044
rect 513514 190400 513574 191044
rect 514250 190400 514310 191044
rect 514986 190400 515046 191044
rect 515722 190400 515782 191044
rect 516458 190400 516518 191080
rect 517194 190400 517254 191080
rect 517930 190400 517990 191080
rect 518666 190400 518726 191080
rect 519402 190400 519462 191080
rect 520138 190400 520198 191080
rect 520874 190400 520934 191080
rect 521610 190400 521670 191080
rect 522346 190400 522406 191080
rect 523082 190400 523142 191420
rect 523818 190400 523878 191080
rect 524554 190400 524614 191420
rect 525290 190400 525350 191420
rect 526026 190400 526086 191080
rect 526762 190400 526822 191080
rect 527498 190400 527558 191420
rect 528234 190400 528294 191080
rect 528970 190400 529030 191420
rect 529706 190400 529766 191080
rect 530442 190400 530502 191420
rect 531178 190400 531238 191420
rect 531914 190400 531974 191080
rect 532650 190400 532710 191080
rect 533386 190400 533446 191080
rect 534122 190400 534182 191080
rect 534858 190400 534918 191080
rect 535594 190400 535654 191080
rect 536330 190400 536390 191080
rect 537066 190400 537126 191420
rect 537802 190400 537862 191080
rect 538538 190400 538598 191080
rect 539274 190400 539334 191420
rect 542494 190400 542554 191044
rect 543230 190400 543290 191080
rect 543966 190060 544026 191420
rect 544702 190060 544762 191420
rect 545438 190060 545498 191044
rect 546174 190400 546234 191044
rect 546910 190060 546970 191044
rect 547646 190060 547706 191044
rect 548382 190060 548442 191044
rect 549118 190400 549178 191044
rect 549854 190060 549914 191044
rect 550590 190060 550650 191080
rect 551326 190060 551386 191080
rect 552062 190060 552122 191080
rect 552798 190400 552858 191080
rect 553534 190400 553594 191080
rect 554270 190400 554330 191080
rect 555006 190060 555066 191080
rect 555742 190060 555802 191080
rect 556478 190400 556538 191080
rect 557214 190400 557274 191420
rect 557950 190400 558010 191080
rect 558686 190400 558746 191420
rect 559422 190400 559482 191420
rect 560158 190400 560218 191080
rect 560894 190400 560954 191080
rect 561630 190400 561690 191420
rect 562366 190400 562426 191080
rect 563102 190400 563162 191420
rect 563838 190400 563898 191080
rect 564574 190400 564634 191420
rect 565310 190400 565370 191420
rect 566046 190400 566106 191080
rect 566782 190400 566842 191080
rect 567518 190400 567578 191080
rect 568254 190400 568314 191080
rect 568990 190400 569050 191080
rect 569726 190400 569786 191080
rect 570462 190400 570522 191080
rect 571198 190400 571258 191420
rect 571934 190400 571994 191080
rect 572670 190400 572730 191080
rect 573406 190400 573466 191420
rect 301451 189276 301517 189277
rect 301451 189212 301452 189276
rect 301516 189212 301517 189276
rect 301451 189211 301517 189212
rect 301267 189140 301333 189141
rect 301267 189076 301268 189140
rect 301332 189076 301333 189140
rect 301267 189075 301333 189076
rect 301083 188324 301149 188325
rect 301083 188260 301084 188324
rect 301148 188260 301149 188324
rect 301083 188259 301149 188260
rect 300899 187508 300965 187509
rect 300899 187444 300900 187508
rect 300964 187444 300965 187508
rect 300899 187443 300965 187444
rect 300899 187372 300965 187373
rect 299246 187310 299490 187370
rect 299243 186964 299309 186965
rect 299243 186900 299244 186964
rect 299308 186900 299309 186964
rect 299243 186899 299309 186900
rect 299059 179484 299125 179485
rect 299059 179420 299060 179484
rect 299124 179420 299125 179484
rect 299059 179419 299125 179420
rect 299059 176764 299125 176765
rect 299059 176700 299060 176764
rect 299124 176700 299125 176764
rect 299059 176699 299125 176700
rect 299062 157453 299122 176699
rect 299059 157452 299125 157453
rect 299059 157388 299060 157452
rect 299124 157388 299125 157452
rect 299059 157387 299125 157388
rect 299246 65620 299306 186899
rect 299430 185469 299490 187310
rect 300899 187308 300900 187372
rect 300964 187308 300965 187372
rect 300899 187307 300965 187308
rect 299979 187236 300045 187237
rect 299979 187172 299980 187236
rect 300044 187172 300045 187236
rect 299979 187171 300045 187172
rect 299611 186692 299677 186693
rect 299611 186628 299612 186692
rect 299676 186628 299677 186692
rect 299611 186627 299677 186628
rect 299427 185468 299493 185469
rect 299427 185404 299428 185468
rect 299492 185404 299493 185468
rect 299427 185403 299493 185404
rect 299614 182477 299674 186627
rect 299795 185740 299861 185741
rect 299795 185676 299796 185740
rect 299860 185676 299861 185740
rect 299795 185675 299861 185676
rect 299611 182476 299677 182477
rect 299611 182412 299612 182476
rect 299676 182412 299677 182476
rect 299611 182411 299677 182412
rect 299798 180810 299858 185675
rect 299614 180750 299858 180810
rect 299614 65620 299674 180750
rect 299982 65620 300042 187171
rect 300902 181930 300962 187307
rect 301086 184789 301146 188259
rect 301270 186693 301330 189075
rect 301454 187373 301514 189211
rect 337147 188174 337467 188206
rect 337147 187938 337189 188174
rect 337425 187938 337467 188174
rect 337147 187854 337467 187938
rect 337147 187618 337189 187854
rect 337425 187618 337467 187854
rect 337147 187586 337467 187618
rect 404744 188174 405064 188206
rect 404744 187938 404786 188174
rect 405022 187938 405064 188174
rect 404744 187854 405064 187938
rect 404744 187618 404786 187854
rect 405022 187618 405064 187854
rect 404744 187586 405064 187618
rect 472341 188174 472661 188206
rect 472341 187938 472383 188174
rect 472619 187938 472661 188174
rect 472341 187854 472661 187938
rect 472341 187618 472383 187854
rect 472619 187618 472661 187854
rect 472341 187586 472661 187618
rect 539938 188174 540258 188206
rect 539938 187938 539980 188174
rect 540216 187938 540258 188174
rect 539938 187854 540258 187938
rect 539938 187618 539980 187854
rect 540216 187618 540258 187854
rect 539938 187586 540258 187618
rect 301451 187372 301517 187373
rect 301451 187308 301452 187372
rect 301516 187308 301517 187372
rect 301451 187307 301517 187308
rect 301267 186692 301333 186693
rect 301267 186628 301268 186692
rect 301332 186628 301333 186692
rect 301267 186627 301333 186628
rect 301083 184788 301149 184789
rect 301083 184724 301084 184788
rect 301148 184724 301149 184788
rect 301083 184723 301149 184724
rect 301270 184650 301330 186627
rect 300718 181870 300962 181930
rect 301086 184590 301330 184650
rect 300531 179892 300597 179893
rect 300531 179828 300532 179892
rect 300596 179828 300597 179892
rect 300531 179827 300597 179828
rect 300534 178805 300594 179827
rect 300163 178804 300229 178805
rect 300163 178740 300164 178804
rect 300228 178740 300229 178804
rect 300163 178739 300229 178740
rect 300531 178804 300597 178805
rect 300531 178740 300532 178804
rect 300596 178740 300597 178804
rect 300531 178739 300597 178740
rect 300166 157453 300226 178739
rect 300718 161490 300778 181870
rect 300899 181388 300965 181389
rect 300899 181324 300900 181388
rect 300964 181324 300965 181388
rect 300899 181323 300965 181324
rect 300902 180437 300962 181323
rect 300899 180436 300965 180437
rect 300899 180372 300900 180436
rect 300964 180372 300965 180436
rect 300899 180371 300965 180372
rect 301086 176765 301146 184590
rect 303349 184454 303669 184486
rect 303349 184218 303391 184454
rect 303627 184218 303669 184454
rect 303349 184134 303669 184218
rect 303349 183898 303391 184134
rect 303627 183898 303669 184134
rect 303349 183866 303669 183898
rect 370946 184454 371266 184486
rect 370946 184218 370988 184454
rect 371224 184218 371266 184454
rect 370946 184134 371266 184218
rect 370946 183898 370988 184134
rect 371224 183898 371266 184134
rect 370946 183866 371266 183898
rect 438543 184454 438863 184486
rect 438543 184218 438585 184454
rect 438821 184218 438863 184454
rect 438543 184134 438863 184218
rect 438543 183898 438585 184134
rect 438821 183898 438863 184134
rect 438543 183866 438863 183898
rect 506140 184454 506460 184486
rect 506140 184218 506182 184454
rect 506418 184218 506460 184454
rect 506140 184134 506460 184218
rect 506140 183898 506182 184134
rect 506418 183898 506460 184134
rect 506140 183866 506460 183898
rect 301267 182612 301333 182613
rect 301267 182548 301268 182612
rect 301332 182548 301333 182612
rect 301267 182547 301333 182548
rect 301270 177445 301330 182547
rect 302371 180028 302437 180029
rect 302371 179964 302372 180028
rect 302436 179964 302437 180028
rect 302371 179963 302437 179964
rect 302374 179890 302434 179963
rect 302374 179830 302618 179890
rect 302371 179484 302437 179485
rect 302371 179420 302372 179484
rect 302436 179420 302437 179484
rect 302371 179419 302437 179420
rect 301635 179348 301701 179349
rect 301635 179284 301636 179348
rect 301700 179284 301701 179348
rect 301635 179283 301701 179284
rect 301267 177444 301333 177445
rect 301267 177380 301268 177444
rect 301332 177380 301333 177444
rect 301267 177379 301333 177380
rect 301451 177308 301517 177309
rect 301451 177244 301452 177308
rect 301516 177244 301517 177308
rect 301451 177243 301517 177244
rect 301083 176764 301149 176765
rect 301083 176700 301084 176764
rect 301148 176700 301149 176764
rect 301083 176699 301149 176700
rect 300534 161430 300778 161490
rect 300163 157452 300229 157453
rect 300163 157388 300164 157452
rect 300228 157388 300229 157452
rect 300163 157387 300229 157388
rect 300534 156637 300594 161430
rect 300531 156636 300597 156637
rect 300531 156572 300532 156636
rect 300596 156572 300597 156636
rect 300531 156571 300597 156572
rect 300715 74628 300781 74629
rect 300715 74564 300716 74628
rect 300780 74564 300781 74628
rect 300715 74563 300781 74564
rect 300347 68780 300413 68781
rect 300347 68716 300348 68780
rect 300412 68716 300413 68780
rect 300347 68715 300413 68716
rect 300350 65620 300410 68715
rect 300718 65620 300778 74563
rect 301454 68917 301514 177243
rect 301638 158133 301698 179283
rect 301635 158132 301701 158133
rect 301635 158068 301636 158132
rect 301700 158068 301701 158132
rect 301635 158067 301701 158068
rect 301819 74764 301885 74765
rect 301819 74700 301820 74764
rect 301884 74700 301885 74764
rect 301819 74699 301885 74700
rect 301083 68916 301149 68917
rect 301083 68852 301084 68916
rect 301148 68852 301149 68916
rect 301083 68851 301149 68852
rect 301451 68916 301517 68917
rect 301451 68852 301452 68916
rect 301516 68852 301517 68916
rect 301451 68851 301517 68852
rect 301086 65620 301146 68851
rect 301451 67012 301517 67013
rect 301451 66948 301452 67012
rect 301516 66948 301517 67012
rect 301451 66947 301517 66948
rect 301454 65620 301514 66947
rect 301822 65620 301882 74699
rect 302374 65650 302434 179419
rect 302558 171150 302618 179830
rect 303570 178876 303630 179520
rect 304306 178840 304366 179520
rect 305042 178500 305102 179520
rect 305778 178500 305838 179520
rect 306514 178876 306574 179520
rect 307250 178876 307310 179520
rect 307986 178876 308046 179520
rect 308722 178876 308782 179520
rect 309458 178876 309518 179520
rect 310194 178876 310254 179520
rect 310930 178876 310990 179520
rect 311666 178840 311726 179520
rect 312402 178840 312462 179520
rect 313138 178840 313198 179520
rect 313874 178840 313934 179520
rect 314610 178840 314670 179520
rect 315346 178840 315406 179520
rect 316082 178840 316142 179520
rect 316818 178840 316878 179520
rect 317554 178840 317614 179520
rect 318290 178500 318350 179520
rect 319026 178840 319086 179520
rect 319762 178500 319822 179520
rect 320498 178500 320558 179520
rect 321234 178840 321294 179520
rect 321970 178840 322030 179520
rect 322706 178500 322766 179520
rect 323442 178840 323502 179520
rect 324178 178500 324238 179520
rect 324914 178840 324974 179520
rect 325650 178500 325710 179520
rect 326386 178500 326446 179520
rect 327122 178840 327182 179520
rect 327858 178840 327918 179520
rect 328594 178840 328654 179520
rect 329330 178840 329390 179520
rect 330066 178840 330126 179520
rect 330802 178840 330862 179520
rect 331538 178840 331598 179520
rect 332274 178500 332334 179520
rect 333010 178840 333070 179520
rect 333746 178840 333806 179520
rect 334482 178500 334542 179520
rect 337702 178876 337762 179520
rect 338438 178840 338498 179520
rect 334755 178804 334821 178805
rect 334755 178740 334756 178804
rect 334820 178740 334821 178804
rect 334755 178739 334821 178740
rect 307365 177879 307685 177936
rect 307365 177643 307407 177879
rect 307643 177643 307685 177879
rect 307365 177586 307685 177643
rect 315207 177879 315527 177936
rect 315207 177643 315249 177879
rect 315485 177643 315527 177879
rect 315207 177586 315527 177643
rect 323049 177879 323369 177936
rect 323049 177643 323091 177879
rect 323327 177643 323369 177879
rect 323049 177586 323369 177643
rect 330891 177879 331211 177936
rect 330891 177643 330933 177879
rect 331169 177643 331211 177879
rect 330891 177586 331211 177643
rect 303107 174588 303173 174589
rect 303107 174524 303108 174588
rect 303172 174524 303173 174588
rect 303107 174523 303173 174524
rect 302558 171090 302802 171150
rect 302742 157181 302802 171090
rect 302739 157180 302805 157181
rect 302739 157116 302740 157180
rect 302804 157116 302805 157180
rect 302739 157115 302805 157116
rect 303110 74550 303170 174523
rect 303444 174454 303764 174486
rect 303444 174218 303486 174454
rect 303722 174218 303764 174454
rect 303444 174134 303764 174218
rect 303444 173898 303486 174134
rect 303722 173898 303764 174134
rect 303444 173866 303764 173898
rect 311286 174454 311606 174486
rect 311286 174218 311328 174454
rect 311564 174218 311606 174454
rect 311286 174134 311606 174218
rect 311286 173898 311328 174134
rect 311564 173898 311606 174134
rect 311286 173866 311606 173898
rect 319128 174454 319448 174486
rect 319128 174218 319170 174454
rect 319406 174218 319448 174454
rect 319128 174134 319448 174218
rect 319128 173898 319170 174134
rect 319406 173898 319448 174134
rect 319128 173866 319448 173898
rect 326970 174454 327290 174486
rect 326970 174218 327012 174454
rect 327248 174218 327290 174454
rect 326970 174134 327290 174218
rect 326970 173898 327012 174134
rect 327248 173898 327290 174134
rect 326970 173866 327290 173898
rect 307365 168174 307685 168206
rect 307365 167938 307407 168174
rect 307643 167938 307685 168174
rect 307365 167854 307685 167938
rect 307365 167618 307407 167854
rect 307643 167618 307685 167854
rect 307365 167586 307685 167618
rect 315207 168174 315527 168206
rect 315207 167938 315249 168174
rect 315485 167938 315527 168174
rect 315207 167854 315527 167938
rect 315207 167618 315249 167854
rect 315485 167618 315527 167854
rect 315207 167586 315527 167618
rect 323049 168174 323369 168206
rect 323049 167938 323091 168174
rect 323327 167938 323369 168174
rect 323049 167854 323369 167938
rect 323049 167618 323091 167854
rect 323327 167618 323369 167854
rect 323049 167586 323369 167618
rect 330891 168174 331211 168206
rect 330891 167938 330933 168174
rect 331169 167938 331211 168174
rect 330891 167854 331211 167938
rect 330891 167618 330933 167854
rect 331169 167618 331211 167854
rect 330891 167586 331211 167618
rect 303444 164454 303764 164486
rect 303444 164218 303486 164454
rect 303722 164218 303764 164454
rect 303444 164134 303764 164218
rect 303444 163898 303486 164134
rect 303722 163898 303764 164134
rect 303444 163866 303764 163898
rect 311286 164454 311606 164486
rect 311286 164218 311328 164454
rect 311564 164218 311606 164454
rect 311286 164134 311606 164218
rect 311286 163898 311328 164134
rect 311564 163898 311606 164134
rect 311286 163866 311606 163898
rect 319128 164454 319448 164486
rect 319128 164218 319170 164454
rect 319406 164218 319448 164454
rect 319128 164134 319448 164218
rect 319128 163898 319170 164134
rect 319406 163898 319448 164134
rect 319128 163866 319448 163898
rect 326970 164454 327290 164486
rect 326970 164218 327012 164454
rect 327248 164218 327290 164454
rect 326970 164134 327290 164218
rect 326970 163898 327012 164134
rect 327248 163898 327290 164134
rect 326970 163866 327290 163898
rect 307707 158132 307773 158133
rect 307707 158068 307708 158132
rect 307772 158068 307773 158132
rect 307707 158067 307773 158068
rect 303659 157452 303725 157453
rect 303659 157388 303660 157452
rect 303724 157388 303725 157452
rect 303659 157387 303725 157388
rect 303110 74490 303538 74550
rect 302555 68372 302621 68373
rect 302555 68308 302556 68372
rect 302620 68308 302621 68372
rect 302555 68307 302621 68308
rect 302220 65590 302434 65650
rect 302558 65620 302618 68307
rect 303478 65620 303538 74490
rect 303662 68237 303722 157387
rect 306419 157180 306485 157181
rect 306419 157116 306420 157180
rect 306484 157116 306485 157180
rect 306419 157115 306485 157116
rect 305683 156908 305749 156909
rect 305683 156844 305684 156908
rect 305748 156844 305749 156908
rect 305683 156843 305749 156844
rect 303843 156636 303909 156637
rect 303843 156572 303844 156636
rect 303908 156572 303909 156636
rect 303843 156571 303909 156572
rect 303846 68781 303906 156571
rect 304211 68916 304277 68917
rect 304211 68852 304212 68916
rect 304276 68852 304277 68916
rect 304211 68851 304277 68852
rect 305315 68916 305381 68917
rect 305315 68852 305316 68916
rect 305380 68852 305381 68916
rect 305315 68851 305381 68852
rect 303843 68780 303909 68781
rect 303843 68716 303844 68780
rect 303908 68716 303909 68780
rect 303843 68715 303909 68716
rect 303659 68236 303725 68237
rect 303659 68172 303660 68236
rect 303724 68172 303725 68236
rect 303659 68171 303725 68172
rect 303843 67148 303909 67149
rect 303843 67084 303844 67148
rect 303908 67084 303909 67148
rect 303843 67083 303909 67084
rect 303846 65620 303906 67083
rect 304214 65620 304274 68851
rect 304579 68508 304645 68509
rect 304579 68444 304580 68508
rect 304644 68444 304645 68508
rect 304579 68443 304645 68444
rect 304582 65620 304642 68443
rect 304947 66876 305013 66877
rect 304947 66812 304948 66876
rect 305012 66812 305013 66876
rect 304947 66811 305013 66812
rect 304950 65620 305010 66811
rect 305318 65620 305378 68851
rect 305686 65620 305746 156843
rect 306422 74629 306482 157115
rect 307710 74765 307770 158067
rect 311939 156772 312005 156773
rect 311939 156708 311940 156772
rect 312004 156708 312005 156772
rect 311939 156707 312005 156708
rect 307891 156636 307957 156637
rect 307891 156572 307892 156636
rect 307956 156572 307957 156636
rect 307891 156571 307957 156572
rect 307707 74764 307773 74765
rect 307707 74700 307708 74764
rect 307772 74700 307773 74764
rect 307707 74699 307773 74700
rect 306419 74628 306485 74629
rect 306419 74564 306420 74628
rect 306484 74564 306485 74628
rect 306419 74563 306485 74564
rect 307155 73812 307221 73813
rect 307155 73748 307156 73812
rect 307220 73748 307221 73812
rect 307155 73747 307221 73748
rect 306235 69596 306301 69597
rect 306235 69532 306236 69596
rect 306300 69532 306301 69596
rect 306235 69531 306301 69532
rect 306238 67650 306298 69531
rect 306787 68236 306853 68237
rect 306787 68172 306788 68236
rect 306852 68172 306853 68236
rect 306787 68171 306853 68172
rect 306238 67590 306482 67650
rect 306051 67556 306117 67557
rect 306051 67492 306052 67556
rect 306116 67492 306117 67556
rect 306051 67491 306117 67492
rect 306054 65620 306114 67491
rect 306422 65620 306482 67590
rect 306790 65620 306850 68171
rect 307158 65620 307218 73747
rect 307523 72452 307589 72453
rect 307523 72388 307524 72452
rect 307588 72388 307589 72452
rect 307523 72387 307589 72388
rect 307526 65620 307586 72387
rect 307894 65620 307954 156571
rect 311019 155276 311085 155277
rect 311019 155212 311020 155276
rect 311084 155212 311085 155276
rect 311019 155211 311085 155212
rect 309363 153780 309429 153781
rect 309363 153716 309364 153780
rect 309428 153716 309429 153780
rect 309363 153715 309429 153716
rect 308995 75172 309061 75173
rect 308995 75108 308996 75172
rect 309060 75108 309061 75172
rect 308995 75107 309061 75108
rect 308259 71092 308325 71093
rect 308259 71028 308260 71092
rect 308324 71028 308325 71092
rect 308259 71027 308325 71028
rect 308262 65620 308322 71027
rect 308627 69596 308693 69597
rect 308627 69532 308628 69596
rect 308692 69532 308693 69596
rect 308627 69531 308693 69532
rect 308630 65620 308690 69531
rect 308998 65620 309058 75107
rect 309366 65620 309426 153715
rect 292992 64171 293312 64240
rect 292992 63935 293034 64171
rect 293270 63935 293312 64171
rect 292992 63866 293312 63935
rect 277632 58174 277952 58206
rect 277632 57938 277674 58174
rect 277910 57938 277952 58174
rect 277632 57854 277952 57938
rect 277632 57618 277674 57854
rect 277910 57618 277952 57854
rect 277632 57586 277952 57618
rect 308352 58174 308672 58206
rect 308352 57938 308394 58174
rect 308630 57938 308672 58174
rect 308352 57854 308672 57938
rect 308352 57618 308394 57854
rect 308630 57618 308672 57854
rect 308352 57586 308672 57618
rect 292992 54454 293312 54486
rect 292992 54218 293034 54454
rect 293270 54218 293312 54454
rect 292992 54134 293312 54218
rect 292992 53898 293034 54134
rect 293270 53898 293312 54134
rect 292992 53866 293312 53898
rect 277632 48174 277952 48206
rect 277632 47938 277674 48174
rect 277910 47938 277952 48174
rect 277632 47854 277952 47938
rect 277632 47618 277674 47854
rect 277910 47618 277952 47854
rect 277632 47586 277952 47618
rect 308352 48174 308672 48206
rect 308352 47938 308394 48174
rect 308630 47938 308672 48174
rect 308352 47854 308672 47938
rect 308352 47618 308394 47854
rect 308630 47618 308672 47854
rect 308352 47586 308672 47618
rect 292992 44454 293312 44486
rect 292992 44218 293034 44454
rect 293270 44218 293312 44454
rect 292992 44134 293312 44218
rect 292992 43898 293034 44134
rect 293270 43898 293312 44134
rect 292992 43866 293312 43898
rect 277632 38174 277952 38206
rect 277632 37938 277674 38174
rect 277910 37938 277952 38174
rect 277632 37854 277952 37938
rect 277632 37618 277674 37854
rect 277910 37618 277952 37854
rect 277632 37586 277952 37618
rect 308352 38174 308672 38206
rect 308352 37938 308394 38174
rect 308630 37938 308672 38174
rect 308352 37854 308672 37938
rect 308352 37618 308394 37854
rect 308630 37618 308672 37854
rect 308352 37586 308672 37618
rect 292992 34454 293312 34486
rect 292992 34218 293034 34454
rect 293270 34218 293312 34454
rect 292992 34134 293312 34218
rect 292992 33898 293034 34134
rect 293270 33898 293312 34134
rect 292992 33866 293312 33898
rect 273299 22676 273365 22677
rect 273299 22612 273300 22676
rect 273364 22612 273365 22676
rect 273299 22611 273365 22612
rect 273302 20637 273362 22611
rect 275510 22070 275724 22130
rect 276092 22070 276306 22130
rect 275510 21861 275570 22070
rect 276246 21997 276306 22070
rect 276614 22070 276828 22130
rect 276243 21996 276309 21997
rect 276243 21932 276244 21996
rect 276308 21932 276309 21996
rect 276243 21931 276309 21932
rect 275507 21860 275573 21861
rect 275507 21796 275508 21860
rect 275572 21796 275573 21860
rect 275507 21795 275573 21796
rect 273299 20636 273365 20637
rect 273299 20572 273300 20636
rect 273364 20572 273365 20636
rect 273299 20571 273365 20572
rect 275326 20093 275386 21760
rect 275323 20092 275389 20093
rect 275323 20028 275324 20092
rect 275388 20028 275389 20092
rect 275323 20027 275389 20028
rect 276430 19277 276490 21760
rect 276614 21725 276674 22070
rect 276611 21724 276677 21725
rect 276611 21660 276612 21724
rect 276676 21660 276677 21724
rect 276611 21659 276677 21660
rect 277166 20365 277226 22100
rect 306268 22070 306482 22130
rect 306422 21997 306482 22070
rect 306419 21996 306485 21997
rect 306419 21932 306420 21996
rect 306484 21932 306485 21996
rect 306419 21931 306485 21932
rect 277163 20364 277229 20365
rect 277163 20300 277164 20364
rect 277228 20300 277229 20364
rect 277163 20299 277229 20300
rect 277534 20229 277594 21760
rect 277902 20501 277962 21760
rect 278270 20637 278330 21760
rect 278267 20636 278333 20637
rect 278267 20572 278268 20636
rect 278332 20572 278333 20636
rect 278267 20571 278333 20572
rect 277899 20500 277965 20501
rect 277899 20436 277900 20500
rect 277964 20436 277965 20500
rect 277899 20435 277965 20436
rect 277531 20228 277597 20229
rect 277531 20164 277532 20228
rect 277596 20164 277597 20228
rect 277531 20163 277597 20164
rect 276427 19276 276493 19277
rect 276427 19212 276428 19276
rect 276492 19212 276493 19276
rect 276427 19211 276493 19212
rect 278638 19141 278698 21760
rect 279006 19277 279066 21760
rect 306606 20637 306666 21760
rect 311022 20637 311082 155211
rect 311942 68645 312002 156707
rect 311939 68644 312005 68645
rect 311939 68580 311940 68644
rect 312004 68580 312005 68644
rect 311939 68579 312005 68580
rect 334758 68373 334818 178739
rect 339174 178500 339234 179860
rect 339910 178500 339970 179520
rect 340646 178876 340706 179520
rect 341382 178876 341442 179520
rect 342118 178876 342178 179520
rect 342854 178876 342914 179520
rect 343590 178876 343650 179520
rect 344326 178876 344386 179520
rect 345062 178876 345122 179520
rect 345798 178840 345858 179520
rect 346534 178840 346594 179520
rect 347270 178840 347330 179520
rect 348006 178840 348066 179520
rect 348742 178840 348802 179860
rect 349478 178840 349538 179520
rect 350214 178840 350274 179860
rect 350950 178840 351010 179520
rect 351686 178840 351746 179860
rect 352422 178500 352482 179520
rect 353158 178840 353218 179520
rect 353894 178500 353954 179520
rect 354630 178500 354690 179520
rect 355366 178840 355426 179520
rect 356102 178840 356162 179520
rect 356838 178500 356898 179520
rect 357574 178840 357634 179520
rect 358310 178500 358370 179520
rect 359046 178840 359106 179520
rect 359782 178500 359842 179520
rect 360518 178500 360578 179520
rect 361254 178840 361314 179520
rect 361990 178840 362050 179520
rect 362726 178840 362786 179520
rect 363462 178840 363522 179520
rect 364198 178840 364258 179520
rect 364934 178840 364994 179520
rect 365670 178840 365730 179520
rect 366406 178500 366466 179520
rect 367142 178840 367202 179520
rect 367878 178840 367938 179520
rect 368614 178500 368674 179520
rect 371834 178876 371894 179520
rect 372570 178840 372630 179520
rect 373306 178500 373366 179520
rect 374042 178500 374102 179520
rect 374778 178876 374838 179520
rect 375514 178876 375574 179520
rect 376250 178876 376310 179520
rect 376986 178876 377046 179520
rect 377722 178876 377782 179520
rect 378458 178876 378518 179520
rect 379194 178876 379254 179520
rect 379930 178840 379990 179520
rect 380666 178840 380726 179520
rect 381402 178840 381462 179520
rect 382138 178840 382198 179520
rect 382874 178840 382934 179520
rect 383610 178840 383670 179520
rect 384346 178840 384406 179520
rect 385082 178840 385142 179520
rect 385818 178840 385878 179520
rect 386554 178500 386614 179520
rect 387290 178840 387350 179520
rect 388026 178500 388086 179520
rect 388762 178500 388822 179520
rect 389498 178840 389558 179520
rect 390234 178840 390294 179520
rect 390970 178500 391030 179520
rect 391706 178840 391766 179520
rect 392442 178500 392502 179520
rect 393178 178840 393238 179520
rect 393914 178500 393974 179520
rect 394650 178500 394710 179520
rect 395386 178840 395446 179520
rect 396122 178840 396182 179520
rect 396858 178840 396918 179520
rect 397594 178840 397654 179520
rect 398330 178840 398390 179520
rect 399066 178840 399126 179520
rect 399802 178840 399862 179520
rect 400538 178500 400598 179520
rect 401274 178840 401334 179520
rect 402010 178840 402070 179520
rect 402746 178500 402806 179520
rect 405966 178876 406026 179520
rect 406702 178840 406762 179520
rect 407438 178500 407498 179520
rect 408174 178500 408234 179520
rect 408910 178876 408970 179520
rect 409646 178876 409706 179520
rect 410382 178876 410442 179520
rect 411118 178876 411178 179520
rect 411854 178876 411914 179520
rect 412590 178876 412650 179520
rect 413326 178876 413386 179520
rect 414062 178840 414122 179520
rect 414798 178840 414858 179520
rect 415534 178840 415594 179860
rect 416270 178840 416330 179520
rect 417006 178840 417066 179520
rect 417742 178840 417802 179860
rect 418478 178840 418538 179520
rect 419214 178840 419274 179520
rect 419950 178840 420010 179520
rect 420686 178500 420746 179520
rect 421422 178840 421482 179520
rect 422158 178500 422218 179520
rect 422894 178500 422954 179520
rect 423630 178840 423690 179520
rect 424366 178840 424426 179520
rect 425102 178500 425162 179520
rect 425838 178840 425898 179520
rect 426574 178500 426634 179520
rect 427310 178840 427370 179520
rect 428046 178500 428106 179520
rect 428782 178500 428842 179520
rect 429518 178840 429578 179520
rect 430254 178840 430314 179520
rect 430990 178840 431050 179520
rect 431726 178840 431786 179520
rect 432462 178840 432522 179520
rect 433198 178840 433258 179520
rect 433934 178840 433994 179520
rect 434670 178500 434730 179520
rect 435406 178840 435466 179520
rect 436142 178840 436202 179520
rect 436878 178500 436938 179520
rect 440098 178876 440158 179520
rect 440834 178840 440894 179520
rect 441570 178500 441630 179520
rect 442306 178500 442366 179520
rect 443042 178876 443102 179520
rect 443778 178876 443838 179520
rect 444514 178876 444574 179520
rect 445250 178876 445310 179520
rect 445986 178876 446046 179520
rect 446722 178876 446782 179520
rect 447458 178876 447518 179520
rect 448194 178840 448254 179520
rect 448930 178840 448990 179520
rect 449666 178840 449726 179520
rect 450402 178840 450462 179520
rect 451138 178840 451198 179520
rect 451874 178840 451934 179520
rect 452610 178840 452670 179520
rect 453346 178840 453406 179520
rect 454082 178840 454142 179520
rect 454818 178500 454878 179520
rect 455554 178840 455614 179520
rect 456290 178500 456350 179520
rect 457026 178500 457086 179520
rect 457762 178840 457822 179520
rect 458498 178840 458558 179520
rect 459234 178500 459294 179520
rect 459970 178840 460030 179520
rect 460706 178500 460766 179520
rect 461442 178840 461502 179520
rect 462178 178500 462238 179520
rect 462914 178500 462974 179520
rect 463650 178840 463710 179520
rect 464386 178840 464446 179520
rect 465122 178840 465182 179520
rect 465858 178840 465918 179520
rect 466594 178840 466654 179520
rect 467330 178840 467390 179520
rect 468066 178840 468126 179520
rect 468802 178500 468862 179520
rect 469538 178840 469598 179520
rect 470274 178840 470334 179520
rect 471010 178500 471070 179520
rect 474230 178876 474290 179520
rect 474966 178840 475026 179520
rect 475702 178500 475762 179520
rect 476438 178500 476498 179520
rect 477174 178876 477234 179520
rect 477910 178876 477970 179520
rect 478646 178876 478706 179520
rect 479382 178876 479442 179520
rect 480118 178876 480178 179520
rect 480854 178876 480914 179520
rect 481590 178876 481650 179520
rect 482326 178840 482386 179520
rect 483062 178840 483122 179520
rect 483798 178840 483858 179520
rect 484534 178840 484594 179520
rect 485270 178840 485330 179520
rect 486006 178840 486066 179520
rect 486742 178840 486802 179520
rect 487478 178840 487538 179520
rect 488214 178840 488274 179520
rect 488950 178500 489010 179520
rect 489686 178840 489746 179520
rect 490422 178500 490482 179520
rect 491158 178500 491218 179520
rect 491894 178840 491954 179520
rect 492630 178840 492690 179520
rect 493366 178500 493426 179520
rect 494102 178840 494162 179520
rect 494838 178500 494898 179520
rect 495574 178840 495634 179520
rect 496310 178500 496370 179520
rect 497046 178500 497106 179520
rect 497782 178840 497842 179520
rect 498518 178840 498578 179520
rect 499254 178840 499314 179520
rect 499990 178840 500050 179520
rect 500726 178840 500786 179520
rect 501462 178840 501522 179520
rect 502198 178840 502258 179520
rect 502934 178500 502994 179520
rect 503670 178840 503730 179520
rect 504406 178840 504466 179520
rect 505142 178500 505202 179520
rect 508362 178876 508422 179520
rect 509098 178840 509158 179520
rect 509834 178500 509894 179520
rect 510570 178500 510630 179520
rect 511306 178876 511366 179520
rect 512042 178876 512102 179520
rect 512778 178876 512838 179520
rect 513514 178876 513574 179520
rect 514250 178876 514310 179520
rect 514986 178876 515046 179520
rect 515722 178876 515782 179520
rect 516458 178840 516518 179520
rect 517194 178840 517254 179520
rect 517930 178840 517990 179520
rect 518666 178840 518726 179520
rect 519402 178840 519462 179520
rect 520138 178840 520198 179520
rect 520874 178840 520934 179520
rect 521610 178840 521670 179520
rect 522346 178840 522406 179520
rect 523082 178500 523142 179520
rect 523818 178840 523878 179520
rect 524554 178500 524614 179520
rect 525290 178500 525350 179520
rect 526026 178840 526086 179520
rect 526762 178840 526822 179520
rect 527498 178500 527558 179520
rect 528234 178840 528294 179520
rect 528970 178500 529030 179520
rect 529706 178840 529766 179520
rect 530442 178500 530502 179520
rect 531178 178500 531238 179520
rect 531914 178840 531974 179520
rect 532650 178840 532710 179520
rect 533386 178840 533446 179520
rect 534122 178840 534182 179520
rect 534858 178840 534918 179520
rect 535594 178840 535654 179520
rect 536330 178840 536390 179520
rect 537066 178500 537126 179520
rect 537802 178840 537862 179520
rect 538538 178840 538598 179520
rect 539274 178500 539334 179520
rect 542494 178876 542554 179520
rect 543230 178840 543290 179520
rect 543966 178500 544026 179520
rect 544702 178500 544762 179520
rect 545438 178876 545498 179520
rect 546174 178876 546234 179520
rect 546910 178876 546970 179520
rect 547646 178876 547706 179520
rect 548382 178876 548442 179520
rect 549118 178876 549178 179520
rect 549854 178876 549914 179860
rect 550590 178840 550650 179860
rect 551326 178840 551386 179520
rect 552062 178840 552122 179860
rect 552798 178840 552858 179860
rect 553534 178840 553594 179520
rect 554270 178840 554330 179520
rect 555006 178840 555066 179860
rect 555742 178840 555802 179860
rect 556478 178840 556538 179520
rect 557214 178500 557274 179520
rect 557950 178840 558010 179520
rect 558686 178500 558746 179520
rect 559422 178500 559482 179520
rect 560158 178840 560218 179520
rect 560894 178840 560954 179520
rect 561630 178500 561690 179520
rect 562366 178840 562426 179520
rect 563102 178500 563162 179520
rect 563838 178840 563898 179520
rect 564574 178500 564634 179520
rect 565310 178500 565370 179520
rect 566046 178840 566106 179520
rect 566782 178840 566842 179520
rect 567518 178840 567578 179520
rect 568254 178840 568314 179520
rect 568990 178840 569050 179520
rect 569726 178840 569786 179520
rect 570462 178840 570522 179520
rect 571198 178500 571258 179520
rect 571934 178840 571994 179520
rect 572670 178840 572730 179520
rect 573406 178500 573466 179520
rect 341497 177879 341817 177936
rect 341497 177643 341539 177879
rect 341775 177643 341817 177879
rect 341497 177586 341817 177643
rect 349339 177879 349659 177936
rect 349339 177643 349381 177879
rect 349617 177643 349659 177879
rect 349339 177586 349659 177643
rect 357181 177879 357501 177936
rect 357181 177643 357223 177879
rect 357459 177643 357501 177879
rect 357181 177586 357501 177643
rect 365023 177879 365343 177936
rect 365023 177643 365065 177879
rect 365301 177643 365343 177879
rect 365023 177586 365343 177643
rect 375629 177879 375949 177936
rect 375629 177643 375671 177879
rect 375907 177643 375949 177879
rect 375629 177586 375949 177643
rect 383471 177879 383791 177936
rect 383471 177643 383513 177879
rect 383749 177643 383791 177879
rect 383471 177586 383791 177643
rect 391313 177879 391633 177936
rect 391313 177643 391355 177879
rect 391591 177643 391633 177879
rect 391313 177586 391633 177643
rect 399155 177879 399475 177936
rect 399155 177643 399197 177879
rect 399433 177643 399475 177879
rect 399155 177586 399475 177643
rect 409761 177879 410081 177936
rect 409761 177643 409803 177879
rect 410039 177643 410081 177879
rect 409761 177586 410081 177643
rect 417603 177879 417923 177936
rect 417603 177643 417645 177879
rect 417881 177643 417923 177879
rect 417603 177586 417923 177643
rect 425445 177879 425765 177936
rect 425445 177643 425487 177879
rect 425723 177643 425765 177879
rect 425445 177586 425765 177643
rect 433287 177879 433607 177936
rect 433287 177643 433329 177879
rect 433565 177643 433607 177879
rect 433287 177586 433607 177643
rect 443893 177879 444213 177936
rect 443893 177643 443935 177879
rect 444171 177643 444213 177879
rect 443893 177586 444213 177643
rect 451735 177879 452055 177936
rect 451735 177643 451777 177879
rect 452013 177643 452055 177879
rect 451735 177586 452055 177643
rect 459577 177879 459897 177936
rect 459577 177643 459619 177879
rect 459855 177643 459897 177879
rect 459577 177586 459897 177643
rect 467419 177879 467739 177936
rect 467419 177643 467461 177879
rect 467697 177643 467739 177879
rect 467419 177586 467739 177643
rect 478025 177879 478345 177936
rect 478025 177643 478067 177879
rect 478303 177643 478345 177879
rect 478025 177586 478345 177643
rect 485867 177879 486187 177936
rect 485867 177643 485909 177879
rect 486145 177643 486187 177879
rect 485867 177586 486187 177643
rect 493709 177879 494029 177936
rect 493709 177643 493751 177879
rect 493987 177643 494029 177879
rect 493709 177586 494029 177643
rect 501551 177879 501871 177936
rect 501551 177643 501593 177879
rect 501829 177643 501871 177879
rect 501551 177586 501871 177643
rect 512157 177879 512477 177936
rect 512157 177643 512199 177879
rect 512435 177643 512477 177879
rect 512157 177586 512477 177643
rect 519999 177879 520319 177936
rect 519999 177643 520041 177879
rect 520277 177643 520319 177879
rect 519999 177586 520319 177643
rect 527841 177879 528161 177936
rect 527841 177643 527883 177879
rect 528119 177643 528161 177879
rect 527841 177586 528161 177643
rect 535683 177879 536003 177936
rect 535683 177643 535725 177879
rect 535961 177643 536003 177879
rect 535683 177586 536003 177643
rect 546289 177879 546609 177936
rect 546289 177643 546331 177879
rect 546567 177643 546609 177879
rect 546289 177586 546609 177643
rect 554131 177879 554451 177936
rect 554131 177643 554173 177879
rect 554409 177643 554451 177879
rect 554131 177586 554451 177643
rect 561973 177879 562293 177936
rect 561973 177643 562015 177879
rect 562251 177643 562293 177879
rect 561973 177586 562293 177643
rect 569815 177879 570135 177936
rect 569815 177643 569857 177879
rect 570093 177643 570135 177879
rect 569815 177586 570135 177643
rect 337576 174454 337896 174486
rect 337576 174218 337618 174454
rect 337854 174218 337896 174454
rect 337576 174134 337896 174218
rect 337576 173898 337618 174134
rect 337854 173898 337896 174134
rect 337576 173866 337896 173898
rect 345418 174454 345738 174486
rect 345418 174218 345460 174454
rect 345696 174218 345738 174454
rect 345418 174134 345738 174218
rect 345418 173898 345460 174134
rect 345696 173898 345738 174134
rect 345418 173866 345738 173898
rect 353260 174454 353580 174486
rect 353260 174218 353302 174454
rect 353538 174218 353580 174454
rect 353260 174134 353580 174218
rect 353260 173898 353302 174134
rect 353538 173898 353580 174134
rect 353260 173866 353580 173898
rect 361102 174454 361422 174486
rect 361102 174218 361144 174454
rect 361380 174218 361422 174454
rect 361102 174134 361422 174218
rect 361102 173898 361144 174134
rect 361380 173898 361422 174134
rect 361102 173866 361422 173898
rect 371708 174454 372028 174486
rect 371708 174218 371750 174454
rect 371986 174218 372028 174454
rect 371708 174134 372028 174218
rect 371708 173898 371750 174134
rect 371986 173898 372028 174134
rect 371708 173866 372028 173898
rect 379550 174454 379870 174486
rect 379550 174218 379592 174454
rect 379828 174218 379870 174454
rect 379550 174134 379870 174218
rect 379550 173898 379592 174134
rect 379828 173898 379870 174134
rect 379550 173866 379870 173898
rect 387392 174454 387712 174486
rect 387392 174218 387434 174454
rect 387670 174218 387712 174454
rect 387392 174134 387712 174218
rect 387392 173898 387434 174134
rect 387670 173898 387712 174134
rect 387392 173866 387712 173898
rect 395234 174454 395554 174486
rect 395234 174218 395276 174454
rect 395512 174218 395554 174454
rect 395234 174134 395554 174218
rect 395234 173898 395276 174134
rect 395512 173898 395554 174134
rect 395234 173866 395554 173898
rect 405840 174454 406160 174486
rect 405840 174218 405882 174454
rect 406118 174218 406160 174454
rect 405840 174134 406160 174218
rect 405840 173898 405882 174134
rect 406118 173898 406160 174134
rect 405840 173866 406160 173898
rect 413682 174454 414002 174486
rect 413682 174218 413724 174454
rect 413960 174218 414002 174454
rect 413682 174134 414002 174218
rect 413682 173898 413724 174134
rect 413960 173898 414002 174134
rect 413682 173866 414002 173898
rect 421524 174454 421844 174486
rect 421524 174218 421566 174454
rect 421802 174218 421844 174454
rect 421524 174134 421844 174218
rect 421524 173898 421566 174134
rect 421802 173898 421844 174134
rect 421524 173866 421844 173898
rect 429366 174454 429686 174486
rect 429366 174218 429408 174454
rect 429644 174218 429686 174454
rect 429366 174134 429686 174218
rect 429366 173898 429408 174134
rect 429644 173898 429686 174134
rect 429366 173866 429686 173898
rect 439972 174454 440292 174486
rect 439972 174218 440014 174454
rect 440250 174218 440292 174454
rect 439972 174134 440292 174218
rect 439972 173898 440014 174134
rect 440250 173898 440292 174134
rect 439972 173866 440292 173898
rect 447814 174454 448134 174486
rect 447814 174218 447856 174454
rect 448092 174218 448134 174454
rect 447814 174134 448134 174218
rect 447814 173898 447856 174134
rect 448092 173898 448134 174134
rect 447814 173866 448134 173898
rect 455656 174454 455976 174486
rect 455656 174218 455698 174454
rect 455934 174218 455976 174454
rect 455656 174134 455976 174218
rect 455656 173898 455698 174134
rect 455934 173898 455976 174134
rect 455656 173866 455976 173898
rect 463498 174454 463818 174486
rect 463498 174218 463540 174454
rect 463776 174218 463818 174454
rect 463498 174134 463818 174218
rect 463498 173898 463540 174134
rect 463776 173898 463818 174134
rect 463498 173866 463818 173898
rect 474104 174454 474424 174486
rect 474104 174218 474146 174454
rect 474382 174218 474424 174454
rect 474104 174134 474424 174218
rect 474104 173898 474146 174134
rect 474382 173898 474424 174134
rect 474104 173866 474424 173898
rect 481946 174454 482266 174486
rect 481946 174218 481988 174454
rect 482224 174218 482266 174454
rect 481946 174134 482266 174218
rect 481946 173898 481988 174134
rect 482224 173898 482266 174134
rect 481946 173866 482266 173898
rect 489788 174454 490108 174486
rect 489788 174218 489830 174454
rect 490066 174218 490108 174454
rect 489788 174134 490108 174218
rect 489788 173898 489830 174134
rect 490066 173898 490108 174134
rect 489788 173866 490108 173898
rect 497630 174454 497950 174486
rect 497630 174218 497672 174454
rect 497908 174218 497950 174454
rect 497630 174134 497950 174218
rect 497630 173898 497672 174134
rect 497908 173898 497950 174134
rect 497630 173866 497950 173898
rect 508236 174454 508556 174486
rect 508236 174218 508278 174454
rect 508514 174218 508556 174454
rect 508236 174134 508556 174218
rect 508236 173898 508278 174134
rect 508514 173898 508556 174134
rect 508236 173866 508556 173898
rect 516078 174454 516398 174486
rect 516078 174218 516120 174454
rect 516356 174218 516398 174454
rect 516078 174134 516398 174218
rect 516078 173898 516120 174134
rect 516356 173898 516398 174134
rect 516078 173866 516398 173898
rect 523920 174454 524240 174486
rect 523920 174218 523962 174454
rect 524198 174218 524240 174454
rect 523920 174134 524240 174218
rect 523920 173898 523962 174134
rect 524198 173898 524240 174134
rect 523920 173866 524240 173898
rect 531762 174454 532082 174486
rect 531762 174218 531804 174454
rect 532040 174218 532082 174454
rect 531762 174134 532082 174218
rect 531762 173898 531804 174134
rect 532040 173898 532082 174134
rect 531762 173866 532082 173898
rect 542368 174454 542688 174486
rect 542368 174218 542410 174454
rect 542646 174218 542688 174454
rect 542368 174134 542688 174218
rect 542368 173898 542410 174134
rect 542646 173898 542688 174134
rect 542368 173866 542688 173898
rect 550210 174454 550530 174486
rect 550210 174218 550252 174454
rect 550488 174218 550530 174454
rect 550210 174134 550530 174218
rect 550210 173898 550252 174134
rect 550488 173898 550530 174134
rect 550210 173866 550530 173898
rect 558052 174454 558372 174486
rect 558052 174218 558094 174454
rect 558330 174218 558372 174454
rect 558052 174134 558372 174218
rect 558052 173898 558094 174134
rect 558330 173898 558372 174134
rect 558052 173866 558372 173898
rect 565894 174454 566214 174486
rect 565894 174218 565936 174454
rect 566172 174218 566214 174454
rect 565894 174134 566214 174218
rect 565894 173898 565936 174134
rect 566172 173898 566214 174134
rect 565894 173866 566214 173898
rect 341497 168174 341817 168206
rect 341497 167938 341539 168174
rect 341775 167938 341817 168174
rect 341497 167854 341817 167938
rect 341497 167618 341539 167854
rect 341775 167618 341817 167854
rect 341497 167586 341817 167618
rect 349339 168174 349659 168206
rect 349339 167938 349381 168174
rect 349617 167938 349659 168174
rect 349339 167854 349659 167938
rect 349339 167618 349381 167854
rect 349617 167618 349659 167854
rect 349339 167586 349659 167618
rect 357181 168174 357501 168206
rect 357181 167938 357223 168174
rect 357459 167938 357501 168174
rect 357181 167854 357501 167938
rect 357181 167618 357223 167854
rect 357459 167618 357501 167854
rect 357181 167586 357501 167618
rect 365023 168174 365343 168206
rect 365023 167938 365065 168174
rect 365301 167938 365343 168174
rect 365023 167854 365343 167938
rect 365023 167618 365065 167854
rect 365301 167618 365343 167854
rect 365023 167586 365343 167618
rect 375629 168174 375949 168206
rect 375629 167938 375671 168174
rect 375907 167938 375949 168174
rect 375629 167854 375949 167938
rect 375629 167618 375671 167854
rect 375907 167618 375949 167854
rect 375629 167586 375949 167618
rect 383471 168174 383791 168206
rect 383471 167938 383513 168174
rect 383749 167938 383791 168174
rect 383471 167854 383791 167938
rect 383471 167618 383513 167854
rect 383749 167618 383791 167854
rect 383471 167586 383791 167618
rect 391313 168174 391633 168206
rect 391313 167938 391355 168174
rect 391591 167938 391633 168174
rect 391313 167854 391633 167938
rect 391313 167618 391355 167854
rect 391591 167618 391633 167854
rect 391313 167586 391633 167618
rect 399155 168174 399475 168206
rect 399155 167938 399197 168174
rect 399433 167938 399475 168174
rect 399155 167854 399475 167938
rect 399155 167618 399197 167854
rect 399433 167618 399475 167854
rect 399155 167586 399475 167618
rect 409761 168174 410081 168206
rect 409761 167938 409803 168174
rect 410039 167938 410081 168174
rect 409761 167854 410081 167938
rect 409761 167618 409803 167854
rect 410039 167618 410081 167854
rect 409761 167586 410081 167618
rect 417603 168174 417923 168206
rect 417603 167938 417645 168174
rect 417881 167938 417923 168174
rect 417603 167854 417923 167938
rect 417603 167618 417645 167854
rect 417881 167618 417923 167854
rect 417603 167586 417923 167618
rect 425445 168174 425765 168206
rect 425445 167938 425487 168174
rect 425723 167938 425765 168174
rect 425445 167854 425765 167938
rect 425445 167618 425487 167854
rect 425723 167618 425765 167854
rect 425445 167586 425765 167618
rect 433287 168174 433607 168206
rect 433287 167938 433329 168174
rect 433565 167938 433607 168174
rect 433287 167854 433607 167938
rect 433287 167618 433329 167854
rect 433565 167618 433607 167854
rect 433287 167586 433607 167618
rect 443893 168174 444213 168206
rect 443893 167938 443935 168174
rect 444171 167938 444213 168174
rect 443893 167854 444213 167938
rect 443893 167618 443935 167854
rect 444171 167618 444213 167854
rect 443893 167586 444213 167618
rect 451735 168174 452055 168206
rect 451735 167938 451777 168174
rect 452013 167938 452055 168174
rect 451735 167854 452055 167938
rect 451735 167618 451777 167854
rect 452013 167618 452055 167854
rect 451735 167586 452055 167618
rect 459577 168174 459897 168206
rect 459577 167938 459619 168174
rect 459855 167938 459897 168174
rect 459577 167854 459897 167938
rect 459577 167618 459619 167854
rect 459855 167618 459897 167854
rect 459577 167586 459897 167618
rect 467419 168174 467739 168206
rect 467419 167938 467461 168174
rect 467697 167938 467739 168174
rect 467419 167854 467739 167938
rect 467419 167618 467461 167854
rect 467697 167618 467739 167854
rect 467419 167586 467739 167618
rect 478025 168174 478345 168206
rect 478025 167938 478067 168174
rect 478303 167938 478345 168174
rect 478025 167854 478345 167938
rect 478025 167618 478067 167854
rect 478303 167618 478345 167854
rect 478025 167586 478345 167618
rect 485867 168174 486187 168206
rect 485867 167938 485909 168174
rect 486145 167938 486187 168174
rect 485867 167854 486187 167938
rect 485867 167618 485909 167854
rect 486145 167618 486187 167854
rect 485867 167586 486187 167618
rect 493709 168174 494029 168206
rect 493709 167938 493751 168174
rect 493987 167938 494029 168174
rect 493709 167854 494029 167938
rect 493709 167618 493751 167854
rect 493987 167618 494029 167854
rect 493709 167586 494029 167618
rect 501551 168174 501871 168206
rect 501551 167938 501593 168174
rect 501829 167938 501871 168174
rect 501551 167854 501871 167938
rect 501551 167618 501593 167854
rect 501829 167618 501871 167854
rect 501551 167586 501871 167618
rect 512157 168174 512477 168206
rect 512157 167938 512199 168174
rect 512435 167938 512477 168174
rect 512157 167854 512477 167938
rect 512157 167618 512199 167854
rect 512435 167618 512477 167854
rect 512157 167586 512477 167618
rect 519999 168174 520319 168206
rect 519999 167938 520041 168174
rect 520277 167938 520319 168174
rect 519999 167854 520319 167938
rect 519999 167618 520041 167854
rect 520277 167618 520319 167854
rect 519999 167586 520319 167618
rect 527841 168174 528161 168206
rect 527841 167938 527883 168174
rect 528119 167938 528161 168174
rect 527841 167854 528161 167938
rect 527841 167618 527883 167854
rect 528119 167618 528161 167854
rect 527841 167586 528161 167618
rect 535683 168174 536003 168206
rect 535683 167938 535725 168174
rect 535961 167938 536003 168174
rect 535683 167854 536003 167938
rect 535683 167618 535725 167854
rect 535961 167618 536003 167854
rect 535683 167586 536003 167618
rect 546289 168174 546609 168206
rect 546289 167938 546331 168174
rect 546567 167938 546609 168174
rect 546289 167854 546609 167938
rect 546289 167618 546331 167854
rect 546567 167618 546609 167854
rect 546289 167586 546609 167618
rect 554131 168174 554451 168206
rect 554131 167938 554173 168174
rect 554409 167938 554451 168174
rect 554131 167854 554451 167938
rect 554131 167618 554173 167854
rect 554409 167618 554451 167854
rect 554131 167586 554451 167618
rect 561973 168174 562293 168206
rect 561973 167938 562015 168174
rect 562251 167938 562293 168174
rect 561973 167854 562293 167938
rect 561973 167618 562015 167854
rect 562251 167618 562293 167854
rect 561973 167586 562293 167618
rect 569815 168174 570135 168206
rect 569815 167938 569857 168174
rect 570093 167938 570135 168174
rect 569815 167854 570135 167938
rect 569815 167618 569857 167854
rect 570093 167618 570135 167854
rect 569815 167586 570135 167618
rect 337576 164454 337896 164486
rect 337576 164218 337618 164454
rect 337854 164218 337896 164454
rect 337576 164134 337896 164218
rect 337576 163898 337618 164134
rect 337854 163898 337896 164134
rect 337576 163866 337896 163898
rect 345418 164454 345738 164486
rect 345418 164218 345460 164454
rect 345696 164218 345738 164454
rect 345418 164134 345738 164218
rect 345418 163898 345460 164134
rect 345696 163898 345738 164134
rect 345418 163866 345738 163898
rect 353260 164454 353580 164486
rect 353260 164218 353302 164454
rect 353538 164218 353580 164454
rect 353260 164134 353580 164218
rect 353260 163898 353302 164134
rect 353538 163898 353580 164134
rect 353260 163866 353580 163898
rect 361102 164454 361422 164486
rect 361102 164218 361144 164454
rect 361380 164218 361422 164454
rect 361102 164134 361422 164218
rect 361102 163898 361144 164134
rect 361380 163898 361422 164134
rect 361102 163866 361422 163898
rect 371708 164454 372028 164486
rect 371708 164218 371750 164454
rect 371986 164218 372028 164454
rect 371708 164134 372028 164218
rect 371708 163898 371750 164134
rect 371986 163898 372028 164134
rect 371708 163866 372028 163898
rect 379550 164454 379870 164486
rect 379550 164218 379592 164454
rect 379828 164218 379870 164454
rect 379550 164134 379870 164218
rect 379550 163898 379592 164134
rect 379828 163898 379870 164134
rect 379550 163866 379870 163898
rect 387392 164454 387712 164486
rect 387392 164218 387434 164454
rect 387670 164218 387712 164454
rect 387392 164134 387712 164218
rect 387392 163898 387434 164134
rect 387670 163898 387712 164134
rect 387392 163866 387712 163898
rect 395234 164454 395554 164486
rect 395234 164218 395276 164454
rect 395512 164218 395554 164454
rect 395234 164134 395554 164218
rect 395234 163898 395276 164134
rect 395512 163898 395554 164134
rect 395234 163866 395554 163898
rect 405840 164454 406160 164486
rect 405840 164218 405882 164454
rect 406118 164218 406160 164454
rect 405840 164134 406160 164218
rect 405840 163898 405882 164134
rect 406118 163898 406160 164134
rect 405840 163866 406160 163898
rect 413682 164454 414002 164486
rect 413682 164218 413724 164454
rect 413960 164218 414002 164454
rect 413682 164134 414002 164218
rect 413682 163898 413724 164134
rect 413960 163898 414002 164134
rect 413682 163866 414002 163898
rect 421524 164454 421844 164486
rect 421524 164218 421566 164454
rect 421802 164218 421844 164454
rect 421524 164134 421844 164218
rect 421524 163898 421566 164134
rect 421802 163898 421844 164134
rect 421524 163866 421844 163898
rect 429366 164454 429686 164486
rect 429366 164218 429408 164454
rect 429644 164218 429686 164454
rect 429366 164134 429686 164218
rect 429366 163898 429408 164134
rect 429644 163898 429686 164134
rect 429366 163866 429686 163898
rect 439972 164454 440292 164486
rect 439972 164218 440014 164454
rect 440250 164218 440292 164454
rect 439972 164134 440292 164218
rect 439972 163898 440014 164134
rect 440250 163898 440292 164134
rect 439972 163866 440292 163898
rect 447814 164454 448134 164486
rect 447814 164218 447856 164454
rect 448092 164218 448134 164454
rect 447814 164134 448134 164218
rect 447814 163898 447856 164134
rect 448092 163898 448134 164134
rect 447814 163866 448134 163898
rect 455656 164454 455976 164486
rect 455656 164218 455698 164454
rect 455934 164218 455976 164454
rect 455656 164134 455976 164218
rect 455656 163898 455698 164134
rect 455934 163898 455976 164134
rect 455656 163866 455976 163898
rect 463498 164454 463818 164486
rect 463498 164218 463540 164454
rect 463776 164218 463818 164454
rect 463498 164134 463818 164218
rect 463498 163898 463540 164134
rect 463776 163898 463818 164134
rect 463498 163866 463818 163898
rect 474104 164454 474424 164486
rect 474104 164218 474146 164454
rect 474382 164218 474424 164454
rect 474104 164134 474424 164218
rect 474104 163898 474146 164134
rect 474382 163898 474424 164134
rect 474104 163866 474424 163898
rect 481946 164454 482266 164486
rect 481946 164218 481988 164454
rect 482224 164218 482266 164454
rect 481946 164134 482266 164218
rect 481946 163898 481988 164134
rect 482224 163898 482266 164134
rect 481946 163866 482266 163898
rect 489788 164454 490108 164486
rect 489788 164218 489830 164454
rect 490066 164218 490108 164454
rect 489788 164134 490108 164218
rect 489788 163898 489830 164134
rect 490066 163898 490108 164134
rect 489788 163866 490108 163898
rect 497630 164454 497950 164486
rect 497630 164218 497672 164454
rect 497908 164218 497950 164454
rect 497630 164134 497950 164218
rect 497630 163898 497672 164134
rect 497908 163898 497950 164134
rect 497630 163866 497950 163898
rect 508236 164454 508556 164486
rect 508236 164218 508278 164454
rect 508514 164218 508556 164454
rect 508236 164134 508556 164218
rect 508236 163898 508278 164134
rect 508514 163898 508556 164134
rect 508236 163866 508556 163898
rect 516078 164454 516398 164486
rect 516078 164218 516120 164454
rect 516356 164218 516398 164454
rect 516078 164134 516398 164218
rect 516078 163898 516120 164134
rect 516356 163898 516398 164134
rect 516078 163866 516398 163898
rect 523920 164454 524240 164486
rect 523920 164218 523962 164454
rect 524198 164218 524240 164454
rect 523920 164134 524240 164218
rect 523920 163898 523962 164134
rect 524198 163898 524240 164134
rect 523920 163866 524240 163898
rect 531762 164454 532082 164486
rect 531762 164218 531804 164454
rect 532040 164218 532082 164454
rect 531762 164134 532082 164218
rect 531762 163898 531804 164134
rect 532040 163898 532082 164134
rect 531762 163866 532082 163898
rect 542368 164454 542688 164486
rect 542368 164218 542410 164454
rect 542646 164218 542688 164454
rect 542368 164134 542688 164218
rect 542368 163898 542410 164134
rect 542646 163898 542688 164134
rect 542368 163866 542688 163898
rect 550210 164454 550530 164486
rect 550210 164218 550252 164454
rect 550488 164218 550530 164454
rect 550210 164134 550530 164218
rect 550210 163898 550252 164134
rect 550488 163898 550530 164134
rect 550210 163866 550530 163898
rect 558052 164454 558372 164486
rect 558052 164218 558094 164454
rect 558330 164218 558372 164454
rect 558052 164134 558372 164218
rect 558052 163898 558094 164134
rect 558330 163898 558372 164134
rect 558052 163866 558372 163898
rect 565894 164454 566214 164486
rect 565894 164218 565936 164454
rect 566172 164218 566214 164454
rect 565894 164134 566214 164218
rect 565894 163898 565936 164134
rect 566172 163898 566214 164134
rect 565894 163866 566214 163898
rect 574694 73813 574754 670651
rect 585310 668174 585930 677618
rect 585310 667938 585342 668174
rect 585578 667938 585662 668174
rect 585898 667938 585930 668174
rect 585310 667854 585930 667938
rect 585310 667618 585342 667854
rect 585578 667618 585662 667854
rect 585898 667618 585930 667854
rect 585310 658174 585930 667618
rect 585310 657938 585342 658174
rect 585578 657938 585662 658174
rect 585898 657938 585930 658174
rect 585310 657854 585930 657938
rect 585310 657618 585342 657854
rect 585578 657618 585662 657854
rect 585898 657618 585930 657854
rect 585310 648174 585930 657618
rect 585310 647938 585342 648174
rect 585578 647938 585662 648174
rect 585898 647938 585930 648174
rect 585310 647854 585930 647938
rect 585310 647618 585342 647854
rect 585578 647618 585662 647854
rect 585898 647618 585930 647854
rect 585310 638174 585930 647618
rect 585310 637938 585342 638174
rect 585578 637938 585662 638174
rect 585898 637938 585930 638174
rect 585310 637854 585930 637938
rect 585310 637618 585342 637854
rect 585578 637618 585662 637854
rect 585898 637618 585930 637854
rect 585310 628174 585930 637618
rect 585310 627938 585342 628174
rect 585578 627938 585662 628174
rect 585898 627938 585930 628174
rect 585310 627854 585930 627938
rect 585310 627618 585342 627854
rect 585578 627618 585662 627854
rect 585898 627618 585930 627854
rect 585310 618174 585930 627618
rect 585310 617938 585342 618174
rect 585578 617938 585662 618174
rect 585898 617938 585930 618174
rect 585310 617854 585930 617938
rect 585310 617618 585342 617854
rect 585578 617618 585662 617854
rect 585898 617618 585930 617854
rect 575979 617540 576045 617541
rect 575979 617476 575980 617540
rect 576044 617476 576045 617540
rect 575979 617475 576045 617476
rect 574875 511324 574941 511325
rect 574875 511260 574876 511324
rect 574940 511260 574941 511324
rect 574875 511259 574941 511260
rect 574691 73812 574757 73813
rect 574691 73748 574692 73812
rect 574756 73748 574757 73812
rect 574691 73747 574757 73748
rect 574878 71093 574938 511259
rect 575982 72453 576042 617475
rect 585310 608174 585930 617618
rect 585310 607938 585342 608174
rect 585578 607938 585662 608174
rect 585898 607938 585930 608174
rect 585310 607854 585930 607938
rect 585310 607618 585342 607854
rect 585578 607618 585662 607854
rect 585898 607618 585930 607854
rect 585310 598174 585930 607618
rect 585310 597938 585342 598174
rect 585578 597938 585662 598174
rect 585898 597938 585930 598174
rect 585310 597854 585930 597938
rect 585310 597618 585342 597854
rect 585578 597618 585662 597854
rect 585898 597618 585930 597854
rect 585310 588174 585930 597618
rect 585310 587938 585342 588174
rect 585578 587938 585662 588174
rect 585898 587938 585930 588174
rect 585310 587854 585930 587938
rect 585310 587618 585342 587854
rect 585578 587618 585662 587854
rect 585898 587618 585930 587854
rect 585310 578174 585930 587618
rect 585310 577938 585342 578174
rect 585578 577938 585662 578174
rect 585898 577938 585930 578174
rect 585310 577854 585930 577938
rect 585310 577618 585342 577854
rect 585578 577618 585662 577854
rect 585898 577618 585930 577854
rect 585310 568174 585930 577618
rect 585310 567938 585342 568174
rect 585578 567938 585662 568174
rect 585898 567938 585930 568174
rect 585310 567854 585930 567938
rect 585310 567618 585342 567854
rect 585578 567618 585662 567854
rect 585898 567618 585930 567854
rect 578739 564364 578805 564365
rect 578739 564300 578740 564364
rect 578804 564300 578805 564364
rect 578739 564299 578805 564300
rect 577451 404972 577517 404973
rect 577451 404908 577452 404972
rect 577516 404908 577517 404972
rect 577451 404907 577517 404908
rect 576163 245580 576229 245581
rect 576163 245516 576164 245580
rect 576228 245516 576229 245580
rect 576163 245515 576229 245516
rect 575979 72452 576045 72453
rect 575979 72388 575980 72452
rect 576044 72388 576045 72452
rect 575979 72387 576045 72388
rect 574875 71092 574941 71093
rect 574875 71028 574876 71092
rect 574940 71028 574941 71092
rect 574875 71027 574941 71028
rect 334755 68372 334821 68373
rect 334755 68308 334756 68372
rect 334820 68308 334821 68372
rect 334755 68307 334821 68308
rect 576166 21997 576226 245515
rect 577454 75173 577514 404907
rect 577635 351932 577701 351933
rect 577635 351868 577636 351932
rect 577700 351868 577701 351932
rect 577635 351867 577701 351868
rect 577638 153781 577698 351867
rect 578742 156637 578802 564299
rect 585310 558174 585930 567618
rect 585310 557938 585342 558174
rect 585578 557938 585662 558174
rect 585898 557938 585930 558174
rect 585310 557854 585930 557938
rect 585310 557618 585342 557854
rect 585578 557618 585662 557854
rect 585898 557618 585930 557854
rect 585310 548174 585930 557618
rect 585310 547938 585342 548174
rect 585578 547938 585662 548174
rect 585898 547938 585930 548174
rect 585310 547854 585930 547938
rect 585310 547618 585342 547854
rect 585578 547618 585662 547854
rect 585898 547618 585930 547854
rect 585310 538174 585930 547618
rect 585310 537938 585342 538174
rect 585578 537938 585662 538174
rect 585898 537938 585930 538174
rect 585310 537854 585930 537938
rect 585310 537618 585342 537854
rect 585578 537618 585662 537854
rect 585898 537618 585930 537854
rect 585310 528174 585930 537618
rect 585310 527938 585342 528174
rect 585578 527938 585662 528174
rect 585898 527938 585930 528174
rect 585310 527854 585930 527938
rect 585310 527618 585342 527854
rect 585578 527618 585662 527854
rect 585898 527618 585930 527854
rect 585310 518174 585930 527618
rect 585310 517938 585342 518174
rect 585578 517938 585662 518174
rect 585898 517938 585930 518174
rect 585310 517854 585930 517938
rect 585310 517618 585342 517854
rect 585578 517618 585662 517854
rect 585898 517618 585930 517854
rect 585310 508174 585930 517618
rect 585310 507938 585342 508174
rect 585578 507938 585662 508174
rect 585898 507938 585930 508174
rect 585310 507854 585930 507938
rect 585310 507618 585342 507854
rect 585578 507618 585662 507854
rect 585898 507618 585930 507854
rect 585310 498174 585930 507618
rect 585310 497938 585342 498174
rect 585578 497938 585662 498174
rect 585898 497938 585930 498174
rect 585310 497854 585930 497938
rect 585310 497618 585342 497854
rect 585578 497618 585662 497854
rect 585898 497618 585930 497854
rect 585310 488174 585930 497618
rect 585310 487938 585342 488174
rect 585578 487938 585662 488174
rect 585898 487938 585930 488174
rect 585310 487854 585930 487938
rect 585310 487618 585342 487854
rect 585578 487618 585662 487854
rect 585898 487618 585930 487854
rect 585310 478174 585930 487618
rect 585310 477938 585342 478174
rect 585578 477938 585662 478174
rect 585898 477938 585930 478174
rect 585310 477854 585930 477938
rect 585310 477618 585342 477854
rect 585578 477618 585662 477854
rect 585898 477618 585930 477854
rect 585310 468174 585930 477618
rect 585310 467938 585342 468174
rect 585578 467938 585662 468174
rect 585898 467938 585930 468174
rect 585310 467854 585930 467938
rect 585310 467618 585342 467854
rect 585578 467618 585662 467854
rect 585898 467618 585930 467854
rect 585310 458174 585930 467618
rect 578923 458148 578989 458149
rect 578923 458084 578924 458148
rect 578988 458084 578989 458148
rect 578923 458083 578989 458084
rect 578739 156636 578805 156637
rect 578739 156572 578740 156636
rect 578804 156572 578805 156636
rect 578739 156571 578805 156572
rect 577635 153780 577701 153781
rect 577635 153716 577636 153780
rect 577700 153716 577701 153780
rect 577635 153715 577701 153716
rect 577451 75172 577517 75173
rect 577451 75108 577452 75172
rect 577516 75108 577517 75172
rect 577451 75107 577517 75108
rect 578926 69597 578986 458083
rect 585310 457938 585342 458174
rect 585578 457938 585662 458174
rect 585898 457938 585930 458174
rect 585310 457854 585930 457938
rect 585310 457618 585342 457854
rect 585578 457618 585662 457854
rect 585898 457618 585930 457854
rect 585310 448174 585930 457618
rect 585310 447938 585342 448174
rect 585578 447938 585662 448174
rect 585898 447938 585930 448174
rect 585310 447854 585930 447938
rect 585310 447618 585342 447854
rect 585578 447618 585662 447854
rect 585898 447618 585930 447854
rect 585310 438174 585930 447618
rect 585310 437938 585342 438174
rect 585578 437938 585662 438174
rect 585898 437938 585930 438174
rect 585310 437854 585930 437938
rect 585310 437618 585342 437854
rect 585578 437618 585662 437854
rect 585898 437618 585930 437854
rect 585310 428174 585930 437618
rect 585310 427938 585342 428174
rect 585578 427938 585662 428174
rect 585898 427938 585930 428174
rect 585310 427854 585930 427938
rect 585310 427618 585342 427854
rect 585578 427618 585662 427854
rect 585898 427618 585930 427854
rect 585310 418174 585930 427618
rect 585310 417938 585342 418174
rect 585578 417938 585662 418174
rect 585898 417938 585930 418174
rect 585310 417854 585930 417938
rect 585310 417618 585342 417854
rect 585578 417618 585662 417854
rect 585898 417618 585930 417854
rect 585310 408174 585930 417618
rect 585310 407938 585342 408174
rect 585578 407938 585662 408174
rect 585898 407938 585930 408174
rect 585310 407854 585930 407938
rect 585310 407618 585342 407854
rect 585578 407618 585662 407854
rect 585898 407618 585930 407854
rect 585310 398174 585930 407618
rect 585310 397938 585342 398174
rect 585578 397938 585662 398174
rect 585898 397938 585930 398174
rect 585310 397854 585930 397938
rect 585310 397618 585342 397854
rect 585578 397618 585662 397854
rect 585898 397618 585930 397854
rect 585310 388174 585930 397618
rect 585310 387938 585342 388174
rect 585578 387938 585662 388174
rect 585898 387938 585930 388174
rect 585310 387854 585930 387938
rect 585310 387618 585342 387854
rect 585578 387618 585662 387854
rect 585898 387618 585930 387854
rect 585310 378174 585930 387618
rect 585310 377938 585342 378174
rect 585578 377938 585662 378174
rect 585898 377938 585930 378174
rect 585310 377854 585930 377938
rect 585310 377618 585342 377854
rect 585578 377618 585662 377854
rect 585898 377618 585930 377854
rect 585310 368174 585930 377618
rect 585310 367938 585342 368174
rect 585578 367938 585662 368174
rect 585898 367938 585930 368174
rect 585310 367854 585930 367938
rect 585310 367618 585342 367854
rect 585578 367618 585662 367854
rect 585898 367618 585930 367854
rect 585310 358174 585930 367618
rect 585310 357938 585342 358174
rect 585578 357938 585662 358174
rect 585898 357938 585930 358174
rect 585310 357854 585930 357938
rect 585310 357618 585342 357854
rect 585578 357618 585662 357854
rect 585898 357618 585930 357854
rect 585310 348174 585930 357618
rect 585310 347938 585342 348174
rect 585578 347938 585662 348174
rect 585898 347938 585930 348174
rect 585310 347854 585930 347938
rect 585310 347618 585342 347854
rect 585578 347618 585662 347854
rect 585898 347618 585930 347854
rect 585310 338174 585930 347618
rect 585310 337938 585342 338174
rect 585578 337938 585662 338174
rect 585898 337938 585930 338174
rect 585310 337854 585930 337938
rect 585310 337618 585342 337854
rect 585578 337618 585662 337854
rect 585898 337618 585930 337854
rect 585310 328174 585930 337618
rect 585310 327938 585342 328174
rect 585578 327938 585662 328174
rect 585898 327938 585930 328174
rect 585310 327854 585930 327938
rect 585310 327618 585342 327854
rect 585578 327618 585662 327854
rect 585898 327618 585930 327854
rect 585310 318174 585930 327618
rect 585310 317938 585342 318174
rect 585578 317938 585662 318174
rect 585898 317938 585930 318174
rect 585310 317854 585930 317938
rect 585310 317618 585342 317854
rect 585578 317618 585662 317854
rect 585898 317618 585930 317854
rect 585310 308174 585930 317618
rect 585310 307938 585342 308174
rect 585578 307938 585662 308174
rect 585898 307938 585930 308174
rect 585310 307854 585930 307938
rect 585310 307618 585342 307854
rect 585578 307618 585662 307854
rect 585898 307618 585930 307854
rect 580211 298756 580277 298757
rect 580211 298692 580212 298756
rect 580276 298692 580277 298756
rect 580211 298691 580277 298692
rect 580214 155277 580274 298691
rect 585310 298174 585930 307618
rect 585310 297938 585342 298174
rect 585578 297938 585662 298174
rect 585898 297938 585930 298174
rect 585310 297854 585930 297938
rect 585310 297618 585342 297854
rect 585578 297618 585662 297854
rect 585898 297618 585930 297854
rect 585310 288174 585930 297618
rect 585310 287938 585342 288174
rect 585578 287938 585662 288174
rect 585898 287938 585930 288174
rect 585310 287854 585930 287938
rect 585310 287618 585342 287854
rect 585578 287618 585662 287854
rect 585898 287618 585930 287854
rect 585310 278174 585930 287618
rect 585310 277938 585342 278174
rect 585578 277938 585662 278174
rect 585898 277938 585930 278174
rect 585310 277854 585930 277938
rect 585310 277618 585342 277854
rect 585578 277618 585662 277854
rect 585898 277618 585930 277854
rect 585310 268174 585930 277618
rect 585310 267938 585342 268174
rect 585578 267938 585662 268174
rect 585898 267938 585930 268174
rect 585310 267854 585930 267938
rect 585310 267618 585342 267854
rect 585578 267618 585662 267854
rect 585898 267618 585930 267854
rect 585310 258174 585930 267618
rect 585310 257938 585342 258174
rect 585578 257938 585662 258174
rect 585898 257938 585930 258174
rect 585310 257854 585930 257938
rect 585310 257618 585342 257854
rect 585578 257618 585662 257854
rect 585898 257618 585930 257854
rect 585310 248174 585930 257618
rect 585310 247938 585342 248174
rect 585578 247938 585662 248174
rect 585898 247938 585930 248174
rect 585310 247854 585930 247938
rect 585310 247618 585342 247854
rect 585578 247618 585662 247854
rect 585898 247618 585930 247854
rect 585310 238174 585930 247618
rect 585310 237938 585342 238174
rect 585578 237938 585662 238174
rect 585898 237938 585930 238174
rect 585310 237854 585930 237938
rect 585310 237618 585342 237854
rect 585578 237618 585662 237854
rect 585898 237618 585930 237854
rect 580579 232388 580645 232389
rect 580579 232324 580580 232388
rect 580644 232324 580645 232388
rect 580579 232323 580645 232324
rect 580582 192541 580642 232323
rect 585310 228174 585930 237618
rect 585310 227938 585342 228174
rect 585578 227938 585662 228174
rect 585898 227938 585930 228174
rect 585310 227854 585930 227938
rect 585310 227618 585342 227854
rect 585578 227618 585662 227854
rect 585898 227618 585930 227854
rect 580763 219060 580829 219061
rect 580763 218996 580764 219060
rect 580828 218996 580829 219060
rect 580763 218995 580829 218996
rect 580579 192540 580645 192541
rect 580579 192476 580580 192540
rect 580644 192476 580645 192540
rect 580579 192475 580645 192476
rect 580582 179213 580642 192475
rect 580579 179212 580645 179213
rect 580579 179148 580580 179212
rect 580644 179148 580645 179212
rect 580579 179147 580645 179148
rect 580582 174589 580642 179147
rect 580579 174588 580645 174589
rect 580579 174524 580580 174588
rect 580644 174524 580645 174588
rect 580579 174523 580645 174524
rect 580211 155276 580277 155277
rect 580211 155212 580212 155276
rect 580276 155212 580277 155276
rect 580211 155211 580277 155212
rect 578923 69596 578989 69597
rect 578923 69532 578924 69596
rect 578988 69532 578989 69596
rect 578923 69531 578989 69532
rect 576163 21996 576229 21997
rect 576163 21932 576164 21996
rect 576228 21932 576229 21996
rect 576163 21931 576229 21932
rect 306603 20636 306669 20637
rect 306603 20572 306604 20636
rect 306668 20572 306669 20636
rect 306603 20571 306669 20572
rect 311019 20636 311085 20637
rect 311019 20572 311020 20636
rect 311084 20572 311085 20636
rect 311019 20571 311085 20572
rect 279003 19276 279069 19277
rect 279003 19212 279004 19276
rect 279068 19212 279069 19276
rect 279003 19211 279069 19212
rect 272379 19140 272445 19141
rect 272379 19076 272380 19140
rect 272444 19076 272445 19140
rect 272379 19075 272445 19076
rect 278635 19140 278701 19141
rect 278635 19076 278636 19140
rect 278700 19076 278701 19140
rect 278635 19075 278701 19076
rect 271091 19004 271157 19005
rect 271091 18940 271092 19004
rect 271156 18940 271157 19004
rect 271091 18939 271157 18940
rect 580766 3501 580826 218995
rect 585310 218174 585930 227618
rect 585310 217938 585342 218174
rect 585578 217938 585662 218174
rect 585898 217938 585930 218174
rect 585310 217854 585930 217938
rect 585310 217618 585342 217854
rect 585578 217618 585662 217854
rect 585898 217618 585930 217854
rect 585310 208174 585930 217618
rect 585310 207938 585342 208174
rect 585578 207938 585662 208174
rect 585898 207938 585930 208174
rect 585310 207854 585930 207938
rect 585310 207618 585342 207854
rect 585578 207618 585662 207854
rect 585898 207618 585930 207854
rect 585310 198174 585930 207618
rect 585310 197938 585342 198174
rect 585578 197938 585662 198174
rect 585898 197938 585930 198174
rect 585310 197854 585930 197938
rect 585310 197618 585342 197854
rect 585578 197618 585662 197854
rect 585898 197618 585930 197854
rect 585310 188174 585930 197618
rect 585310 187938 585342 188174
rect 585578 187938 585662 188174
rect 585898 187938 585930 188174
rect 585310 187854 585930 187938
rect 585310 187618 585342 187854
rect 585578 187618 585662 187854
rect 585898 187618 585930 187854
rect 585310 178174 585930 187618
rect 585310 177938 585342 178174
rect 585578 177938 585662 178174
rect 585898 177938 585930 178174
rect 585310 177854 585930 177938
rect 585310 177618 585342 177854
rect 585578 177618 585662 177854
rect 585898 177618 585930 177854
rect 585310 168174 585930 177618
rect 585310 167938 585342 168174
rect 585578 167938 585662 168174
rect 585898 167938 585930 168174
rect 585310 167854 585930 167938
rect 585310 167618 585342 167854
rect 585578 167618 585662 167854
rect 585898 167618 585930 167854
rect 585310 158174 585930 167618
rect 585310 157938 585342 158174
rect 585578 157938 585662 158174
rect 585898 157938 585930 158174
rect 585310 157854 585930 157938
rect 585310 157618 585342 157854
rect 585578 157618 585662 157854
rect 585898 157618 585930 157854
rect 585310 148174 585930 157618
rect 585310 147938 585342 148174
rect 585578 147938 585662 148174
rect 585898 147938 585930 148174
rect 585310 147854 585930 147938
rect 585310 147618 585342 147854
rect 585578 147618 585662 147854
rect 585898 147618 585930 147854
rect 585310 138174 585930 147618
rect 585310 137938 585342 138174
rect 585578 137938 585662 138174
rect 585898 137938 585930 138174
rect 585310 137854 585930 137938
rect 585310 137618 585342 137854
rect 585578 137618 585662 137854
rect 585898 137618 585930 137854
rect 585310 128174 585930 137618
rect 585310 127938 585342 128174
rect 585578 127938 585662 128174
rect 585898 127938 585930 128174
rect 585310 127854 585930 127938
rect 585310 127618 585342 127854
rect 585578 127618 585662 127854
rect 585898 127618 585930 127854
rect 585310 118174 585930 127618
rect 585310 117938 585342 118174
rect 585578 117938 585662 118174
rect 585898 117938 585930 118174
rect 585310 117854 585930 117938
rect 585310 117618 585342 117854
rect 585578 117618 585662 117854
rect 585898 117618 585930 117854
rect 585310 108174 585930 117618
rect 585310 107938 585342 108174
rect 585578 107938 585662 108174
rect 585898 107938 585930 108174
rect 585310 107854 585930 107938
rect 585310 107618 585342 107854
rect 585578 107618 585662 107854
rect 585898 107618 585930 107854
rect 585310 98174 585930 107618
rect 585310 97938 585342 98174
rect 585578 97938 585662 98174
rect 585898 97938 585930 98174
rect 585310 97854 585930 97938
rect 585310 97618 585342 97854
rect 585578 97618 585662 97854
rect 585898 97618 585930 97854
rect 585310 88174 585930 97618
rect 585310 87938 585342 88174
rect 585578 87938 585662 88174
rect 585898 87938 585930 88174
rect 585310 87854 585930 87938
rect 585310 87618 585342 87854
rect 585578 87618 585662 87854
rect 585898 87618 585930 87854
rect 585310 78174 585930 87618
rect 585310 77938 585342 78174
rect 585578 77938 585662 78174
rect 585898 77938 585930 78174
rect 585310 77854 585930 77938
rect 585310 77618 585342 77854
rect 585578 77618 585662 77854
rect 585898 77618 585930 77854
rect 585310 68174 585930 77618
rect 585310 67938 585342 68174
rect 585578 67938 585662 68174
rect 585898 67938 585930 68174
rect 585310 67854 585930 67938
rect 585310 67618 585342 67854
rect 585578 67618 585662 67854
rect 585898 67618 585930 67854
rect 585310 58174 585930 67618
rect 585310 57938 585342 58174
rect 585578 57938 585662 58174
rect 585898 57938 585930 58174
rect 585310 57854 585930 57938
rect 585310 57618 585342 57854
rect 585578 57618 585662 57854
rect 585898 57618 585930 57854
rect 585310 48174 585930 57618
rect 585310 47938 585342 48174
rect 585578 47938 585662 48174
rect 585898 47938 585930 48174
rect 585310 47854 585930 47938
rect 585310 47618 585342 47854
rect 585578 47618 585662 47854
rect 585898 47618 585930 47854
rect 585310 38174 585930 47618
rect 585310 37938 585342 38174
rect 585578 37938 585662 38174
rect 585898 37938 585930 38174
rect 585310 37854 585930 37938
rect 585310 37618 585342 37854
rect 585578 37618 585662 37854
rect 585898 37618 585930 37854
rect 580763 3500 580829 3501
rect 580763 3436 580764 3500
rect 580828 3436 580829 3500
rect 580763 3435 580829 3436
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 585310 -346 585930 37618
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 694454 586890 705242
rect 586270 694218 586302 694454
rect 586538 694218 586622 694454
rect 586858 694218 586890 694454
rect 586270 694134 586890 694218
rect 586270 693898 586302 694134
rect 586538 693898 586622 694134
rect 586858 693898 586890 694134
rect 586270 684454 586890 693898
rect 586270 684218 586302 684454
rect 586538 684218 586622 684454
rect 586858 684218 586890 684454
rect 586270 684134 586890 684218
rect 586270 683898 586302 684134
rect 586538 683898 586622 684134
rect 586858 683898 586890 684134
rect 586270 674454 586890 683898
rect 586270 674218 586302 674454
rect 586538 674218 586622 674454
rect 586858 674218 586890 674454
rect 586270 674134 586890 674218
rect 586270 673898 586302 674134
rect 586538 673898 586622 674134
rect 586858 673898 586890 674134
rect 586270 664454 586890 673898
rect 586270 664218 586302 664454
rect 586538 664218 586622 664454
rect 586858 664218 586890 664454
rect 586270 664134 586890 664218
rect 586270 663898 586302 664134
rect 586538 663898 586622 664134
rect 586858 663898 586890 664134
rect 586270 654454 586890 663898
rect 586270 654218 586302 654454
rect 586538 654218 586622 654454
rect 586858 654218 586890 654454
rect 586270 654134 586890 654218
rect 586270 653898 586302 654134
rect 586538 653898 586622 654134
rect 586858 653898 586890 654134
rect 586270 644454 586890 653898
rect 586270 644218 586302 644454
rect 586538 644218 586622 644454
rect 586858 644218 586890 644454
rect 586270 644134 586890 644218
rect 586270 643898 586302 644134
rect 586538 643898 586622 644134
rect 586858 643898 586890 644134
rect 586270 634454 586890 643898
rect 586270 634218 586302 634454
rect 586538 634218 586622 634454
rect 586858 634218 586890 634454
rect 586270 634134 586890 634218
rect 586270 633898 586302 634134
rect 586538 633898 586622 634134
rect 586858 633898 586890 634134
rect 586270 624454 586890 633898
rect 586270 624218 586302 624454
rect 586538 624218 586622 624454
rect 586858 624218 586890 624454
rect 586270 624134 586890 624218
rect 586270 623898 586302 624134
rect 586538 623898 586622 624134
rect 586858 623898 586890 624134
rect 586270 614454 586890 623898
rect 586270 614218 586302 614454
rect 586538 614218 586622 614454
rect 586858 614218 586890 614454
rect 586270 614134 586890 614218
rect 586270 613898 586302 614134
rect 586538 613898 586622 614134
rect 586858 613898 586890 614134
rect 586270 604454 586890 613898
rect 586270 604218 586302 604454
rect 586538 604218 586622 604454
rect 586858 604218 586890 604454
rect 586270 604134 586890 604218
rect 586270 603898 586302 604134
rect 586538 603898 586622 604134
rect 586858 603898 586890 604134
rect 586270 594454 586890 603898
rect 586270 594218 586302 594454
rect 586538 594218 586622 594454
rect 586858 594218 586890 594454
rect 586270 594134 586890 594218
rect 586270 593898 586302 594134
rect 586538 593898 586622 594134
rect 586858 593898 586890 594134
rect 586270 584454 586890 593898
rect 586270 584218 586302 584454
rect 586538 584218 586622 584454
rect 586858 584218 586890 584454
rect 586270 584134 586890 584218
rect 586270 583898 586302 584134
rect 586538 583898 586622 584134
rect 586858 583898 586890 584134
rect 586270 574454 586890 583898
rect 586270 574218 586302 574454
rect 586538 574218 586622 574454
rect 586858 574218 586890 574454
rect 586270 574134 586890 574218
rect 586270 573898 586302 574134
rect 586538 573898 586622 574134
rect 586858 573898 586890 574134
rect 586270 564454 586890 573898
rect 586270 564218 586302 564454
rect 586538 564218 586622 564454
rect 586858 564218 586890 564454
rect 586270 564134 586890 564218
rect 586270 563898 586302 564134
rect 586538 563898 586622 564134
rect 586858 563898 586890 564134
rect 586270 554454 586890 563898
rect 586270 554218 586302 554454
rect 586538 554218 586622 554454
rect 586858 554218 586890 554454
rect 586270 554134 586890 554218
rect 586270 553898 586302 554134
rect 586538 553898 586622 554134
rect 586858 553898 586890 554134
rect 586270 544454 586890 553898
rect 586270 544218 586302 544454
rect 586538 544218 586622 544454
rect 586858 544218 586890 544454
rect 586270 544134 586890 544218
rect 586270 543898 586302 544134
rect 586538 543898 586622 544134
rect 586858 543898 586890 544134
rect 586270 534454 586890 543898
rect 586270 534218 586302 534454
rect 586538 534218 586622 534454
rect 586858 534218 586890 534454
rect 586270 534134 586890 534218
rect 586270 533898 586302 534134
rect 586538 533898 586622 534134
rect 586858 533898 586890 534134
rect 586270 524454 586890 533898
rect 586270 524218 586302 524454
rect 586538 524218 586622 524454
rect 586858 524218 586890 524454
rect 586270 524134 586890 524218
rect 586270 523898 586302 524134
rect 586538 523898 586622 524134
rect 586858 523898 586890 524134
rect 586270 514454 586890 523898
rect 586270 514218 586302 514454
rect 586538 514218 586622 514454
rect 586858 514218 586890 514454
rect 586270 514134 586890 514218
rect 586270 513898 586302 514134
rect 586538 513898 586622 514134
rect 586858 513898 586890 514134
rect 586270 504454 586890 513898
rect 586270 504218 586302 504454
rect 586538 504218 586622 504454
rect 586858 504218 586890 504454
rect 586270 504134 586890 504218
rect 586270 503898 586302 504134
rect 586538 503898 586622 504134
rect 586858 503898 586890 504134
rect 586270 494454 586890 503898
rect 586270 494218 586302 494454
rect 586538 494218 586622 494454
rect 586858 494218 586890 494454
rect 586270 494134 586890 494218
rect 586270 493898 586302 494134
rect 586538 493898 586622 494134
rect 586858 493898 586890 494134
rect 586270 484454 586890 493898
rect 586270 484218 586302 484454
rect 586538 484218 586622 484454
rect 586858 484218 586890 484454
rect 586270 484134 586890 484218
rect 586270 483898 586302 484134
rect 586538 483898 586622 484134
rect 586858 483898 586890 484134
rect 586270 474454 586890 483898
rect 586270 474218 586302 474454
rect 586538 474218 586622 474454
rect 586858 474218 586890 474454
rect 586270 474134 586890 474218
rect 586270 473898 586302 474134
rect 586538 473898 586622 474134
rect 586858 473898 586890 474134
rect 586270 464454 586890 473898
rect 586270 464218 586302 464454
rect 586538 464218 586622 464454
rect 586858 464218 586890 464454
rect 586270 464134 586890 464218
rect 586270 463898 586302 464134
rect 586538 463898 586622 464134
rect 586858 463898 586890 464134
rect 586270 454454 586890 463898
rect 586270 454218 586302 454454
rect 586538 454218 586622 454454
rect 586858 454218 586890 454454
rect 586270 454134 586890 454218
rect 586270 453898 586302 454134
rect 586538 453898 586622 454134
rect 586858 453898 586890 454134
rect 586270 444454 586890 453898
rect 586270 444218 586302 444454
rect 586538 444218 586622 444454
rect 586858 444218 586890 444454
rect 586270 444134 586890 444218
rect 586270 443898 586302 444134
rect 586538 443898 586622 444134
rect 586858 443898 586890 444134
rect 586270 434454 586890 443898
rect 586270 434218 586302 434454
rect 586538 434218 586622 434454
rect 586858 434218 586890 434454
rect 586270 434134 586890 434218
rect 586270 433898 586302 434134
rect 586538 433898 586622 434134
rect 586858 433898 586890 434134
rect 586270 424454 586890 433898
rect 586270 424218 586302 424454
rect 586538 424218 586622 424454
rect 586858 424218 586890 424454
rect 586270 424134 586890 424218
rect 586270 423898 586302 424134
rect 586538 423898 586622 424134
rect 586858 423898 586890 424134
rect 586270 414454 586890 423898
rect 586270 414218 586302 414454
rect 586538 414218 586622 414454
rect 586858 414218 586890 414454
rect 586270 414134 586890 414218
rect 586270 413898 586302 414134
rect 586538 413898 586622 414134
rect 586858 413898 586890 414134
rect 586270 404454 586890 413898
rect 586270 404218 586302 404454
rect 586538 404218 586622 404454
rect 586858 404218 586890 404454
rect 586270 404134 586890 404218
rect 586270 403898 586302 404134
rect 586538 403898 586622 404134
rect 586858 403898 586890 404134
rect 586270 394454 586890 403898
rect 586270 394218 586302 394454
rect 586538 394218 586622 394454
rect 586858 394218 586890 394454
rect 586270 394134 586890 394218
rect 586270 393898 586302 394134
rect 586538 393898 586622 394134
rect 586858 393898 586890 394134
rect 586270 384454 586890 393898
rect 586270 384218 586302 384454
rect 586538 384218 586622 384454
rect 586858 384218 586890 384454
rect 586270 384134 586890 384218
rect 586270 383898 586302 384134
rect 586538 383898 586622 384134
rect 586858 383898 586890 384134
rect 586270 374454 586890 383898
rect 586270 374218 586302 374454
rect 586538 374218 586622 374454
rect 586858 374218 586890 374454
rect 586270 374134 586890 374218
rect 586270 373898 586302 374134
rect 586538 373898 586622 374134
rect 586858 373898 586890 374134
rect 586270 364454 586890 373898
rect 586270 364218 586302 364454
rect 586538 364218 586622 364454
rect 586858 364218 586890 364454
rect 586270 364134 586890 364218
rect 586270 363898 586302 364134
rect 586538 363898 586622 364134
rect 586858 363898 586890 364134
rect 586270 354454 586890 363898
rect 586270 354218 586302 354454
rect 586538 354218 586622 354454
rect 586858 354218 586890 354454
rect 586270 354134 586890 354218
rect 586270 353898 586302 354134
rect 586538 353898 586622 354134
rect 586858 353898 586890 354134
rect 586270 344454 586890 353898
rect 586270 344218 586302 344454
rect 586538 344218 586622 344454
rect 586858 344218 586890 344454
rect 586270 344134 586890 344218
rect 586270 343898 586302 344134
rect 586538 343898 586622 344134
rect 586858 343898 586890 344134
rect 586270 334454 586890 343898
rect 586270 334218 586302 334454
rect 586538 334218 586622 334454
rect 586858 334218 586890 334454
rect 586270 334134 586890 334218
rect 586270 333898 586302 334134
rect 586538 333898 586622 334134
rect 586858 333898 586890 334134
rect 586270 324454 586890 333898
rect 586270 324218 586302 324454
rect 586538 324218 586622 324454
rect 586858 324218 586890 324454
rect 586270 324134 586890 324218
rect 586270 323898 586302 324134
rect 586538 323898 586622 324134
rect 586858 323898 586890 324134
rect 586270 314454 586890 323898
rect 586270 314218 586302 314454
rect 586538 314218 586622 314454
rect 586858 314218 586890 314454
rect 586270 314134 586890 314218
rect 586270 313898 586302 314134
rect 586538 313898 586622 314134
rect 586858 313898 586890 314134
rect 586270 304454 586890 313898
rect 586270 304218 586302 304454
rect 586538 304218 586622 304454
rect 586858 304218 586890 304454
rect 586270 304134 586890 304218
rect 586270 303898 586302 304134
rect 586538 303898 586622 304134
rect 586858 303898 586890 304134
rect 586270 294454 586890 303898
rect 586270 294218 586302 294454
rect 586538 294218 586622 294454
rect 586858 294218 586890 294454
rect 586270 294134 586890 294218
rect 586270 293898 586302 294134
rect 586538 293898 586622 294134
rect 586858 293898 586890 294134
rect 586270 284454 586890 293898
rect 586270 284218 586302 284454
rect 586538 284218 586622 284454
rect 586858 284218 586890 284454
rect 586270 284134 586890 284218
rect 586270 283898 586302 284134
rect 586538 283898 586622 284134
rect 586858 283898 586890 284134
rect 586270 274454 586890 283898
rect 586270 274218 586302 274454
rect 586538 274218 586622 274454
rect 586858 274218 586890 274454
rect 586270 274134 586890 274218
rect 586270 273898 586302 274134
rect 586538 273898 586622 274134
rect 586858 273898 586890 274134
rect 586270 264454 586890 273898
rect 586270 264218 586302 264454
rect 586538 264218 586622 264454
rect 586858 264218 586890 264454
rect 586270 264134 586890 264218
rect 586270 263898 586302 264134
rect 586538 263898 586622 264134
rect 586858 263898 586890 264134
rect 586270 254454 586890 263898
rect 586270 254218 586302 254454
rect 586538 254218 586622 254454
rect 586858 254218 586890 254454
rect 586270 254134 586890 254218
rect 586270 253898 586302 254134
rect 586538 253898 586622 254134
rect 586858 253898 586890 254134
rect 586270 244454 586890 253898
rect 586270 244218 586302 244454
rect 586538 244218 586622 244454
rect 586858 244218 586890 244454
rect 586270 244134 586890 244218
rect 586270 243898 586302 244134
rect 586538 243898 586622 244134
rect 586858 243898 586890 244134
rect 586270 234454 586890 243898
rect 586270 234218 586302 234454
rect 586538 234218 586622 234454
rect 586858 234218 586890 234454
rect 586270 234134 586890 234218
rect 586270 233898 586302 234134
rect 586538 233898 586622 234134
rect 586858 233898 586890 234134
rect 586270 224454 586890 233898
rect 586270 224218 586302 224454
rect 586538 224218 586622 224454
rect 586858 224218 586890 224454
rect 586270 224134 586890 224218
rect 586270 223898 586302 224134
rect 586538 223898 586622 224134
rect 586858 223898 586890 224134
rect 586270 214454 586890 223898
rect 586270 214218 586302 214454
rect 586538 214218 586622 214454
rect 586858 214218 586890 214454
rect 586270 214134 586890 214218
rect 586270 213898 586302 214134
rect 586538 213898 586622 214134
rect 586858 213898 586890 214134
rect 586270 204454 586890 213898
rect 586270 204218 586302 204454
rect 586538 204218 586622 204454
rect 586858 204218 586890 204454
rect 586270 204134 586890 204218
rect 586270 203898 586302 204134
rect 586538 203898 586622 204134
rect 586858 203898 586890 204134
rect 586270 194454 586890 203898
rect 586270 194218 586302 194454
rect 586538 194218 586622 194454
rect 586858 194218 586890 194454
rect 586270 194134 586890 194218
rect 586270 193898 586302 194134
rect 586538 193898 586622 194134
rect 586858 193898 586890 194134
rect 586270 184454 586890 193898
rect 586270 184218 586302 184454
rect 586538 184218 586622 184454
rect 586858 184218 586890 184454
rect 586270 184134 586890 184218
rect 586270 183898 586302 184134
rect 586538 183898 586622 184134
rect 586858 183898 586890 184134
rect 586270 174454 586890 183898
rect 586270 174218 586302 174454
rect 586538 174218 586622 174454
rect 586858 174218 586890 174454
rect 586270 174134 586890 174218
rect 586270 173898 586302 174134
rect 586538 173898 586622 174134
rect 586858 173898 586890 174134
rect 586270 164454 586890 173898
rect 586270 164218 586302 164454
rect 586538 164218 586622 164454
rect 586858 164218 586890 164454
rect 586270 164134 586890 164218
rect 586270 163898 586302 164134
rect 586538 163898 586622 164134
rect 586858 163898 586890 164134
rect 586270 154454 586890 163898
rect 586270 154218 586302 154454
rect 586538 154218 586622 154454
rect 586858 154218 586890 154454
rect 586270 154134 586890 154218
rect 586270 153898 586302 154134
rect 586538 153898 586622 154134
rect 586858 153898 586890 154134
rect 586270 144454 586890 153898
rect 586270 144218 586302 144454
rect 586538 144218 586622 144454
rect 586858 144218 586890 144454
rect 586270 144134 586890 144218
rect 586270 143898 586302 144134
rect 586538 143898 586622 144134
rect 586858 143898 586890 144134
rect 586270 134454 586890 143898
rect 586270 134218 586302 134454
rect 586538 134218 586622 134454
rect 586858 134218 586890 134454
rect 586270 134134 586890 134218
rect 586270 133898 586302 134134
rect 586538 133898 586622 134134
rect 586858 133898 586890 134134
rect 586270 124454 586890 133898
rect 586270 124218 586302 124454
rect 586538 124218 586622 124454
rect 586858 124218 586890 124454
rect 586270 124134 586890 124218
rect 586270 123898 586302 124134
rect 586538 123898 586622 124134
rect 586858 123898 586890 124134
rect 586270 114454 586890 123898
rect 586270 114218 586302 114454
rect 586538 114218 586622 114454
rect 586858 114218 586890 114454
rect 586270 114134 586890 114218
rect 586270 113898 586302 114134
rect 586538 113898 586622 114134
rect 586858 113898 586890 114134
rect 586270 104454 586890 113898
rect 586270 104218 586302 104454
rect 586538 104218 586622 104454
rect 586858 104218 586890 104454
rect 586270 104134 586890 104218
rect 586270 103898 586302 104134
rect 586538 103898 586622 104134
rect 586858 103898 586890 104134
rect 586270 94454 586890 103898
rect 586270 94218 586302 94454
rect 586538 94218 586622 94454
rect 586858 94218 586890 94454
rect 586270 94134 586890 94218
rect 586270 93898 586302 94134
rect 586538 93898 586622 94134
rect 586858 93898 586890 94134
rect 586270 84454 586890 93898
rect 586270 84218 586302 84454
rect 586538 84218 586622 84454
rect 586858 84218 586890 84454
rect 586270 84134 586890 84218
rect 586270 83898 586302 84134
rect 586538 83898 586622 84134
rect 586858 83898 586890 84134
rect 586270 74454 586890 83898
rect 586270 74218 586302 74454
rect 586538 74218 586622 74454
rect 586858 74218 586890 74454
rect 586270 74134 586890 74218
rect 586270 73898 586302 74134
rect 586538 73898 586622 74134
rect 586858 73898 586890 74134
rect 586270 64454 586890 73898
rect 586270 64218 586302 64454
rect 586538 64218 586622 64454
rect 586858 64218 586890 64454
rect 586270 64134 586890 64218
rect 586270 63898 586302 64134
rect 586538 63898 586622 64134
rect 586858 63898 586890 64134
rect 586270 54454 586890 63898
rect 586270 54218 586302 54454
rect 586538 54218 586622 54454
rect 586858 54218 586890 54454
rect 586270 54134 586890 54218
rect 586270 53898 586302 54134
rect 586538 53898 586622 54134
rect 586858 53898 586890 54134
rect 586270 44454 586890 53898
rect 586270 44218 586302 44454
rect 586538 44218 586622 44454
rect 586858 44218 586890 44454
rect 586270 44134 586890 44218
rect 586270 43898 586302 44134
rect 586538 43898 586622 44134
rect 586858 43898 586890 44134
rect 586270 34454 586890 43898
rect 586270 34218 586302 34454
rect 586538 34218 586622 34454
rect 586858 34218 586890 34454
rect 586270 34134 586890 34218
rect 586270 33898 586302 34134
rect 586538 33898 586622 34134
rect 586858 33898 586890 34134
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 586270 -1306 586890 33898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 587230 -2266 587850 706202
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 588190 -3226 588810 707162
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 589150 -4186 589770 708122
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 590110 -5146 590730 709082
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 591070 -6106 591690 710042
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 592030 -7066 592650 711002
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect -2934 694218 -2698 694454
rect -2614 694218 -2378 694454
rect -2934 693898 -2698 694134
rect -2614 693898 -2378 694134
rect -2934 684218 -2698 684454
rect -2614 684218 -2378 684454
rect -2934 683898 -2698 684134
rect -2614 683898 -2378 684134
rect -2934 674218 -2698 674454
rect -2614 674218 -2378 674454
rect -2934 673898 -2698 674134
rect -2614 673898 -2378 674134
rect -2934 664218 -2698 664454
rect -2614 664218 -2378 664454
rect -2934 663898 -2698 664134
rect -2614 663898 -2378 664134
rect -2934 654218 -2698 654454
rect -2614 654218 -2378 654454
rect -2934 653898 -2698 654134
rect -2614 653898 -2378 654134
rect -2934 644218 -2698 644454
rect -2614 644218 -2378 644454
rect -2934 643898 -2698 644134
rect -2614 643898 -2378 644134
rect -2934 634218 -2698 634454
rect -2614 634218 -2378 634454
rect -2934 633898 -2698 634134
rect -2614 633898 -2378 634134
rect -2934 624218 -2698 624454
rect -2614 624218 -2378 624454
rect -2934 623898 -2698 624134
rect -2614 623898 -2378 624134
rect -2934 614218 -2698 614454
rect -2614 614218 -2378 614454
rect -2934 613898 -2698 614134
rect -2614 613898 -2378 614134
rect -2934 604218 -2698 604454
rect -2614 604218 -2378 604454
rect -2934 603898 -2698 604134
rect -2614 603898 -2378 604134
rect -2934 594218 -2698 594454
rect -2614 594218 -2378 594454
rect -2934 593898 -2698 594134
rect -2614 593898 -2378 594134
rect -2934 584218 -2698 584454
rect -2614 584218 -2378 584454
rect -2934 583898 -2698 584134
rect -2614 583898 -2378 584134
rect -2934 574218 -2698 574454
rect -2614 574218 -2378 574454
rect -2934 573898 -2698 574134
rect -2614 573898 -2378 574134
rect -2934 564218 -2698 564454
rect -2614 564218 -2378 564454
rect -2934 563898 -2698 564134
rect -2614 563898 -2378 564134
rect -2934 554218 -2698 554454
rect -2614 554218 -2378 554454
rect -2934 553898 -2698 554134
rect -2614 553898 -2378 554134
rect -2934 544218 -2698 544454
rect -2614 544218 -2378 544454
rect -2934 543898 -2698 544134
rect -2614 543898 -2378 544134
rect -2934 534218 -2698 534454
rect -2614 534218 -2378 534454
rect -2934 533898 -2698 534134
rect -2614 533898 -2378 534134
rect -2934 524218 -2698 524454
rect -2614 524218 -2378 524454
rect -2934 523898 -2698 524134
rect -2614 523898 -2378 524134
rect -2934 514218 -2698 514454
rect -2614 514218 -2378 514454
rect -2934 513898 -2698 514134
rect -2614 513898 -2378 514134
rect -2934 504218 -2698 504454
rect -2614 504218 -2378 504454
rect -2934 503898 -2698 504134
rect -2614 503898 -2378 504134
rect -2934 494218 -2698 494454
rect -2614 494218 -2378 494454
rect -2934 493898 -2698 494134
rect -2614 493898 -2378 494134
rect -2934 484218 -2698 484454
rect -2614 484218 -2378 484454
rect -2934 483898 -2698 484134
rect -2614 483898 -2378 484134
rect -2934 474218 -2698 474454
rect -2614 474218 -2378 474454
rect -2934 473898 -2698 474134
rect -2614 473898 -2378 474134
rect -2934 464218 -2698 464454
rect -2614 464218 -2378 464454
rect -2934 463898 -2698 464134
rect -2614 463898 -2378 464134
rect -2934 454218 -2698 454454
rect -2614 454218 -2378 454454
rect -2934 453898 -2698 454134
rect -2614 453898 -2378 454134
rect -2934 444218 -2698 444454
rect -2614 444218 -2378 444454
rect -2934 443898 -2698 444134
rect -2614 443898 -2378 444134
rect -2934 434218 -2698 434454
rect -2614 434218 -2378 434454
rect -2934 433898 -2698 434134
rect -2614 433898 -2378 434134
rect -2934 424218 -2698 424454
rect -2614 424218 -2378 424454
rect -2934 423898 -2698 424134
rect -2614 423898 -2378 424134
rect -2934 414218 -2698 414454
rect -2614 414218 -2378 414454
rect -2934 413898 -2698 414134
rect -2614 413898 -2378 414134
rect -2934 404218 -2698 404454
rect -2614 404218 -2378 404454
rect -2934 403898 -2698 404134
rect -2614 403898 -2378 404134
rect -2934 394218 -2698 394454
rect -2614 394218 -2378 394454
rect -2934 393898 -2698 394134
rect -2614 393898 -2378 394134
rect -2934 384218 -2698 384454
rect -2614 384218 -2378 384454
rect -2934 383898 -2698 384134
rect -2614 383898 -2378 384134
rect -2934 374218 -2698 374454
rect -2614 374218 -2378 374454
rect -2934 373898 -2698 374134
rect -2614 373898 -2378 374134
rect -2934 364218 -2698 364454
rect -2614 364218 -2378 364454
rect -2934 363898 -2698 364134
rect -2614 363898 -2378 364134
rect -2934 354218 -2698 354454
rect -2614 354218 -2378 354454
rect -2934 353898 -2698 354134
rect -2614 353898 -2378 354134
rect -2934 344218 -2698 344454
rect -2614 344218 -2378 344454
rect -2934 343898 -2698 344134
rect -2614 343898 -2378 344134
rect -2934 334218 -2698 334454
rect -2614 334218 -2378 334454
rect -2934 333898 -2698 334134
rect -2614 333898 -2378 334134
rect -2934 324218 -2698 324454
rect -2614 324218 -2378 324454
rect -2934 323898 -2698 324134
rect -2614 323898 -2378 324134
rect -2934 314218 -2698 314454
rect -2614 314218 -2378 314454
rect -2934 313898 -2698 314134
rect -2614 313898 -2378 314134
rect -2934 304218 -2698 304454
rect -2614 304218 -2378 304454
rect -2934 303898 -2698 304134
rect -2614 303898 -2378 304134
rect -2934 294218 -2698 294454
rect -2614 294218 -2378 294454
rect -2934 293898 -2698 294134
rect -2614 293898 -2378 294134
rect -2934 284218 -2698 284454
rect -2614 284218 -2378 284454
rect -2934 283898 -2698 284134
rect -2614 283898 -2378 284134
rect -2934 274218 -2698 274454
rect -2614 274218 -2378 274454
rect -2934 273898 -2698 274134
rect -2614 273898 -2378 274134
rect -2934 264218 -2698 264454
rect -2614 264218 -2378 264454
rect -2934 263898 -2698 264134
rect -2614 263898 -2378 264134
rect -2934 254218 -2698 254454
rect -2614 254218 -2378 254454
rect -2934 253898 -2698 254134
rect -2614 253898 -2378 254134
rect -2934 244218 -2698 244454
rect -2614 244218 -2378 244454
rect -2934 243898 -2698 244134
rect -2614 243898 -2378 244134
rect -2934 234218 -2698 234454
rect -2614 234218 -2378 234454
rect -2934 233898 -2698 234134
rect -2614 233898 -2378 234134
rect -2934 224218 -2698 224454
rect -2614 224218 -2378 224454
rect -2934 223898 -2698 224134
rect -2614 223898 -2378 224134
rect -2934 214218 -2698 214454
rect -2614 214218 -2378 214454
rect -2934 213898 -2698 214134
rect -2614 213898 -2378 214134
rect -2934 204218 -2698 204454
rect -2614 204218 -2378 204454
rect -2934 203898 -2698 204134
rect -2614 203898 -2378 204134
rect -2934 194218 -2698 194454
rect -2614 194218 -2378 194454
rect -2934 193898 -2698 194134
rect -2614 193898 -2378 194134
rect -2934 184218 -2698 184454
rect -2614 184218 -2378 184454
rect -2934 183898 -2698 184134
rect -2614 183898 -2378 184134
rect -2934 174218 -2698 174454
rect -2614 174218 -2378 174454
rect -2934 173898 -2698 174134
rect -2614 173898 -2378 174134
rect -2934 164218 -2698 164454
rect -2614 164218 -2378 164454
rect -2934 163898 -2698 164134
rect -2614 163898 -2378 164134
rect -2934 154218 -2698 154454
rect -2614 154218 -2378 154454
rect -2934 153898 -2698 154134
rect -2614 153898 -2378 154134
rect -2934 144218 -2698 144454
rect -2614 144218 -2378 144454
rect -2934 143898 -2698 144134
rect -2614 143898 -2378 144134
rect -2934 134218 -2698 134454
rect -2614 134218 -2378 134454
rect -2934 133898 -2698 134134
rect -2614 133898 -2378 134134
rect -2934 124218 -2698 124454
rect -2614 124218 -2378 124454
rect -2934 123898 -2698 124134
rect -2614 123898 -2378 124134
rect -2934 114218 -2698 114454
rect -2614 114218 -2378 114454
rect -2934 113898 -2698 114134
rect -2614 113898 -2378 114134
rect -2934 104218 -2698 104454
rect -2614 104218 -2378 104454
rect -2934 103898 -2698 104134
rect -2614 103898 -2378 104134
rect -2934 94218 -2698 94454
rect -2614 94218 -2378 94454
rect -2934 93898 -2698 94134
rect -2614 93898 -2378 94134
rect -2934 84218 -2698 84454
rect -2614 84218 -2378 84454
rect -2934 83898 -2698 84134
rect -2614 83898 -2378 84134
rect -2934 74218 -2698 74454
rect -2614 74218 -2378 74454
rect -2934 73898 -2698 74134
rect -2614 73898 -2378 74134
rect -2934 64218 -2698 64454
rect -2614 64218 -2378 64454
rect -2934 63898 -2698 64134
rect -2614 63898 -2378 64134
rect -2934 54218 -2698 54454
rect -2614 54218 -2378 54454
rect -2934 53898 -2698 54134
rect -2614 53898 -2378 54134
rect -2934 44218 -2698 44454
rect -2614 44218 -2378 44454
rect -2934 43898 -2698 44134
rect -2614 43898 -2378 44134
rect -2934 34218 -2698 34454
rect -2614 34218 -2378 34454
rect -2934 33898 -2698 34134
rect -2614 33898 -2378 34134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect -1974 697938 -1738 698174
rect -1654 697938 -1418 698174
rect -1974 697618 -1738 697854
rect -1654 697618 -1418 697854
rect -1974 687938 -1738 688174
rect -1654 687938 -1418 688174
rect -1974 687618 -1738 687854
rect -1654 687618 -1418 687854
rect -1974 677938 -1738 678174
rect -1654 677938 -1418 678174
rect -1974 677618 -1738 677854
rect -1654 677618 -1418 677854
rect -1974 667938 -1738 668174
rect -1654 667938 -1418 668174
rect -1974 667618 -1738 667854
rect -1654 667618 -1418 667854
rect -1974 657938 -1738 658174
rect -1654 657938 -1418 658174
rect -1974 657618 -1738 657854
rect -1654 657618 -1418 657854
rect -1974 647938 -1738 648174
rect -1654 647938 -1418 648174
rect -1974 647618 -1738 647854
rect -1654 647618 -1418 647854
rect -1974 637938 -1738 638174
rect -1654 637938 -1418 638174
rect -1974 637618 -1738 637854
rect -1654 637618 -1418 637854
rect -1974 627938 -1738 628174
rect -1654 627938 -1418 628174
rect -1974 627618 -1738 627854
rect -1654 627618 -1418 627854
rect -1974 617938 -1738 618174
rect -1654 617938 -1418 618174
rect -1974 617618 -1738 617854
rect -1654 617618 -1418 617854
rect -1974 607938 -1738 608174
rect -1654 607938 -1418 608174
rect -1974 607618 -1738 607854
rect -1654 607618 -1418 607854
rect -1974 597938 -1738 598174
rect -1654 597938 -1418 598174
rect -1974 597618 -1738 597854
rect -1654 597618 -1418 597854
rect -1974 587938 -1738 588174
rect -1654 587938 -1418 588174
rect -1974 587618 -1738 587854
rect -1654 587618 -1418 587854
rect -1974 577938 -1738 578174
rect -1654 577938 -1418 578174
rect -1974 577618 -1738 577854
rect -1654 577618 -1418 577854
rect -1974 567938 -1738 568174
rect -1654 567938 -1418 568174
rect -1974 567618 -1738 567854
rect -1654 567618 -1418 567854
rect -1974 557938 -1738 558174
rect -1654 557938 -1418 558174
rect -1974 557618 -1738 557854
rect -1654 557618 -1418 557854
rect -1974 547938 -1738 548174
rect -1654 547938 -1418 548174
rect -1974 547618 -1738 547854
rect -1654 547618 -1418 547854
rect -1974 537938 -1738 538174
rect -1654 537938 -1418 538174
rect -1974 537618 -1738 537854
rect -1654 537618 -1418 537854
rect -1974 527938 -1738 528174
rect -1654 527938 -1418 528174
rect -1974 527618 -1738 527854
rect -1654 527618 -1418 527854
rect -1974 517938 -1738 518174
rect -1654 517938 -1418 518174
rect -1974 517618 -1738 517854
rect -1654 517618 -1418 517854
rect -1974 507938 -1738 508174
rect -1654 507938 -1418 508174
rect -1974 507618 -1738 507854
rect -1654 507618 -1418 507854
rect -1974 497938 -1738 498174
rect -1654 497938 -1418 498174
rect -1974 497618 -1738 497854
rect -1654 497618 -1418 497854
rect -1974 487938 -1738 488174
rect -1654 487938 -1418 488174
rect -1974 487618 -1738 487854
rect -1654 487618 -1418 487854
rect -1974 477938 -1738 478174
rect -1654 477938 -1418 478174
rect -1974 477618 -1738 477854
rect -1654 477618 -1418 477854
rect -1974 467938 -1738 468174
rect -1654 467938 -1418 468174
rect -1974 467618 -1738 467854
rect -1654 467618 -1418 467854
rect -1974 457938 -1738 458174
rect -1654 457938 -1418 458174
rect -1974 457618 -1738 457854
rect -1654 457618 -1418 457854
rect -1974 447938 -1738 448174
rect -1654 447938 -1418 448174
rect -1974 447618 -1738 447854
rect -1654 447618 -1418 447854
rect -1974 437938 -1738 438174
rect -1654 437938 -1418 438174
rect -1974 437618 -1738 437854
rect -1654 437618 -1418 437854
rect -1974 427938 -1738 428174
rect -1654 427938 -1418 428174
rect -1974 427618 -1738 427854
rect -1654 427618 -1418 427854
rect -1974 417938 -1738 418174
rect -1654 417938 -1418 418174
rect -1974 417618 -1738 417854
rect -1654 417618 -1418 417854
rect -1974 407938 -1738 408174
rect -1654 407938 -1418 408174
rect -1974 407618 -1738 407854
rect -1654 407618 -1418 407854
rect -1974 397938 -1738 398174
rect -1654 397938 -1418 398174
rect -1974 397618 -1738 397854
rect -1654 397618 -1418 397854
rect -1974 387938 -1738 388174
rect -1654 387938 -1418 388174
rect -1974 387618 -1738 387854
rect -1654 387618 -1418 387854
rect -1974 377938 -1738 378174
rect -1654 377938 -1418 378174
rect -1974 377618 -1738 377854
rect -1654 377618 -1418 377854
rect -1974 367938 -1738 368174
rect -1654 367938 -1418 368174
rect -1974 367618 -1738 367854
rect -1654 367618 -1418 367854
rect -1974 357938 -1738 358174
rect -1654 357938 -1418 358174
rect -1974 357618 -1738 357854
rect -1654 357618 -1418 357854
rect -1974 347938 -1738 348174
rect -1654 347938 -1418 348174
rect -1974 347618 -1738 347854
rect -1654 347618 -1418 347854
rect -1974 337938 -1738 338174
rect -1654 337938 -1418 338174
rect -1974 337618 -1738 337854
rect -1654 337618 -1418 337854
rect -1974 327938 -1738 328174
rect -1654 327938 -1418 328174
rect -1974 327618 -1738 327854
rect -1654 327618 -1418 327854
rect -1974 317938 -1738 318174
rect -1654 317938 -1418 318174
rect -1974 317618 -1738 317854
rect -1654 317618 -1418 317854
rect -1974 307938 -1738 308174
rect -1654 307938 -1418 308174
rect -1974 307618 -1738 307854
rect -1654 307618 -1418 307854
rect -1974 297938 -1738 298174
rect -1654 297938 -1418 298174
rect -1974 297618 -1738 297854
rect -1654 297618 -1418 297854
rect -1974 287938 -1738 288174
rect -1654 287938 -1418 288174
rect -1974 287618 -1738 287854
rect -1654 287618 -1418 287854
rect -1974 277938 -1738 278174
rect -1654 277938 -1418 278174
rect -1974 277618 -1738 277854
rect -1654 277618 -1418 277854
rect -1974 267938 -1738 268174
rect -1654 267938 -1418 268174
rect -1974 267618 -1738 267854
rect -1654 267618 -1418 267854
rect -1974 257938 -1738 258174
rect -1654 257938 -1418 258174
rect -1974 257618 -1738 257854
rect -1654 257618 -1418 257854
rect -1974 247938 -1738 248174
rect -1654 247938 -1418 248174
rect -1974 247618 -1738 247854
rect -1654 247618 -1418 247854
rect -1974 237938 -1738 238174
rect -1654 237938 -1418 238174
rect -1974 237618 -1738 237854
rect -1654 237618 -1418 237854
rect -1974 227938 -1738 228174
rect -1654 227938 -1418 228174
rect -1974 227618 -1738 227854
rect -1654 227618 -1418 227854
rect -1974 217938 -1738 218174
rect -1654 217938 -1418 218174
rect -1974 217618 -1738 217854
rect -1654 217618 -1418 217854
rect -1974 207938 -1738 208174
rect -1654 207938 -1418 208174
rect -1974 207618 -1738 207854
rect -1654 207618 -1418 207854
rect -1974 197938 -1738 198174
rect -1654 197938 -1418 198174
rect -1974 197618 -1738 197854
rect -1654 197618 -1418 197854
rect -1974 187938 -1738 188174
rect -1654 187938 -1418 188174
rect -1974 187618 -1738 187854
rect -1654 187618 -1418 187854
rect -1974 177938 -1738 178174
rect -1654 177938 -1418 178174
rect -1974 177618 -1738 177854
rect -1654 177618 -1418 177854
rect -1974 167938 -1738 168174
rect -1654 167938 -1418 168174
rect -1974 167618 -1738 167854
rect -1654 167618 -1418 167854
rect -1974 157938 -1738 158174
rect -1654 157938 -1418 158174
rect -1974 157618 -1738 157854
rect -1654 157618 -1418 157854
rect -1974 147938 -1738 148174
rect -1654 147938 -1418 148174
rect -1974 147618 -1738 147854
rect -1654 147618 -1418 147854
rect -1974 137938 -1738 138174
rect -1654 137938 -1418 138174
rect -1974 137618 -1738 137854
rect -1654 137618 -1418 137854
rect -1974 127938 -1738 128174
rect -1654 127938 -1418 128174
rect -1974 127618 -1738 127854
rect -1654 127618 -1418 127854
rect -1974 117938 -1738 118174
rect -1654 117938 -1418 118174
rect -1974 117618 -1738 117854
rect -1654 117618 -1418 117854
rect -1974 107938 -1738 108174
rect -1654 107938 -1418 108174
rect -1974 107618 -1738 107854
rect -1654 107618 -1418 107854
rect -1974 97938 -1738 98174
rect -1654 97938 -1418 98174
rect -1974 97618 -1738 97854
rect -1654 97618 -1418 97854
rect -1974 87938 -1738 88174
rect -1654 87938 -1418 88174
rect -1974 87618 -1738 87854
rect -1654 87618 -1418 87854
rect -1974 77938 -1738 78174
rect -1654 77938 -1418 78174
rect -1974 77618 -1738 77854
rect -1654 77618 -1418 77854
rect -1974 67938 -1738 68174
rect -1654 67938 -1418 68174
rect -1974 67618 -1738 67854
rect -1654 67618 -1418 67854
rect -1974 57938 -1738 58174
rect -1654 57938 -1418 58174
rect -1974 57618 -1738 57854
rect -1654 57618 -1418 57854
rect -1974 47938 -1738 48174
rect -1654 47938 -1418 48174
rect -1974 47618 -1738 47854
rect -1654 47618 -1418 47854
rect -1974 37938 -1738 38174
rect -1654 37938 -1418 38174
rect -1974 37618 -1738 37854
rect -1654 37618 -1418 37854
rect 14107 207938 14343 208174
rect 14107 207618 14343 207854
rect 21949 207938 22185 208174
rect 21949 207618 22185 207854
rect 29791 207938 30027 208174
rect 29791 207618 30027 207854
rect 37633 207938 37869 208174
rect 37633 207618 37869 207854
rect 48239 207938 48475 208174
rect 48239 207618 48475 207854
rect 56081 207938 56317 208174
rect 56081 207618 56317 207854
rect 63923 207938 64159 208174
rect 63923 207618 64159 207854
rect 71765 207938 72001 208174
rect 71765 207618 72001 207854
rect 82371 207938 82607 208174
rect 82371 207618 82607 207854
rect 90213 207938 90449 208174
rect 90213 207618 90449 207854
rect 98055 207938 98291 208174
rect 98055 207618 98291 207854
rect 105897 207938 106133 208174
rect 105897 207618 106133 207854
rect 116503 207938 116739 208174
rect 116503 207618 116739 207854
rect 124345 207938 124581 208174
rect 124345 207618 124581 207854
rect 132187 207938 132423 208174
rect 132187 207618 132423 207854
rect 140029 207938 140265 208174
rect 140029 207618 140265 207854
rect 150635 207938 150871 208174
rect 150635 207618 150871 207854
rect 158477 207938 158713 208174
rect 158477 207618 158713 207854
rect 166319 207938 166555 208174
rect 166319 207618 166555 207854
rect 174161 207938 174397 208174
rect 174161 207618 174397 207854
rect 184767 207938 185003 208174
rect 184767 207618 185003 207854
rect 192609 207938 192845 208174
rect 192609 207618 192845 207854
rect 200451 207938 200687 208174
rect 200451 207618 200687 207854
rect 208293 207938 208529 208174
rect 208293 207618 208529 207854
rect 218899 207938 219135 208174
rect 218899 207618 219135 207854
rect 226741 207938 226977 208174
rect 226741 207618 226977 207854
rect 234583 207938 234819 208174
rect 234583 207618 234819 207854
rect 242425 207938 242661 208174
rect 242425 207618 242661 207854
rect 253031 207938 253267 208174
rect 253031 207618 253267 207854
rect 260873 207938 261109 208174
rect 260873 207618 261109 207854
rect 268715 207938 268951 208174
rect 268715 207618 268951 207854
rect 276557 207938 276793 208174
rect 276557 207618 276793 207854
rect 18028 204218 18264 204454
rect 18028 203898 18264 204134
rect 25870 204218 26106 204454
rect 25870 203898 26106 204134
rect 33712 204218 33948 204454
rect 33712 203898 33948 204134
rect 41554 204218 41790 204454
rect 41554 203898 41790 204134
rect 52160 204218 52396 204454
rect 52160 203898 52396 204134
rect 60002 204218 60238 204454
rect 60002 203898 60238 204134
rect 67844 204218 68080 204454
rect 67844 203898 68080 204134
rect 75686 204218 75922 204454
rect 75686 203898 75922 204134
rect 86292 204218 86528 204454
rect 86292 203898 86528 204134
rect 94134 204218 94370 204454
rect 94134 203898 94370 204134
rect 101976 204218 102212 204454
rect 101976 203898 102212 204134
rect 109818 204218 110054 204454
rect 109818 203898 110054 204134
rect 120424 204218 120660 204454
rect 120424 203898 120660 204134
rect 128266 204218 128502 204454
rect 128266 203898 128502 204134
rect 136108 204218 136344 204454
rect 136108 203898 136344 204134
rect 143950 204218 144186 204454
rect 143950 203898 144186 204134
rect 154556 204218 154792 204454
rect 154556 203898 154792 204134
rect 162398 204218 162634 204454
rect 162398 203898 162634 204134
rect 170240 204218 170476 204454
rect 170240 203898 170476 204134
rect 178082 204218 178318 204454
rect 178082 203898 178318 204134
rect 188688 204218 188924 204454
rect 188688 203898 188924 204134
rect 196530 204218 196766 204454
rect 196530 203898 196766 204134
rect 204372 204218 204608 204454
rect 204372 203898 204608 204134
rect 212214 204218 212450 204454
rect 212214 203898 212450 204134
rect 222820 204218 223056 204454
rect 222820 203898 223056 204134
rect 230662 204218 230898 204454
rect 230662 203898 230898 204134
rect 238504 204218 238740 204454
rect 238504 203898 238740 204134
rect 246346 204218 246582 204454
rect 246346 203898 246582 204134
rect 256952 204218 257188 204454
rect 256952 203898 257188 204134
rect 264794 204218 265030 204454
rect 264794 203898 265030 204134
rect 272636 204218 272872 204454
rect 272636 203898 272872 204134
rect 280478 204218 280714 204454
rect 280478 203898 280714 204134
rect 14107 197938 14343 198174
rect 14107 197618 14343 197854
rect 21949 197938 22185 198174
rect 21949 197618 22185 197854
rect 29791 197938 30027 198174
rect 29791 197618 30027 197854
rect 37633 197938 37869 198174
rect 37633 197618 37869 197854
rect 48239 197938 48475 198174
rect 48239 197618 48475 197854
rect 56081 197938 56317 198174
rect 56081 197618 56317 197854
rect 63923 197938 64159 198174
rect 63923 197618 64159 197854
rect 71765 197938 72001 198174
rect 71765 197618 72001 197854
rect 82371 197938 82607 198174
rect 82371 197618 82607 197854
rect 90213 197938 90449 198174
rect 90213 197618 90449 197854
rect 98055 197938 98291 198174
rect 98055 197618 98291 197854
rect 105897 197938 106133 198174
rect 105897 197618 106133 197854
rect 116503 197938 116739 198174
rect 116503 197618 116739 197854
rect 124345 197938 124581 198174
rect 124345 197618 124581 197854
rect 132187 197938 132423 198174
rect 132187 197618 132423 197854
rect 140029 197938 140265 198174
rect 140029 197618 140265 197854
rect 150635 197938 150871 198174
rect 150635 197618 150871 197854
rect 158477 197938 158713 198174
rect 158477 197618 158713 197854
rect 166319 197938 166555 198174
rect 166319 197618 166555 197854
rect 174161 197938 174397 198174
rect 174161 197618 174397 197854
rect 184767 197938 185003 198174
rect 184767 197618 185003 197854
rect 192609 197938 192845 198174
rect 192609 197618 192845 197854
rect 200451 197938 200687 198174
rect 200451 197618 200687 197854
rect 208293 197938 208529 198174
rect 208293 197618 208529 197854
rect 218899 197938 219135 198174
rect 218899 197618 219135 197854
rect 226741 197938 226977 198174
rect 226741 197618 226977 197854
rect 234583 197938 234819 198174
rect 234583 197618 234819 197854
rect 242425 197938 242661 198174
rect 242425 197618 242661 197854
rect 253031 197938 253267 198174
rect 253031 197618 253267 197854
rect 260873 197938 261109 198174
rect 260873 197618 261109 197854
rect 268715 197938 268951 198174
rect 268715 197618 268951 197854
rect 276557 197938 276793 198174
rect 276557 197618 276793 197854
rect 18028 194218 18264 194454
rect 18028 193898 18264 194134
rect 25870 194218 26106 194454
rect 25870 193898 26106 194134
rect 33712 194218 33948 194454
rect 33712 193898 33948 194134
rect 41554 194218 41790 194454
rect 41554 193898 41790 194134
rect 52160 194218 52396 194454
rect 52160 193898 52396 194134
rect 60002 194218 60238 194454
rect 60002 193898 60238 194134
rect 67844 194218 68080 194454
rect 67844 193898 68080 194134
rect 75686 194218 75922 194454
rect 75686 193898 75922 194134
rect 86292 194218 86528 194454
rect 86292 193898 86528 194134
rect 94134 194218 94370 194454
rect 94134 193898 94370 194134
rect 101976 194218 102212 194454
rect 101976 193898 102212 194134
rect 109818 194218 110054 194454
rect 109818 193898 110054 194134
rect 120424 194218 120660 194454
rect 120424 193898 120660 194134
rect 128266 194218 128502 194454
rect 128266 193898 128502 194134
rect 136108 194218 136344 194454
rect 136108 193898 136344 194134
rect 143950 194218 144186 194454
rect 143950 193898 144186 194134
rect 154556 194218 154792 194454
rect 154556 193898 154792 194134
rect 162398 194218 162634 194454
rect 162398 193898 162634 194134
rect 170240 194218 170476 194454
rect 170240 193898 170476 194134
rect 178082 194218 178318 194454
rect 178082 193898 178318 194134
rect 188688 194218 188924 194454
rect 188688 193898 188924 194134
rect 196530 194218 196766 194454
rect 196530 193898 196766 194134
rect 204372 194218 204608 194454
rect 204372 193898 204608 194134
rect 212214 194218 212450 194454
rect 212214 193898 212450 194134
rect 222820 194218 223056 194454
rect 222820 193898 223056 194134
rect 230662 194218 230898 194454
rect 230662 193898 230898 194134
rect 238504 194218 238740 194454
rect 238504 193898 238740 194134
rect 246346 194218 246582 194454
rect 246346 193898 246582 194134
rect 256952 194218 257188 194454
rect 256952 193898 257188 194134
rect 264794 194218 265030 194454
rect 264794 193898 265030 194134
rect 272636 194218 272872 194454
rect 272636 193898 272872 194134
rect 280478 194218 280714 194454
rect 280478 193898 280714 194134
rect 43984 187938 44220 188174
rect 43984 187618 44220 187854
rect 111581 187938 111817 188174
rect 111581 187618 111817 187854
rect 179178 187938 179414 188174
rect 179178 187618 179414 187854
rect 246775 187938 247011 188174
rect 246775 187618 247011 187854
rect 77782 184218 78018 184454
rect 77782 183898 78018 184134
rect 145379 184218 145615 184454
rect 145379 183898 145615 184134
rect 212976 184218 213212 184454
rect 212976 183898 213212 184134
rect 280573 184218 280809 184454
rect 280573 183898 280809 184134
rect 585342 697938 585578 698174
rect 585662 697938 585898 698174
rect 585342 697618 585578 697854
rect 585662 697618 585898 697854
rect 585342 687938 585578 688174
rect 585662 687938 585898 688174
rect 585342 687618 585578 687854
rect 585662 687618 585898 687854
rect 585342 677938 585578 678174
rect 585662 677938 585898 678174
rect 585342 677618 585578 677854
rect 585662 677618 585898 677854
rect 14107 177643 14343 177879
rect 21949 177643 22185 177879
rect 29791 177643 30027 177879
rect 37633 177643 37869 177879
rect 18028 174218 18264 174454
rect 18028 173898 18264 174134
rect 25870 174218 26106 174454
rect 25870 173898 26106 174134
rect 33712 174218 33948 174454
rect 33712 173898 33948 174134
rect 41554 174218 41790 174454
rect 41554 173898 41790 174134
rect 14107 167938 14343 168174
rect 14107 167618 14343 167854
rect 21949 167938 22185 168174
rect 21949 167618 22185 167854
rect 29791 167938 30027 168174
rect 29791 167618 30027 167854
rect 37633 167938 37869 168174
rect 37633 167618 37869 167854
rect 18028 164218 18264 164454
rect 18028 163898 18264 164134
rect 25870 164218 26106 164454
rect 25870 163898 26106 164134
rect 33712 164218 33948 164454
rect 33712 163898 33948 164134
rect 41554 164218 41790 164454
rect 41554 163898 41790 164134
rect 48239 177643 48475 177879
rect 56081 177643 56317 177879
rect 63923 177643 64159 177879
rect 71765 177643 72001 177879
rect 82371 177643 82607 177879
rect 90213 177643 90449 177879
rect 98055 177643 98291 177879
rect 105897 177643 106133 177879
rect 52160 174218 52396 174454
rect 52160 173898 52396 174134
rect 60002 174218 60238 174454
rect 60002 173898 60238 174134
rect 67844 174218 68080 174454
rect 67844 173898 68080 174134
rect 75686 174218 75922 174454
rect 75686 173898 75922 174134
rect 86292 174218 86528 174454
rect 86292 173898 86528 174134
rect 94134 174218 94370 174454
rect 94134 173898 94370 174134
rect 101976 174218 102212 174454
rect 101976 173898 102212 174134
rect 109818 174218 110054 174454
rect 109818 173898 110054 174134
rect 48239 167938 48475 168174
rect 48239 167618 48475 167854
rect 56081 167938 56317 168174
rect 56081 167618 56317 167854
rect 63923 167938 64159 168174
rect 63923 167618 64159 167854
rect 71765 167938 72001 168174
rect 71765 167618 72001 167854
rect 82371 167938 82607 168174
rect 82371 167618 82607 167854
rect 90213 167938 90449 168174
rect 90213 167618 90449 167854
rect 98055 167938 98291 168174
rect 98055 167618 98291 167854
rect 105897 167938 106133 168174
rect 105897 167618 106133 167854
rect 52160 164218 52396 164454
rect 52160 163898 52396 164134
rect 60002 164218 60238 164454
rect 60002 163898 60238 164134
rect 67844 164218 68080 164454
rect 67844 163898 68080 164134
rect 75686 164218 75922 164454
rect 75686 163898 75922 164134
rect 86292 164218 86528 164454
rect 86292 163898 86528 164134
rect 94134 164218 94370 164454
rect 94134 163898 94370 164134
rect 101976 164218 102212 164454
rect 101976 163898 102212 164134
rect 109818 164218 110054 164454
rect 109818 163898 110054 164134
rect 116503 177643 116739 177879
rect 124345 177643 124581 177879
rect 132187 177643 132423 177879
rect 140029 177643 140265 177879
rect 150635 177643 150871 177879
rect 158477 177643 158713 177879
rect 166319 177643 166555 177879
rect 174161 177643 174397 177879
rect 184767 177643 185003 177879
rect 192609 177643 192845 177879
rect 200451 177643 200687 177879
rect 208293 177643 208529 177879
rect 218899 177643 219135 177879
rect 226741 177643 226977 177879
rect 234583 177643 234819 177879
rect 242425 177643 242661 177879
rect 120424 174218 120660 174454
rect 120424 173898 120660 174134
rect 128266 174218 128502 174454
rect 128266 173898 128502 174134
rect 136108 174218 136344 174454
rect 136108 173898 136344 174134
rect 143950 174218 144186 174454
rect 143950 173898 144186 174134
rect 154556 174218 154792 174454
rect 154556 173898 154792 174134
rect 162398 174218 162634 174454
rect 162398 173898 162634 174134
rect 170240 174218 170476 174454
rect 170240 173898 170476 174134
rect 178082 174218 178318 174454
rect 178082 173898 178318 174134
rect 188688 174218 188924 174454
rect 188688 173898 188924 174134
rect 196530 174218 196766 174454
rect 196530 173898 196766 174134
rect 204372 174218 204608 174454
rect 204372 173898 204608 174134
rect 212214 174218 212450 174454
rect 212214 173898 212450 174134
rect 222820 174218 223056 174454
rect 222820 173898 223056 174134
rect 230662 174218 230898 174454
rect 230662 173898 230898 174134
rect 238504 174218 238740 174454
rect 238504 173898 238740 174134
rect 246346 174218 246582 174454
rect 246346 173898 246582 174134
rect 116503 167938 116739 168174
rect 116503 167618 116739 167854
rect 124345 167938 124581 168174
rect 124345 167618 124581 167854
rect 132187 167938 132423 168174
rect 132187 167618 132423 167854
rect 140029 167938 140265 168174
rect 140029 167618 140265 167854
rect 150635 167938 150871 168174
rect 150635 167618 150871 167854
rect 158477 167938 158713 168174
rect 158477 167618 158713 167854
rect 166319 167938 166555 168174
rect 166319 167618 166555 167854
rect 174161 167938 174397 168174
rect 174161 167618 174397 167854
rect 184767 167938 185003 168174
rect 184767 167618 185003 167854
rect 192609 167938 192845 168174
rect 192609 167618 192845 167854
rect 200451 167938 200687 168174
rect 200451 167618 200687 167854
rect 208293 167938 208529 168174
rect 208293 167618 208529 167854
rect 218899 167938 219135 168174
rect 218899 167618 219135 167854
rect 226741 167938 226977 168174
rect 226741 167618 226977 167854
rect 234583 167938 234819 168174
rect 234583 167618 234819 167854
rect 242425 167938 242661 168174
rect 242425 167618 242661 167854
rect 120424 164218 120660 164454
rect 120424 163898 120660 164134
rect 128266 164218 128502 164454
rect 128266 163898 128502 164134
rect 136108 164218 136344 164454
rect 136108 163898 136344 164134
rect 143950 164218 144186 164454
rect 143950 163898 144186 164134
rect 154556 164218 154792 164454
rect 154556 163898 154792 164134
rect 162398 164218 162634 164454
rect 162398 163898 162634 164134
rect 170240 164218 170476 164454
rect 170240 163898 170476 164134
rect 178082 164218 178318 164454
rect 178082 163898 178318 164134
rect 188688 164218 188924 164454
rect 188688 163898 188924 164134
rect 196530 164218 196766 164454
rect 196530 163898 196766 164134
rect 204372 164218 204608 164454
rect 204372 163898 204608 164134
rect 212214 164218 212450 164454
rect 212214 163898 212450 164134
rect 222820 164218 223056 164454
rect 222820 163898 223056 164134
rect 230662 164218 230898 164454
rect 230662 163898 230898 164134
rect 238504 164218 238740 164454
rect 238504 163898 238740 164134
rect 246346 164218 246582 164454
rect 246346 163898 246582 164134
rect 253031 177643 253267 177879
rect 260873 177643 261109 177879
rect 268715 177643 268951 177879
rect 276557 177643 276793 177879
rect 256952 174218 257188 174454
rect 256952 173898 257188 174134
rect 264794 174218 265030 174454
rect 264794 173898 265030 174134
rect 272636 174218 272872 174454
rect 272636 173898 272872 174134
rect 280478 174218 280714 174454
rect 280478 173898 280714 174134
rect 253031 167938 253267 168174
rect 253031 167618 253267 167854
rect 260873 167938 261109 168174
rect 260873 167618 261109 167854
rect 268715 167938 268951 168174
rect 268715 167618 268951 167854
rect 276557 167938 276793 168174
rect 276557 167618 276793 167854
rect 256952 164218 257188 164454
rect 256952 163898 257188 164134
rect 264794 164218 265030 164454
rect 264794 163898 265030 164134
rect 272636 164218 272872 164454
rect 272636 163898 272872 164134
rect 280478 164218 280714 164454
rect 280478 163898 280714 164134
rect 307407 207938 307643 208174
rect 307407 207618 307643 207854
rect 315249 207938 315485 208174
rect 315249 207618 315485 207854
rect 323091 207938 323327 208174
rect 323091 207618 323327 207854
rect 330933 207938 331169 208174
rect 330933 207618 331169 207854
rect 341539 207938 341775 208174
rect 341539 207618 341775 207854
rect 349381 207938 349617 208174
rect 349381 207618 349617 207854
rect 357223 207938 357459 208174
rect 357223 207618 357459 207854
rect 365065 207938 365301 208174
rect 365065 207618 365301 207854
rect 375671 207938 375907 208174
rect 375671 207618 375907 207854
rect 383513 207938 383749 208174
rect 383513 207618 383749 207854
rect 391355 207938 391591 208174
rect 391355 207618 391591 207854
rect 399197 207938 399433 208174
rect 399197 207618 399433 207854
rect 409803 207938 410039 208174
rect 409803 207618 410039 207854
rect 417645 207938 417881 208174
rect 417645 207618 417881 207854
rect 425487 207938 425723 208174
rect 425487 207618 425723 207854
rect 433329 207938 433565 208174
rect 433329 207618 433565 207854
rect 443935 207938 444171 208174
rect 443935 207618 444171 207854
rect 451777 207938 452013 208174
rect 451777 207618 452013 207854
rect 459619 207938 459855 208174
rect 459619 207618 459855 207854
rect 467461 207938 467697 208174
rect 467461 207618 467697 207854
rect 478067 207938 478303 208174
rect 478067 207618 478303 207854
rect 485909 207938 486145 208174
rect 485909 207618 486145 207854
rect 493751 207938 493987 208174
rect 493751 207618 493987 207854
rect 501593 207938 501829 208174
rect 501593 207618 501829 207854
rect 512199 207938 512435 208174
rect 512199 207618 512435 207854
rect 520041 207938 520277 208174
rect 520041 207618 520277 207854
rect 527883 207938 528119 208174
rect 527883 207618 528119 207854
rect 535725 207938 535961 208174
rect 535725 207618 535961 207854
rect 546331 207938 546567 208174
rect 546331 207618 546567 207854
rect 554173 207938 554409 208174
rect 554173 207618 554409 207854
rect 562015 207938 562251 208174
rect 562015 207618 562251 207854
rect 569857 207938 570093 208174
rect 569857 207618 570093 207854
rect 303486 204218 303722 204454
rect 303486 203898 303722 204134
rect 311328 204218 311564 204454
rect 311328 203898 311564 204134
rect 319170 204218 319406 204454
rect 319170 203898 319406 204134
rect 327012 204218 327248 204454
rect 327012 203898 327248 204134
rect 337618 204218 337854 204454
rect 337618 203898 337854 204134
rect 345460 204218 345696 204454
rect 345460 203898 345696 204134
rect 353302 204218 353538 204454
rect 353302 203898 353538 204134
rect 361144 204218 361380 204454
rect 361144 203898 361380 204134
rect 371750 204218 371986 204454
rect 371750 203898 371986 204134
rect 379592 204218 379828 204454
rect 379592 203898 379828 204134
rect 387434 204218 387670 204454
rect 387434 203898 387670 204134
rect 395276 204218 395512 204454
rect 395276 203898 395512 204134
rect 405882 204218 406118 204454
rect 405882 203898 406118 204134
rect 413724 204218 413960 204454
rect 413724 203898 413960 204134
rect 421566 204218 421802 204454
rect 421566 203898 421802 204134
rect 429408 204218 429644 204454
rect 429408 203898 429644 204134
rect 440014 204218 440250 204454
rect 440014 203898 440250 204134
rect 447856 204218 448092 204454
rect 447856 203898 448092 204134
rect 455698 204218 455934 204454
rect 455698 203898 455934 204134
rect 463540 204218 463776 204454
rect 463540 203898 463776 204134
rect 474146 204218 474382 204454
rect 474146 203898 474382 204134
rect 481988 204218 482224 204454
rect 481988 203898 482224 204134
rect 489830 204218 490066 204454
rect 489830 203898 490066 204134
rect 497672 204218 497908 204454
rect 497672 203898 497908 204134
rect 508278 204218 508514 204454
rect 508278 203898 508514 204134
rect 516120 204218 516356 204454
rect 516120 203898 516356 204134
rect 523962 204218 524198 204454
rect 523962 203898 524198 204134
rect 531804 204218 532040 204454
rect 531804 203898 532040 204134
rect 542410 204218 542646 204454
rect 542410 203898 542646 204134
rect 550252 204218 550488 204454
rect 550252 203898 550488 204134
rect 558094 204218 558330 204454
rect 558094 203898 558330 204134
rect 565936 204218 566172 204454
rect 565936 203898 566172 204134
rect 307407 197938 307643 198174
rect 307407 197618 307643 197854
rect 315249 197938 315485 198174
rect 315249 197618 315485 197854
rect 323091 197938 323327 198174
rect 323091 197618 323327 197854
rect 330933 197938 331169 198174
rect 330933 197618 331169 197854
rect 341539 197938 341775 198174
rect 341539 197618 341775 197854
rect 349381 197938 349617 198174
rect 349381 197618 349617 197854
rect 357223 197938 357459 198174
rect 357223 197618 357459 197854
rect 365065 197938 365301 198174
rect 365065 197618 365301 197854
rect 375671 197938 375907 198174
rect 375671 197618 375907 197854
rect 383513 197938 383749 198174
rect 383513 197618 383749 197854
rect 391355 197938 391591 198174
rect 391355 197618 391591 197854
rect 399197 197938 399433 198174
rect 399197 197618 399433 197854
rect 409803 197938 410039 198174
rect 409803 197618 410039 197854
rect 417645 197938 417881 198174
rect 417645 197618 417881 197854
rect 425487 197938 425723 198174
rect 425487 197618 425723 197854
rect 433329 197938 433565 198174
rect 433329 197618 433565 197854
rect 443935 197938 444171 198174
rect 443935 197618 444171 197854
rect 451777 197938 452013 198174
rect 451777 197618 452013 197854
rect 459619 197938 459855 198174
rect 459619 197618 459855 197854
rect 467461 197938 467697 198174
rect 467461 197618 467697 197854
rect 478067 197938 478303 198174
rect 478067 197618 478303 197854
rect 485909 197938 486145 198174
rect 485909 197618 486145 197854
rect 493751 197938 493987 198174
rect 493751 197618 493987 197854
rect 501593 197938 501829 198174
rect 501593 197618 501829 197854
rect 512199 197938 512435 198174
rect 512199 197618 512435 197854
rect 520041 197938 520277 198174
rect 520041 197618 520277 197854
rect 527883 197938 528119 198174
rect 527883 197618 528119 197854
rect 535725 197938 535961 198174
rect 535725 197618 535961 197854
rect 546331 197938 546567 198174
rect 546331 197618 546567 197854
rect 554173 197938 554409 198174
rect 554173 197618 554409 197854
rect 562015 197938 562251 198174
rect 562015 197618 562251 197854
rect 569857 197938 570093 198174
rect 569857 197618 570093 197854
rect 303486 194218 303722 194454
rect 303486 193898 303722 194134
rect 311328 194218 311564 194454
rect 311328 193898 311564 194134
rect 319170 194218 319406 194454
rect 319170 193898 319406 194134
rect 327012 194218 327248 194454
rect 327012 193898 327248 194134
rect 337618 194218 337854 194454
rect 337618 193898 337854 194134
rect 345460 194218 345696 194454
rect 345460 193898 345696 194134
rect 353302 194218 353538 194454
rect 353302 193898 353538 194134
rect 361144 194218 361380 194454
rect 361144 193898 361380 194134
rect 371750 194218 371986 194454
rect 371750 193898 371986 194134
rect 379592 194218 379828 194454
rect 379592 193898 379828 194134
rect 387434 194218 387670 194454
rect 387434 193898 387670 194134
rect 395276 194218 395512 194454
rect 395276 193898 395512 194134
rect 405882 194218 406118 194454
rect 405882 193898 406118 194134
rect 413724 194218 413960 194454
rect 413724 193898 413960 194134
rect 421566 194218 421802 194454
rect 421566 193898 421802 194134
rect 429408 194218 429644 194454
rect 429408 193898 429644 194134
rect 440014 194218 440250 194454
rect 440014 193898 440250 194134
rect 447856 194218 448092 194454
rect 447856 193898 448092 194134
rect 455698 194218 455934 194454
rect 455698 193898 455934 194134
rect 463540 194218 463776 194454
rect 463540 193898 463776 194134
rect 474146 194218 474382 194454
rect 474146 193898 474382 194134
rect 481988 194218 482224 194454
rect 481988 193898 482224 194134
rect 489830 194218 490066 194454
rect 489830 193898 490066 194134
rect 497672 194218 497908 194454
rect 497672 193898 497908 194134
rect 508278 194218 508514 194454
rect 508278 193898 508514 194134
rect 516120 194218 516356 194454
rect 516120 193898 516356 194134
rect 523962 194218 524198 194454
rect 523962 193898 524198 194134
rect 531804 194218 532040 194454
rect 531804 193898 532040 194134
rect 542410 194218 542646 194454
rect 542410 193898 542646 194134
rect 550252 194218 550488 194454
rect 550252 193898 550488 194134
rect 558094 194218 558330 194454
rect 558094 193898 558330 194134
rect 565936 194218 566172 194454
rect 565936 193898 566172 194134
rect 337189 187938 337425 188174
rect 337189 187618 337425 187854
rect 404786 187938 405022 188174
rect 404786 187618 405022 187854
rect 472383 187938 472619 188174
rect 472383 187618 472619 187854
rect 539980 187938 540216 188174
rect 539980 187618 540216 187854
rect 303391 184218 303627 184454
rect 303391 183898 303627 184134
rect 370988 184218 371224 184454
rect 370988 183898 371224 184134
rect 438585 184218 438821 184454
rect 438585 183898 438821 184134
rect 506182 184218 506418 184454
rect 506182 183898 506418 184134
rect 307407 177643 307643 177879
rect 315249 177643 315485 177879
rect 323091 177643 323327 177879
rect 330933 177643 331169 177879
rect 303486 174218 303722 174454
rect 303486 173898 303722 174134
rect 311328 174218 311564 174454
rect 311328 173898 311564 174134
rect 319170 174218 319406 174454
rect 319170 173898 319406 174134
rect 327012 174218 327248 174454
rect 327012 173898 327248 174134
rect 307407 167938 307643 168174
rect 307407 167618 307643 167854
rect 315249 167938 315485 168174
rect 315249 167618 315485 167854
rect 323091 167938 323327 168174
rect 323091 167618 323327 167854
rect 330933 167938 331169 168174
rect 330933 167618 331169 167854
rect 303486 164218 303722 164454
rect 303486 163898 303722 164134
rect 311328 164218 311564 164454
rect 311328 163898 311564 164134
rect 319170 164218 319406 164454
rect 319170 163898 319406 164134
rect 327012 164218 327248 164454
rect 327012 163898 327248 164134
rect 293034 63935 293270 64171
rect 277674 57938 277910 58174
rect 277674 57618 277910 57854
rect 308394 57938 308630 58174
rect 308394 57618 308630 57854
rect 293034 54218 293270 54454
rect 293034 53898 293270 54134
rect 277674 47938 277910 48174
rect 277674 47618 277910 47854
rect 308394 47938 308630 48174
rect 308394 47618 308630 47854
rect 293034 44218 293270 44454
rect 293034 43898 293270 44134
rect 277674 37938 277910 38174
rect 277674 37618 277910 37854
rect 308394 37938 308630 38174
rect 308394 37618 308630 37854
rect 293034 34218 293270 34454
rect 293034 33898 293270 34134
rect 341539 177643 341775 177879
rect 349381 177643 349617 177879
rect 357223 177643 357459 177879
rect 365065 177643 365301 177879
rect 375671 177643 375907 177879
rect 383513 177643 383749 177879
rect 391355 177643 391591 177879
rect 399197 177643 399433 177879
rect 409803 177643 410039 177879
rect 417645 177643 417881 177879
rect 425487 177643 425723 177879
rect 433329 177643 433565 177879
rect 443935 177643 444171 177879
rect 451777 177643 452013 177879
rect 459619 177643 459855 177879
rect 467461 177643 467697 177879
rect 478067 177643 478303 177879
rect 485909 177643 486145 177879
rect 493751 177643 493987 177879
rect 501593 177643 501829 177879
rect 512199 177643 512435 177879
rect 520041 177643 520277 177879
rect 527883 177643 528119 177879
rect 535725 177643 535961 177879
rect 546331 177643 546567 177879
rect 554173 177643 554409 177879
rect 562015 177643 562251 177879
rect 569857 177643 570093 177879
rect 337618 174218 337854 174454
rect 337618 173898 337854 174134
rect 345460 174218 345696 174454
rect 345460 173898 345696 174134
rect 353302 174218 353538 174454
rect 353302 173898 353538 174134
rect 361144 174218 361380 174454
rect 361144 173898 361380 174134
rect 371750 174218 371986 174454
rect 371750 173898 371986 174134
rect 379592 174218 379828 174454
rect 379592 173898 379828 174134
rect 387434 174218 387670 174454
rect 387434 173898 387670 174134
rect 395276 174218 395512 174454
rect 395276 173898 395512 174134
rect 405882 174218 406118 174454
rect 405882 173898 406118 174134
rect 413724 174218 413960 174454
rect 413724 173898 413960 174134
rect 421566 174218 421802 174454
rect 421566 173898 421802 174134
rect 429408 174218 429644 174454
rect 429408 173898 429644 174134
rect 440014 174218 440250 174454
rect 440014 173898 440250 174134
rect 447856 174218 448092 174454
rect 447856 173898 448092 174134
rect 455698 174218 455934 174454
rect 455698 173898 455934 174134
rect 463540 174218 463776 174454
rect 463540 173898 463776 174134
rect 474146 174218 474382 174454
rect 474146 173898 474382 174134
rect 481988 174218 482224 174454
rect 481988 173898 482224 174134
rect 489830 174218 490066 174454
rect 489830 173898 490066 174134
rect 497672 174218 497908 174454
rect 497672 173898 497908 174134
rect 508278 174218 508514 174454
rect 508278 173898 508514 174134
rect 516120 174218 516356 174454
rect 516120 173898 516356 174134
rect 523962 174218 524198 174454
rect 523962 173898 524198 174134
rect 531804 174218 532040 174454
rect 531804 173898 532040 174134
rect 542410 174218 542646 174454
rect 542410 173898 542646 174134
rect 550252 174218 550488 174454
rect 550252 173898 550488 174134
rect 558094 174218 558330 174454
rect 558094 173898 558330 174134
rect 565936 174218 566172 174454
rect 565936 173898 566172 174134
rect 341539 167938 341775 168174
rect 341539 167618 341775 167854
rect 349381 167938 349617 168174
rect 349381 167618 349617 167854
rect 357223 167938 357459 168174
rect 357223 167618 357459 167854
rect 365065 167938 365301 168174
rect 365065 167618 365301 167854
rect 375671 167938 375907 168174
rect 375671 167618 375907 167854
rect 383513 167938 383749 168174
rect 383513 167618 383749 167854
rect 391355 167938 391591 168174
rect 391355 167618 391591 167854
rect 399197 167938 399433 168174
rect 399197 167618 399433 167854
rect 409803 167938 410039 168174
rect 409803 167618 410039 167854
rect 417645 167938 417881 168174
rect 417645 167618 417881 167854
rect 425487 167938 425723 168174
rect 425487 167618 425723 167854
rect 433329 167938 433565 168174
rect 433329 167618 433565 167854
rect 443935 167938 444171 168174
rect 443935 167618 444171 167854
rect 451777 167938 452013 168174
rect 451777 167618 452013 167854
rect 459619 167938 459855 168174
rect 459619 167618 459855 167854
rect 467461 167938 467697 168174
rect 467461 167618 467697 167854
rect 478067 167938 478303 168174
rect 478067 167618 478303 167854
rect 485909 167938 486145 168174
rect 485909 167618 486145 167854
rect 493751 167938 493987 168174
rect 493751 167618 493987 167854
rect 501593 167938 501829 168174
rect 501593 167618 501829 167854
rect 512199 167938 512435 168174
rect 512199 167618 512435 167854
rect 520041 167938 520277 168174
rect 520041 167618 520277 167854
rect 527883 167938 528119 168174
rect 527883 167618 528119 167854
rect 535725 167938 535961 168174
rect 535725 167618 535961 167854
rect 546331 167938 546567 168174
rect 546331 167618 546567 167854
rect 554173 167938 554409 168174
rect 554173 167618 554409 167854
rect 562015 167938 562251 168174
rect 562015 167618 562251 167854
rect 569857 167938 570093 168174
rect 569857 167618 570093 167854
rect 337618 164218 337854 164454
rect 337618 163898 337854 164134
rect 345460 164218 345696 164454
rect 345460 163898 345696 164134
rect 353302 164218 353538 164454
rect 353302 163898 353538 164134
rect 361144 164218 361380 164454
rect 361144 163898 361380 164134
rect 371750 164218 371986 164454
rect 371750 163898 371986 164134
rect 379592 164218 379828 164454
rect 379592 163898 379828 164134
rect 387434 164218 387670 164454
rect 387434 163898 387670 164134
rect 395276 164218 395512 164454
rect 395276 163898 395512 164134
rect 405882 164218 406118 164454
rect 405882 163898 406118 164134
rect 413724 164218 413960 164454
rect 413724 163898 413960 164134
rect 421566 164218 421802 164454
rect 421566 163898 421802 164134
rect 429408 164218 429644 164454
rect 429408 163898 429644 164134
rect 440014 164218 440250 164454
rect 440014 163898 440250 164134
rect 447856 164218 448092 164454
rect 447856 163898 448092 164134
rect 455698 164218 455934 164454
rect 455698 163898 455934 164134
rect 463540 164218 463776 164454
rect 463540 163898 463776 164134
rect 474146 164218 474382 164454
rect 474146 163898 474382 164134
rect 481988 164218 482224 164454
rect 481988 163898 482224 164134
rect 489830 164218 490066 164454
rect 489830 163898 490066 164134
rect 497672 164218 497908 164454
rect 497672 163898 497908 164134
rect 508278 164218 508514 164454
rect 508278 163898 508514 164134
rect 516120 164218 516356 164454
rect 516120 163898 516356 164134
rect 523962 164218 524198 164454
rect 523962 163898 524198 164134
rect 531804 164218 532040 164454
rect 531804 163898 532040 164134
rect 542410 164218 542646 164454
rect 542410 163898 542646 164134
rect 550252 164218 550488 164454
rect 550252 163898 550488 164134
rect 558094 164218 558330 164454
rect 558094 163898 558330 164134
rect 565936 164218 566172 164454
rect 565936 163898 566172 164134
rect 585342 667938 585578 668174
rect 585662 667938 585898 668174
rect 585342 667618 585578 667854
rect 585662 667618 585898 667854
rect 585342 657938 585578 658174
rect 585662 657938 585898 658174
rect 585342 657618 585578 657854
rect 585662 657618 585898 657854
rect 585342 647938 585578 648174
rect 585662 647938 585898 648174
rect 585342 647618 585578 647854
rect 585662 647618 585898 647854
rect 585342 637938 585578 638174
rect 585662 637938 585898 638174
rect 585342 637618 585578 637854
rect 585662 637618 585898 637854
rect 585342 627938 585578 628174
rect 585662 627938 585898 628174
rect 585342 627618 585578 627854
rect 585662 627618 585898 627854
rect 585342 617938 585578 618174
rect 585662 617938 585898 618174
rect 585342 617618 585578 617854
rect 585662 617618 585898 617854
rect 585342 607938 585578 608174
rect 585662 607938 585898 608174
rect 585342 607618 585578 607854
rect 585662 607618 585898 607854
rect 585342 597938 585578 598174
rect 585662 597938 585898 598174
rect 585342 597618 585578 597854
rect 585662 597618 585898 597854
rect 585342 587938 585578 588174
rect 585662 587938 585898 588174
rect 585342 587618 585578 587854
rect 585662 587618 585898 587854
rect 585342 577938 585578 578174
rect 585662 577938 585898 578174
rect 585342 577618 585578 577854
rect 585662 577618 585898 577854
rect 585342 567938 585578 568174
rect 585662 567938 585898 568174
rect 585342 567618 585578 567854
rect 585662 567618 585898 567854
rect 585342 557938 585578 558174
rect 585662 557938 585898 558174
rect 585342 557618 585578 557854
rect 585662 557618 585898 557854
rect 585342 547938 585578 548174
rect 585662 547938 585898 548174
rect 585342 547618 585578 547854
rect 585662 547618 585898 547854
rect 585342 537938 585578 538174
rect 585662 537938 585898 538174
rect 585342 537618 585578 537854
rect 585662 537618 585898 537854
rect 585342 527938 585578 528174
rect 585662 527938 585898 528174
rect 585342 527618 585578 527854
rect 585662 527618 585898 527854
rect 585342 517938 585578 518174
rect 585662 517938 585898 518174
rect 585342 517618 585578 517854
rect 585662 517618 585898 517854
rect 585342 507938 585578 508174
rect 585662 507938 585898 508174
rect 585342 507618 585578 507854
rect 585662 507618 585898 507854
rect 585342 497938 585578 498174
rect 585662 497938 585898 498174
rect 585342 497618 585578 497854
rect 585662 497618 585898 497854
rect 585342 487938 585578 488174
rect 585662 487938 585898 488174
rect 585342 487618 585578 487854
rect 585662 487618 585898 487854
rect 585342 477938 585578 478174
rect 585662 477938 585898 478174
rect 585342 477618 585578 477854
rect 585662 477618 585898 477854
rect 585342 467938 585578 468174
rect 585662 467938 585898 468174
rect 585342 467618 585578 467854
rect 585662 467618 585898 467854
rect 585342 457938 585578 458174
rect 585662 457938 585898 458174
rect 585342 457618 585578 457854
rect 585662 457618 585898 457854
rect 585342 447938 585578 448174
rect 585662 447938 585898 448174
rect 585342 447618 585578 447854
rect 585662 447618 585898 447854
rect 585342 437938 585578 438174
rect 585662 437938 585898 438174
rect 585342 437618 585578 437854
rect 585662 437618 585898 437854
rect 585342 427938 585578 428174
rect 585662 427938 585898 428174
rect 585342 427618 585578 427854
rect 585662 427618 585898 427854
rect 585342 417938 585578 418174
rect 585662 417938 585898 418174
rect 585342 417618 585578 417854
rect 585662 417618 585898 417854
rect 585342 407938 585578 408174
rect 585662 407938 585898 408174
rect 585342 407618 585578 407854
rect 585662 407618 585898 407854
rect 585342 397938 585578 398174
rect 585662 397938 585898 398174
rect 585342 397618 585578 397854
rect 585662 397618 585898 397854
rect 585342 387938 585578 388174
rect 585662 387938 585898 388174
rect 585342 387618 585578 387854
rect 585662 387618 585898 387854
rect 585342 377938 585578 378174
rect 585662 377938 585898 378174
rect 585342 377618 585578 377854
rect 585662 377618 585898 377854
rect 585342 367938 585578 368174
rect 585662 367938 585898 368174
rect 585342 367618 585578 367854
rect 585662 367618 585898 367854
rect 585342 357938 585578 358174
rect 585662 357938 585898 358174
rect 585342 357618 585578 357854
rect 585662 357618 585898 357854
rect 585342 347938 585578 348174
rect 585662 347938 585898 348174
rect 585342 347618 585578 347854
rect 585662 347618 585898 347854
rect 585342 337938 585578 338174
rect 585662 337938 585898 338174
rect 585342 337618 585578 337854
rect 585662 337618 585898 337854
rect 585342 327938 585578 328174
rect 585662 327938 585898 328174
rect 585342 327618 585578 327854
rect 585662 327618 585898 327854
rect 585342 317938 585578 318174
rect 585662 317938 585898 318174
rect 585342 317618 585578 317854
rect 585662 317618 585898 317854
rect 585342 307938 585578 308174
rect 585662 307938 585898 308174
rect 585342 307618 585578 307854
rect 585662 307618 585898 307854
rect 585342 297938 585578 298174
rect 585662 297938 585898 298174
rect 585342 297618 585578 297854
rect 585662 297618 585898 297854
rect 585342 287938 585578 288174
rect 585662 287938 585898 288174
rect 585342 287618 585578 287854
rect 585662 287618 585898 287854
rect 585342 277938 585578 278174
rect 585662 277938 585898 278174
rect 585342 277618 585578 277854
rect 585662 277618 585898 277854
rect 585342 267938 585578 268174
rect 585662 267938 585898 268174
rect 585342 267618 585578 267854
rect 585662 267618 585898 267854
rect 585342 257938 585578 258174
rect 585662 257938 585898 258174
rect 585342 257618 585578 257854
rect 585662 257618 585898 257854
rect 585342 247938 585578 248174
rect 585662 247938 585898 248174
rect 585342 247618 585578 247854
rect 585662 247618 585898 247854
rect 585342 237938 585578 238174
rect 585662 237938 585898 238174
rect 585342 237618 585578 237854
rect 585662 237618 585898 237854
rect 585342 227938 585578 228174
rect 585662 227938 585898 228174
rect 585342 227618 585578 227854
rect 585662 227618 585898 227854
rect 585342 217938 585578 218174
rect 585662 217938 585898 218174
rect 585342 217618 585578 217854
rect 585662 217618 585898 217854
rect 585342 207938 585578 208174
rect 585662 207938 585898 208174
rect 585342 207618 585578 207854
rect 585662 207618 585898 207854
rect 585342 197938 585578 198174
rect 585662 197938 585898 198174
rect 585342 197618 585578 197854
rect 585662 197618 585898 197854
rect 585342 187938 585578 188174
rect 585662 187938 585898 188174
rect 585342 187618 585578 187854
rect 585662 187618 585898 187854
rect 585342 177938 585578 178174
rect 585662 177938 585898 178174
rect 585342 177618 585578 177854
rect 585662 177618 585898 177854
rect 585342 167938 585578 168174
rect 585662 167938 585898 168174
rect 585342 167618 585578 167854
rect 585662 167618 585898 167854
rect 585342 157938 585578 158174
rect 585662 157938 585898 158174
rect 585342 157618 585578 157854
rect 585662 157618 585898 157854
rect 585342 147938 585578 148174
rect 585662 147938 585898 148174
rect 585342 147618 585578 147854
rect 585662 147618 585898 147854
rect 585342 137938 585578 138174
rect 585662 137938 585898 138174
rect 585342 137618 585578 137854
rect 585662 137618 585898 137854
rect 585342 127938 585578 128174
rect 585662 127938 585898 128174
rect 585342 127618 585578 127854
rect 585662 127618 585898 127854
rect 585342 117938 585578 118174
rect 585662 117938 585898 118174
rect 585342 117618 585578 117854
rect 585662 117618 585898 117854
rect 585342 107938 585578 108174
rect 585662 107938 585898 108174
rect 585342 107618 585578 107854
rect 585662 107618 585898 107854
rect 585342 97938 585578 98174
rect 585662 97938 585898 98174
rect 585342 97618 585578 97854
rect 585662 97618 585898 97854
rect 585342 87938 585578 88174
rect 585662 87938 585898 88174
rect 585342 87618 585578 87854
rect 585662 87618 585898 87854
rect 585342 77938 585578 78174
rect 585662 77938 585898 78174
rect 585342 77618 585578 77854
rect 585662 77618 585898 77854
rect 585342 67938 585578 68174
rect 585662 67938 585898 68174
rect 585342 67618 585578 67854
rect 585662 67618 585898 67854
rect 585342 57938 585578 58174
rect 585662 57938 585898 58174
rect 585342 57618 585578 57854
rect 585662 57618 585898 57854
rect 585342 47938 585578 48174
rect 585662 47938 585898 48174
rect 585342 47618 585578 47854
rect 585662 47618 585898 47854
rect 585342 37938 585578 38174
rect 585662 37938 585898 38174
rect 585342 37618 585578 37854
rect 585662 37618 585898 37854
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 694218 586538 694454
rect 586622 694218 586858 694454
rect 586302 693898 586538 694134
rect 586622 693898 586858 694134
rect 586302 684218 586538 684454
rect 586622 684218 586858 684454
rect 586302 683898 586538 684134
rect 586622 683898 586858 684134
rect 586302 674218 586538 674454
rect 586622 674218 586858 674454
rect 586302 673898 586538 674134
rect 586622 673898 586858 674134
rect 586302 664218 586538 664454
rect 586622 664218 586858 664454
rect 586302 663898 586538 664134
rect 586622 663898 586858 664134
rect 586302 654218 586538 654454
rect 586622 654218 586858 654454
rect 586302 653898 586538 654134
rect 586622 653898 586858 654134
rect 586302 644218 586538 644454
rect 586622 644218 586858 644454
rect 586302 643898 586538 644134
rect 586622 643898 586858 644134
rect 586302 634218 586538 634454
rect 586622 634218 586858 634454
rect 586302 633898 586538 634134
rect 586622 633898 586858 634134
rect 586302 624218 586538 624454
rect 586622 624218 586858 624454
rect 586302 623898 586538 624134
rect 586622 623898 586858 624134
rect 586302 614218 586538 614454
rect 586622 614218 586858 614454
rect 586302 613898 586538 614134
rect 586622 613898 586858 614134
rect 586302 604218 586538 604454
rect 586622 604218 586858 604454
rect 586302 603898 586538 604134
rect 586622 603898 586858 604134
rect 586302 594218 586538 594454
rect 586622 594218 586858 594454
rect 586302 593898 586538 594134
rect 586622 593898 586858 594134
rect 586302 584218 586538 584454
rect 586622 584218 586858 584454
rect 586302 583898 586538 584134
rect 586622 583898 586858 584134
rect 586302 574218 586538 574454
rect 586622 574218 586858 574454
rect 586302 573898 586538 574134
rect 586622 573898 586858 574134
rect 586302 564218 586538 564454
rect 586622 564218 586858 564454
rect 586302 563898 586538 564134
rect 586622 563898 586858 564134
rect 586302 554218 586538 554454
rect 586622 554218 586858 554454
rect 586302 553898 586538 554134
rect 586622 553898 586858 554134
rect 586302 544218 586538 544454
rect 586622 544218 586858 544454
rect 586302 543898 586538 544134
rect 586622 543898 586858 544134
rect 586302 534218 586538 534454
rect 586622 534218 586858 534454
rect 586302 533898 586538 534134
rect 586622 533898 586858 534134
rect 586302 524218 586538 524454
rect 586622 524218 586858 524454
rect 586302 523898 586538 524134
rect 586622 523898 586858 524134
rect 586302 514218 586538 514454
rect 586622 514218 586858 514454
rect 586302 513898 586538 514134
rect 586622 513898 586858 514134
rect 586302 504218 586538 504454
rect 586622 504218 586858 504454
rect 586302 503898 586538 504134
rect 586622 503898 586858 504134
rect 586302 494218 586538 494454
rect 586622 494218 586858 494454
rect 586302 493898 586538 494134
rect 586622 493898 586858 494134
rect 586302 484218 586538 484454
rect 586622 484218 586858 484454
rect 586302 483898 586538 484134
rect 586622 483898 586858 484134
rect 586302 474218 586538 474454
rect 586622 474218 586858 474454
rect 586302 473898 586538 474134
rect 586622 473898 586858 474134
rect 586302 464218 586538 464454
rect 586622 464218 586858 464454
rect 586302 463898 586538 464134
rect 586622 463898 586858 464134
rect 586302 454218 586538 454454
rect 586622 454218 586858 454454
rect 586302 453898 586538 454134
rect 586622 453898 586858 454134
rect 586302 444218 586538 444454
rect 586622 444218 586858 444454
rect 586302 443898 586538 444134
rect 586622 443898 586858 444134
rect 586302 434218 586538 434454
rect 586622 434218 586858 434454
rect 586302 433898 586538 434134
rect 586622 433898 586858 434134
rect 586302 424218 586538 424454
rect 586622 424218 586858 424454
rect 586302 423898 586538 424134
rect 586622 423898 586858 424134
rect 586302 414218 586538 414454
rect 586622 414218 586858 414454
rect 586302 413898 586538 414134
rect 586622 413898 586858 414134
rect 586302 404218 586538 404454
rect 586622 404218 586858 404454
rect 586302 403898 586538 404134
rect 586622 403898 586858 404134
rect 586302 394218 586538 394454
rect 586622 394218 586858 394454
rect 586302 393898 586538 394134
rect 586622 393898 586858 394134
rect 586302 384218 586538 384454
rect 586622 384218 586858 384454
rect 586302 383898 586538 384134
rect 586622 383898 586858 384134
rect 586302 374218 586538 374454
rect 586622 374218 586858 374454
rect 586302 373898 586538 374134
rect 586622 373898 586858 374134
rect 586302 364218 586538 364454
rect 586622 364218 586858 364454
rect 586302 363898 586538 364134
rect 586622 363898 586858 364134
rect 586302 354218 586538 354454
rect 586622 354218 586858 354454
rect 586302 353898 586538 354134
rect 586622 353898 586858 354134
rect 586302 344218 586538 344454
rect 586622 344218 586858 344454
rect 586302 343898 586538 344134
rect 586622 343898 586858 344134
rect 586302 334218 586538 334454
rect 586622 334218 586858 334454
rect 586302 333898 586538 334134
rect 586622 333898 586858 334134
rect 586302 324218 586538 324454
rect 586622 324218 586858 324454
rect 586302 323898 586538 324134
rect 586622 323898 586858 324134
rect 586302 314218 586538 314454
rect 586622 314218 586858 314454
rect 586302 313898 586538 314134
rect 586622 313898 586858 314134
rect 586302 304218 586538 304454
rect 586622 304218 586858 304454
rect 586302 303898 586538 304134
rect 586622 303898 586858 304134
rect 586302 294218 586538 294454
rect 586622 294218 586858 294454
rect 586302 293898 586538 294134
rect 586622 293898 586858 294134
rect 586302 284218 586538 284454
rect 586622 284218 586858 284454
rect 586302 283898 586538 284134
rect 586622 283898 586858 284134
rect 586302 274218 586538 274454
rect 586622 274218 586858 274454
rect 586302 273898 586538 274134
rect 586622 273898 586858 274134
rect 586302 264218 586538 264454
rect 586622 264218 586858 264454
rect 586302 263898 586538 264134
rect 586622 263898 586858 264134
rect 586302 254218 586538 254454
rect 586622 254218 586858 254454
rect 586302 253898 586538 254134
rect 586622 253898 586858 254134
rect 586302 244218 586538 244454
rect 586622 244218 586858 244454
rect 586302 243898 586538 244134
rect 586622 243898 586858 244134
rect 586302 234218 586538 234454
rect 586622 234218 586858 234454
rect 586302 233898 586538 234134
rect 586622 233898 586858 234134
rect 586302 224218 586538 224454
rect 586622 224218 586858 224454
rect 586302 223898 586538 224134
rect 586622 223898 586858 224134
rect 586302 214218 586538 214454
rect 586622 214218 586858 214454
rect 586302 213898 586538 214134
rect 586622 213898 586858 214134
rect 586302 204218 586538 204454
rect 586622 204218 586858 204454
rect 586302 203898 586538 204134
rect 586622 203898 586858 204134
rect 586302 194218 586538 194454
rect 586622 194218 586858 194454
rect 586302 193898 586538 194134
rect 586622 193898 586858 194134
rect 586302 184218 586538 184454
rect 586622 184218 586858 184454
rect 586302 183898 586538 184134
rect 586622 183898 586858 184134
rect 586302 174218 586538 174454
rect 586622 174218 586858 174454
rect 586302 173898 586538 174134
rect 586622 173898 586858 174134
rect 586302 164218 586538 164454
rect 586622 164218 586858 164454
rect 586302 163898 586538 164134
rect 586622 163898 586858 164134
rect 586302 154218 586538 154454
rect 586622 154218 586858 154454
rect 586302 153898 586538 154134
rect 586622 153898 586858 154134
rect 586302 144218 586538 144454
rect 586622 144218 586858 144454
rect 586302 143898 586538 144134
rect 586622 143898 586858 144134
rect 586302 134218 586538 134454
rect 586622 134218 586858 134454
rect 586302 133898 586538 134134
rect 586622 133898 586858 134134
rect 586302 124218 586538 124454
rect 586622 124218 586858 124454
rect 586302 123898 586538 124134
rect 586622 123898 586858 124134
rect 586302 114218 586538 114454
rect 586622 114218 586858 114454
rect 586302 113898 586538 114134
rect 586622 113898 586858 114134
rect 586302 104218 586538 104454
rect 586622 104218 586858 104454
rect 586302 103898 586538 104134
rect 586622 103898 586858 104134
rect 586302 94218 586538 94454
rect 586622 94218 586858 94454
rect 586302 93898 586538 94134
rect 586622 93898 586858 94134
rect 586302 84218 586538 84454
rect 586622 84218 586858 84454
rect 586302 83898 586538 84134
rect 586622 83898 586858 84134
rect 586302 74218 586538 74454
rect 586622 74218 586858 74454
rect 586302 73898 586538 74134
rect 586622 73898 586858 74134
rect 586302 64218 586538 64454
rect 586622 64218 586858 64454
rect 586302 63898 586538 64134
rect 586622 63898 586858 64134
rect 586302 54218 586538 54454
rect 586622 54218 586858 54454
rect 586302 53898 586538 54134
rect 586622 53898 586858 54134
rect 586302 44218 586538 44454
rect 586622 44218 586858 44454
rect 586302 43898 586538 44134
rect 586622 43898 586858 44134
rect 586302 34218 586538 34454
rect 586622 34218 586858 34454
rect 586302 33898 586538 34134
rect 586622 33898 586858 34134
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698174 592650 698206
rect -8726 697938 -1974 698174
rect -1738 697938 -1654 698174
rect -1418 697938 585342 698174
rect 585578 697938 585662 698174
rect 585898 697938 592650 698174
rect -8726 697854 592650 697938
rect -8726 697618 -1974 697854
rect -1738 697618 -1654 697854
rect -1418 697618 585342 697854
rect 585578 697618 585662 697854
rect 585898 697618 592650 697854
rect -8726 697586 592650 697618
rect -8726 694454 592650 694486
rect -8726 694218 -2934 694454
rect -2698 694218 -2614 694454
rect -2378 694218 586302 694454
rect 586538 694218 586622 694454
rect 586858 694218 592650 694454
rect -8726 694134 592650 694218
rect -8726 693898 -2934 694134
rect -2698 693898 -2614 694134
rect -2378 693898 586302 694134
rect 586538 693898 586622 694134
rect 586858 693898 592650 694134
rect -8726 693866 592650 693898
rect -8726 688174 592650 688206
rect -8726 687938 -1974 688174
rect -1738 687938 -1654 688174
rect -1418 687938 585342 688174
rect 585578 687938 585662 688174
rect 585898 687938 592650 688174
rect -8726 687854 592650 687938
rect -8726 687618 -1974 687854
rect -1738 687618 -1654 687854
rect -1418 687618 585342 687854
rect 585578 687618 585662 687854
rect 585898 687618 592650 687854
rect -8726 687586 592650 687618
rect -8726 684454 592650 684486
rect -8726 684218 -2934 684454
rect -2698 684218 -2614 684454
rect -2378 684218 586302 684454
rect 586538 684218 586622 684454
rect 586858 684218 592650 684454
rect -8726 684134 592650 684218
rect -8726 683898 -2934 684134
rect -2698 683898 -2614 684134
rect -2378 683898 586302 684134
rect 586538 683898 586622 684134
rect 586858 683898 592650 684134
rect -8726 683866 592650 683898
rect -8726 678174 592650 678206
rect -8726 677938 -1974 678174
rect -1738 677938 -1654 678174
rect -1418 677938 585342 678174
rect 585578 677938 585662 678174
rect 585898 677938 592650 678174
rect -8726 677854 592650 677938
rect -8726 677618 -1974 677854
rect -1738 677618 -1654 677854
rect -1418 677618 585342 677854
rect 585578 677618 585662 677854
rect 585898 677618 592650 677854
rect -8726 677586 592650 677618
rect -8726 674454 592650 674486
rect -8726 674218 -2934 674454
rect -2698 674218 -2614 674454
rect -2378 674218 586302 674454
rect 586538 674218 586622 674454
rect 586858 674218 592650 674454
rect -8726 674134 592650 674218
rect -8726 673898 -2934 674134
rect -2698 673898 -2614 674134
rect -2378 673898 586302 674134
rect 586538 673898 586622 674134
rect 586858 673898 592650 674134
rect -8726 673866 592650 673898
rect -8726 668174 592650 668206
rect -8726 667938 -1974 668174
rect -1738 667938 -1654 668174
rect -1418 667938 585342 668174
rect 585578 667938 585662 668174
rect 585898 667938 592650 668174
rect -8726 667854 592650 667938
rect -8726 667618 -1974 667854
rect -1738 667618 -1654 667854
rect -1418 667618 585342 667854
rect 585578 667618 585662 667854
rect 585898 667618 592650 667854
rect -8726 667586 592650 667618
rect -8726 664454 592650 664486
rect -8726 664218 -2934 664454
rect -2698 664218 -2614 664454
rect -2378 664218 586302 664454
rect 586538 664218 586622 664454
rect 586858 664218 592650 664454
rect -8726 664134 592650 664218
rect -8726 663898 -2934 664134
rect -2698 663898 -2614 664134
rect -2378 663898 586302 664134
rect 586538 663898 586622 664134
rect 586858 663898 592650 664134
rect -8726 663866 592650 663898
rect -8726 658174 592650 658206
rect -8726 657938 -1974 658174
rect -1738 657938 -1654 658174
rect -1418 657938 585342 658174
rect 585578 657938 585662 658174
rect 585898 657938 592650 658174
rect -8726 657854 592650 657938
rect -8726 657618 -1974 657854
rect -1738 657618 -1654 657854
rect -1418 657618 585342 657854
rect 585578 657618 585662 657854
rect 585898 657618 592650 657854
rect -8726 657586 592650 657618
rect -8726 654454 592650 654486
rect -8726 654218 -2934 654454
rect -2698 654218 -2614 654454
rect -2378 654218 586302 654454
rect 586538 654218 586622 654454
rect 586858 654218 592650 654454
rect -8726 654134 592650 654218
rect -8726 653898 -2934 654134
rect -2698 653898 -2614 654134
rect -2378 653898 586302 654134
rect 586538 653898 586622 654134
rect 586858 653898 592650 654134
rect -8726 653866 592650 653898
rect -8726 648174 592650 648206
rect -8726 647938 -1974 648174
rect -1738 647938 -1654 648174
rect -1418 647938 585342 648174
rect 585578 647938 585662 648174
rect 585898 647938 592650 648174
rect -8726 647854 592650 647938
rect -8726 647618 -1974 647854
rect -1738 647618 -1654 647854
rect -1418 647618 585342 647854
rect 585578 647618 585662 647854
rect 585898 647618 592650 647854
rect -8726 647586 592650 647618
rect -8726 644454 592650 644486
rect -8726 644218 -2934 644454
rect -2698 644218 -2614 644454
rect -2378 644218 586302 644454
rect 586538 644218 586622 644454
rect 586858 644218 592650 644454
rect -8726 644134 592650 644218
rect -8726 643898 -2934 644134
rect -2698 643898 -2614 644134
rect -2378 643898 586302 644134
rect 586538 643898 586622 644134
rect 586858 643898 592650 644134
rect -8726 643866 592650 643898
rect -8726 638174 592650 638206
rect -8726 637938 -1974 638174
rect -1738 637938 -1654 638174
rect -1418 637938 585342 638174
rect 585578 637938 585662 638174
rect 585898 637938 592650 638174
rect -8726 637854 592650 637938
rect -8726 637618 -1974 637854
rect -1738 637618 -1654 637854
rect -1418 637618 585342 637854
rect 585578 637618 585662 637854
rect 585898 637618 592650 637854
rect -8726 637586 592650 637618
rect -8726 634454 592650 634486
rect -8726 634218 -2934 634454
rect -2698 634218 -2614 634454
rect -2378 634218 586302 634454
rect 586538 634218 586622 634454
rect 586858 634218 592650 634454
rect -8726 634134 592650 634218
rect -8726 633898 -2934 634134
rect -2698 633898 -2614 634134
rect -2378 633898 586302 634134
rect 586538 633898 586622 634134
rect 586858 633898 592650 634134
rect -8726 633866 592650 633898
rect -8726 628174 592650 628206
rect -8726 627938 -1974 628174
rect -1738 627938 -1654 628174
rect -1418 627938 585342 628174
rect 585578 627938 585662 628174
rect 585898 627938 592650 628174
rect -8726 627854 592650 627938
rect -8726 627618 -1974 627854
rect -1738 627618 -1654 627854
rect -1418 627618 585342 627854
rect 585578 627618 585662 627854
rect 585898 627618 592650 627854
rect -8726 627586 592650 627618
rect -8726 624454 592650 624486
rect -8726 624218 -2934 624454
rect -2698 624218 -2614 624454
rect -2378 624218 586302 624454
rect 586538 624218 586622 624454
rect 586858 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -2934 624134
rect -2698 623898 -2614 624134
rect -2378 623898 586302 624134
rect 586538 623898 586622 624134
rect 586858 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 618174 592650 618206
rect -8726 617938 -1974 618174
rect -1738 617938 -1654 618174
rect -1418 617938 585342 618174
rect 585578 617938 585662 618174
rect 585898 617938 592650 618174
rect -8726 617854 592650 617938
rect -8726 617618 -1974 617854
rect -1738 617618 -1654 617854
rect -1418 617618 585342 617854
rect 585578 617618 585662 617854
rect 585898 617618 592650 617854
rect -8726 617586 592650 617618
rect -8726 614454 592650 614486
rect -8726 614218 -2934 614454
rect -2698 614218 -2614 614454
rect -2378 614218 586302 614454
rect 586538 614218 586622 614454
rect 586858 614218 592650 614454
rect -8726 614134 592650 614218
rect -8726 613898 -2934 614134
rect -2698 613898 -2614 614134
rect -2378 613898 586302 614134
rect 586538 613898 586622 614134
rect 586858 613898 592650 614134
rect -8726 613866 592650 613898
rect -8726 608174 592650 608206
rect -8726 607938 -1974 608174
rect -1738 607938 -1654 608174
rect -1418 607938 585342 608174
rect 585578 607938 585662 608174
rect 585898 607938 592650 608174
rect -8726 607854 592650 607938
rect -8726 607618 -1974 607854
rect -1738 607618 -1654 607854
rect -1418 607618 585342 607854
rect 585578 607618 585662 607854
rect 585898 607618 592650 607854
rect -8726 607586 592650 607618
rect -8726 604454 592650 604486
rect -8726 604218 -2934 604454
rect -2698 604218 -2614 604454
rect -2378 604218 586302 604454
rect 586538 604218 586622 604454
rect 586858 604218 592650 604454
rect -8726 604134 592650 604218
rect -8726 603898 -2934 604134
rect -2698 603898 -2614 604134
rect -2378 603898 586302 604134
rect 586538 603898 586622 604134
rect 586858 603898 592650 604134
rect -8726 603866 592650 603898
rect -8726 598174 592650 598206
rect -8726 597938 -1974 598174
rect -1738 597938 -1654 598174
rect -1418 597938 585342 598174
rect 585578 597938 585662 598174
rect 585898 597938 592650 598174
rect -8726 597854 592650 597938
rect -8726 597618 -1974 597854
rect -1738 597618 -1654 597854
rect -1418 597618 585342 597854
rect 585578 597618 585662 597854
rect 585898 597618 592650 597854
rect -8726 597586 592650 597618
rect -8726 594454 592650 594486
rect -8726 594218 -2934 594454
rect -2698 594218 -2614 594454
rect -2378 594218 586302 594454
rect 586538 594218 586622 594454
rect 586858 594218 592650 594454
rect -8726 594134 592650 594218
rect -8726 593898 -2934 594134
rect -2698 593898 -2614 594134
rect -2378 593898 586302 594134
rect 586538 593898 586622 594134
rect 586858 593898 592650 594134
rect -8726 593866 592650 593898
rect -8726 588174 592650 588206
rect -8726 587938 -1974 588174
rect -1738 587938 -1654 588174
rect -1418 587938 585342 588174
rect 585578 587938 585662 588174
rect 585898 587938 592650 588174
rect -8726 587854 592650 587938
rect -8726 587618 -1974 587854
rect -1738 587618 -1654 587854
rect -1418 587618 585342 587854
rect 585578 587618 585662 587854
rect 585898 587618 592650 587854
rect -8726 587586 592650 587618
rect -8726 584454 592650 584486
rect -8726 584218 -2934 584454
rect -2698 584218 -2614 584454
rect -2378 584218 586302 584454
rect 586538 584218 586622 584454
rect 586858 584218 592650 584454
rect -8726 584134 592650 584218
rect -8726 583898 -2934 584134
rect -2698 583898 -2614 584134
rect -2378 583898 586302 584134
rect 586538 583898 586622 584134
rect 586858 583898 592650 584134
rect -8726 583866 592650 583898
rect -8726 578174 592650 578206
rect -8726 577938 -1974 578174
rect -1738 577938 -1654 578174
rect -1418 577938 585342 578174
rect 585578 577938 585662 578174
rect 585898 577938 592650 578174
rect -8726 577854 592650 577938
rect -8726 577618 -1974 577854
rect -1738 577618 -1654 577854
rect -1418 577618 585342 577854
rect 585578 577618 585662 577854
rect 585898 577618 592650 577854
rect -8726 577586 592650 577618
rect -8726 574454 592650 574486
rect -8726 574218 -2934 574454
rect -2698 574218 -2614 574454
rect -2378 574218 586302 574454
rect 586538 574218 586622 574454
rect 586858 574218 592650 574454
rect -8726 574134 592650 574218
rect -8726 573898 -2934 574134
rect -2698 573898 -2614 574134
rect -2378 573898 586302 574134
rect 586538 573898 586622 574134
rect 586858 573898 592650 574134
rect -8726 573866 592650 573898
rect -8726 568174 592650 568206
rect -8726 567938 -1974 568174
rect -1738 567938 -1654 568174
rect -1418 567938 585342 568174
rect 585578 567938 585662 568174
rect 585898 567938 592650 568174
rect -8726 567854 592650 567938
rect -8726 567618 -1974 567854
rect -1738 567618 -1654 567854
rect -1418 567618 585342 567854
rect 585578 567618 585662 567854
rect 585898 567618 592650 567854
rect -8726 567586 592650 567618
rect -8726 564454 592650 564486
rect -8726 564218 -2934 564454
rect -2698 564218 -2614 564454
rect -2378 564218 586302 564454
rect 586538 564218 586622 564454
rect 586858 564218 592650 564454
rect -8726 564134 592650 564218
rect -8726 563898 -2934 564134
rect -2698 563898 -2614 564134
rect -2378 563898 586302 564134
rect 586538 563898 586622 564134
rect 586858 563898 592650 564134
rect -8726 563866 592650 563898
rect -8726 558174 592650 558206
rect -8726 557938 -1974 558174
rect -1738 557938 -1654 558174
rect -1418 557938 585342 558174
rect 585578 557938 585662 558174
rect 585898 557938 592650 558174
rect -8726 557854 592650 557938
rect -8726 557618 -1974 557854
rect -1738 557618 -1654 557854
rect -1418 557618 585342 557854
rect 585578 557618 585662 557854
rect 585898 557618 592650 557854
rect -8726 557586 592650 557618
rect -8726 554454 592650 554486
rect -8726 554218 -2934 554454
rect -2698 554218 -2614 554454
rect -2378 554218 586302 554454
rect 586538 554218 586622 554454
rect 586858 554218 592650 554454
rect -8726 554134 592650 554218
rect -8726 553898 -2934 554134
rect -2698 553898 -2614 554134
rect -2378 553898 586302 554134
rect 586538 553898 586622 554134
rect 586858 553898 592650 554134
rect -8726 553866 592650 553898
rect -8726 548174 592650 548206
rect -8726 547938 -1974 548174
rect -1738 547938 -1654 548174
rect -1418 547938 585342 548174
rect 585578 547938 585662 548174
rect 585898 547938 592650 548174
rect -8726 547854 592650 547938
rect -8726 547618 -1974 547854
rect -1738 547618 -1654 547854
rect -1418 547618 585342 547854
rect 585578 547618 585662 547854
rect 585898 547618 592650 547854
rect -8726 547586 592650 547618
rect -8726 544454 592650 544486
rect -8726 544218 -2934 544454
rect -2698 544218 -2614 544454
rect -2378 544218 586302 544454
rect 586538 544218 586622 544454
rect 586858 544218 592650 544454
rect -8726 544134 592650 544218
rect -8726 543898 -2934 544134
rect -2698 543898 -2614 544134
rect -2378 543898 586302 544134
rect 586538 543898 586622 544134
rect 586858 543898 592650 544134
rect -8726 543866 592650 543898
rect -8726 538174 592650 538206
rect -8726 537938 -1974 538174
rect -1738 537938 -1654 538174
rect -1418 537938 585342 538174
rect 585578 537938 585662 538174
rect 585898 537938 592650 538174
rect -8726 537854 592650 537938
rect -8726 537618 -1974 537854
rect -1738 537618 -1654 537854
rect -1418 537618 585342 537854
rect 585578 537618 585662 537854
rect 585898 537618 592650 537854
rect -8726 537586 592650 537618
rect -8726 534454 592650 534486
rect -8726 534218 -2934 534454
rect -2698 534218 -2614 534454
rect -2378 534218 586302 534454
rect 586538 534218 586622 534454
rect 586858 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -2934 534134
rect -2698 533898 -2614 534134
rect -2378 533898 586302 534134
rect 586538 533898 586622 534134
rect 586858 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 528174 592650 528206
rect -8726 527938 -1974 528174
rect -1738 527938 -1654 528174
rect -1418 527938 585342 528174
rect 585578 527938 585662 528174
rect 585898 527938 592650 528174
rect -8726 527854 592650 527938
rect -8726 527618 -1974 527854
rect -1738 527618 -1654 527854
rect -1418 527618 585342 527854
rect 585578 527618 585662 527854
rect 585898 527618 592650 527854
rect -8726 527586 592650 527618
rect -8726 524454 592650 524486
rect -8726 524218 -2934 524454
rect -2698 524218 -2614 524454
rect -2378 524218 586302 524454
rect 586538 524218 586622 524454
rect 586858 524218 592650 524454
rect -8726 524134 592650 524218
rect -8726 523898 -2934 524134
rect -2698 523898 -2614 524134
rect -2378 523898 586302 524134
rect 586538 523898 586622 524134
rect 586858 523898 592650 524134
rect -8726 523866 592650 523898
rect -8726 518174 592650 518206
rect -8726 517938 -1974 518174
rect -1738 517938 -1654 518174
rect -1418 517938 585342 518174
rect 585578 517938 585662 518174
rect 585898 517938 592650 518174
rect -8726 517854 592650 517938
rect -8726 517618 -1974 517854
rect -1738 517618 -1654 517854
rect -1418 517618 585342 517854
rect 585578 517618 585662 517854
rect 585898 517618 592650 517854
rect -8726 517586 592650 517618
rect -8726 514454 592650 514486
rect -8726 514218 -2934 514454
rect -2698 514218 -2614 514454
rect -2378 514218 586302 514454
rect 586538 514218 586622 514454
rect 586858 514218 592650 514454
rect -8726 514134 592650 514218
rect -8726 513898 -2934 514134
rect -2698 513898 -2614 514134
rect -2378 513898 586302 514134
rect 586538 513898 586622 514134
rect 586858 513898 592650 514134
rect -8726 513866 592650 513898
rect -8726 508174 592650 508206
rect -8726 507938 -1974 508174
rect -1738 507938 -1654 508174
rect -1418 507938 585342 508174
rect 585578 507938 585662 508174
rect 585898 507938 592650 508174
rect -8726 507854 592650 507938
rect -8726 507618 -1974 507854
rect -1738 507618 -1654 507854
rect -1418 507618 585342 507854
rect 585578 507618 585662 507854
rect 585898 507618 592650 507854
rect -8726 507586 592650 507618
rect -8726 504454 592650 504486
rect -8726 504218 -2934 504454
rect -2698 504218 -2614 504454
rect -2378 504218 586302 504454
rect 586538 504218 586622 504454
rect 586858 504218 592650 504454
rect -8726 504134 592650 504218
rect -8726 503898 -2934 504134
rect -2698 503898 -2614 504134
rect -2378 503898 586302 504134
rect 586538 503898 586622 504134
rect 586858 503898 592650 504134
rect -8726 503866 592650 503898
rect -8726 498174 592650 498206
rect -8726 497938 -1974 498174
rect -1738 497938 -1654 498174
rect -1418 497938 585342 498174
rect 585578 497938 585662 498174
rect 585898 497938 592650 498174
rect -8726 497854 592650 497938
rect -8726 497618 -1974 497854
rect -1738 497618 -1654 497854
rect -1418 497618 585342 497854
rect 585578 497618 585662 497854
rect 585898 497618 592650 497854
rect -8726 497586 592650 497618
rect -8726 494454 592650 494486
rect -8726 494218 -2934 494454
rect -2698 494218 -2614 494454
rect -2378 494218 586302 494454
rect 586538 494218 586622 494454
rect 586858 494218 592650 494454
rect -8726 494134 592650 494218
rect -8726 493898 -2934 494134
rect -2698 493898 -2614 494134
rect -2378 493898 586302 494134
rect 586538 493898 586622 494134
rect 586858 493898 592650 494134
rect -8726 493866 592650 493898
rect -8726 488174 592650 488206
rect -8726 487938 -1974 488174
rect -1738 487938 -1654 488174
rect -1418 487938 585342 488174
rect 585578 487938 585662 488174
rect 585898 487938 592650 488174
rect -8726 487854 592650 487938
rect -8726 487618 -1974 487854
rect -1738 487618 -1654 487854
rect -1418 487618 585342 487854
rect 585578 487618 585662 487854
rect 585898 487618 592650 487854
rect -8726 487586 592650 487618
rect -8726 484454 592650 484486
rect -8726 484218 -2934 484454
rect -2698 484218 -2614 484454
rect -2378 484218 586302 484454
rect 586538 484218 586622 484454
rect 586858 484218 592650 484454
rect -8726 484134 592650 484218
rect -8726 483898 -2934 484134
rect -2698 483898 -2614 484134
rect -2378 483898 586302 484134
rect 586538 483898 586622 484134
rect 586858 483898 592650 484134
rect -8726 483866 592650 483898
rect -8726 478174 592650 478206
rect -8726 477938 -1974 478174
rect -1738 477938 -1654 478174
rect -1418 477938 585342 478174
rect 585578 477938 585662 478174
rect 585898 477938 592650 478174
rect -8726 477854 592650 477938
rect -8726 477618 -1974 477854
rect -1738 477618 -1654 477854
rect -1418 477618 585342 477854
rect 585578 477618 585662 477854
rect 585898 477618 592650 477854
rect -8726 477586 592650 477618
rect -8726 474454 592650 474486
rect -8726 474218 -2934 474454
rect -2698 474218 -2614 474454
rect -2378 474218 586302 474454
rect 586538 474218 586622 474454
rect 586858 474218 592650 474454
rect -8726 474134 592650 474218
rect -8726 473898 -2934 474134
rect -2698 473898 -2614 474134
rect -2378 473898 586302 474134
rect 586538 473898 586622 474134
rect 586858 473898 592650 474134
rect -8726 473866 592650 473898
rect -8726 468174 592650 468206
rect -8726 467938 -1974 468174
rect -1738 467938 -1654 468174
rect -1418 467938 585342 468174
rect 585578 467938 585662 468174
rect 585898 467938 592650 468174
rect -8726 467854 592650 467938
rect -8726 467618 -1974 467854
rect -1738 467618 -1654 467854
rect -1418 467618 585342 467854
rect 585578 467618 585662 467854
rect 585898 467618 592650 467854
rect -8726 467586 592650 467618
rect -8726 464454 592650 464486
rect -8726 464218 -2934 464454
rect -2698 464218 -2614 464454
rect -2378 464218 586302 464454
rect 586538 464218 586622 464454
rect 586858 464218 592650 464454
rect -8726 464134 592650 464218
rect -8726 463898 -2934 464134
rect -2698 463898 -2614 464134
rect -2378 463898 586302 464134
rect 586538 463898 586622 464134
rect 586858 463898 592650 464134
rect -8726 463866 592650 463898
rect -8726 458174 592650 458206
rect -8726 457938 -1974 458174
rect -1738 457938 -1654 458174
rect -1418 457938 585342 458174
rect 585578 457938 585662 458174
rect 585898 457938 592650 458174
rect -8726 457854 592650 457938
rect -8726 457618 -1974 457854
rect -1738 457618 -1654 457854
rect -1418 457618 585342 457854
rect 585578 457618 585662 457854
rect 585898 457618 592650 457854
rect -8726 457586 592650 457618
rect -8726 454454 592650 454486
rect -8726 454218 -2934 454454
rect -2698 454218 -2614 454454
rect -2378 454218 586302 454454
rect 586538 454218 586622 454454
rect 586858 454218 592650 454454
rect -8726 454134 592650 454218
rect -8726 453898 -2934 454134
rect -2698 453898 -2614 454134
rect -2378 453898 586302 454134
rect 586538 453898 586622 454134
rect 586858 453898 592650 454134
rect -8726 453866 592650 453898
rect -8726 448174 592650 448206
rect -8726 447938 -1974 448174
rect -1738 447938 -1654 448174
rect -1418 447938 585342 448174
rect 585578 447938 585662 448174
rect 585898 447938 592650 448174
rect -8726 447854 592650 447938
rect -8726 447618 -1974 447854
rect -1738 447618 -1654 447854
rect -1418 447618 585342 447854
rect 585578 447618 585662 447854
rect 585898 447618 592650 447854
rect -8726 447586 592650 447618
rect -8726 444454 592650 444486
rect -8726 444218 -2934 444454
rect -2698 444218 -2614 444454
rect -2378 444218 586302 444454
rect 586538 444218 586622 444454
rect 586858 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -2934 444134
rect -2698 443898 -2614 444134
rect -2378 443898 586302 444134
rect 586538 443898 586622 444134
rect 586858 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 438174 592650 438206
rect -8726 437938 -1974 438174
rect -1738 437938 -1654 438174
rect -1418 437938 585342 438174
rect 585578 437938 585662 438174
rect 585898 437938 592650 438174
rect -8726 437854 592650 437938
rect -8726 437618 -1974 437854
rect -1738 437618 -1654 437854
rect -1418 437618 585342 437854
rect 585578 437618 585662 437854
rect 585898 437618 592650 437854
rect -8726 437586 592650 437618
rect -8726 434454 592650 434486
rect -8726 434218 -2934 434454
rect -2698 434218 -2614 434454
rect -2378 434218 586302 434454
rect 586538 434218 586622 434454
rect 586858 434218 592650 434454
rect -8726 434134 592650 434218
rect -8726 433898 -2934 434134
rect -2698 433898 -2614 434134
rect -2378 433898 586302 434134
rect 586538 433898 586622 434134
rect 586858 433898 592650 434134
rect -8726 433866 592650 433898
rect -8726 428174 592650 428206
rect -8726 427938 -1974 428174
rect -1738 427938 -1654 428174
rect -1418 427938 585342 428174
rect 585578 427938 585662 428174
rect 585898 427938 592650 428174
rect -8726 427854 592650 427938
rect -8726 427618 -1974 427854
rect -1738 427618 -1654 427854
rect -1418 427618 585342 427854
rect 585578 427618 585662 427854
rect 585898 427618 592650 427854
rect -8726 427586 592650 427618
rect -8726 424454 592650 424486
rect -8726 424218 -2934 424454
rect -2698 424218 -2614 424454
rect -2378 424218 586302 424454
rect 586538 424218 586622 424454
rect 586858 424218 592650 424454
rect -8726 424134 592650 424218
rect -8726 423898 -2934 424134
rect -2698 423898 -2614 424134
rect -2378 423898 586302 424134
rect 586538 423898 586622 424134
rect 586858 423898 592650 424134
rect -8726 423866 592650 423898
rect -8726 418174 592650 418206
rect -8726 417938 -1974 418174
rect -1738 417938 -1654 418174
rect -1418 417938 585342 418174
rect 585578 417938 585662 418174
rect 585898 417938 592650 418174
rect -8726 417854 592650 417938
rect -8726 417618 -1974 417854
rect -1738 417618 -1654 417854
rect -1418 417618 585342 417854
rect 585578 417618 585662 417854
rect 585898 417618 592650 417854
rect -8726 417586 592650 417618
rect -8726 414454 592650 414486
rect -8726 414218 -2934 414454
rect -2698 414218 -2614 414454
rect -2378 414218 586302 414454
rect 586538 414218 586622 414454
rect 586858 414218 592650 414454
rect -8726 414134 592650 414218
rect -8726 413898 -2934 414134
rect -2698 413898 -2614 414134
rect -2378 413898 586302 414134
rect 586538 413898 586622 414134
rect 586858 413898 592650 414134
rect -8726 413866 592650 413898
rect -8726 408174 592650 408206
rect -8726 407938 -1974 408174
rect -1738 407938 -1654 408174
rect -1418 407938 585342 408174
rect 585578 407938 585662 408174
rect 585898 407938 592650 408174
rect -8726 407854 592650 407938
rect -8726 407618 -1974 407854
rect -1738 407618 -1654 407854
rect -1418 407618 585342 407854
rect 585578 407618 585662 407854
rect 585898 407618 592650 407854
rect -8726 407586 592650 407618
rect -8726 404454 592650 404486
rect -8726 404218 -2934 404454
rect -2698 404218 -2614 404454
rect -2378 404218 586302 404454
rect 586538 404218 586622 404454
rect 586858 404218 592650 404454
rect -8726 404134 592650 404218
rect -8726 403898 -2934 404134
rect -2698 403898 -2614 404134
rect -2378 403898 586302 404134
rect 586538 403898 586622 404134
rect 586858 403898 592650 404134
rect -8726 403866 592650 403898
rect -8726 398174 592650 398206
rect -8726 397938 -1974 398174
rect -1738 397938 -1654 398174
rect -1418 397938 585342 398174
rect 585578 397938 585662 398174
rect 585898 397938 592650 398174
rect -8726 397854 592650 397938
rect -8726 397618 -1974 397854
rect -1738 397618 -1654 397854
rect -1418 397618 585342 397854
rect 585578 397618 585662 397854
rect 585898 397618 592650 397854
rect -8726 397586 592650 397618
rect -8726 394454 592650 394486
rect -8726 394218 -2934 394454
rect -2698 394218 -2614 394454
rect -2378 394218 586302 394454
rect 586538 394218 586622 394454
rect 586858 394218 592650 394454
rect -8726 394134 592650 394218
rect -8726 393898 -2934 394134
rect -2698 393898 -2614 394134
rect -2378 393898 586302 394134
rect 586538 393898 586622 394134
rect 586858 393898 592650 394134
rect -8726 393866 592650 393898
rect -8726 388174 592650 388206
rect -8726 387938 -1974 388174
rect -1738 387938 -1654 388174
rect -1418 387938 585342 388174
rect 585578 387938 585662 388174
rect 585898 387938 592650 388174
rect -8726 387854 592650 387938
rect -8726 387618 -1974 387854
rect -1738 387618 -1654 387854
rect -1418 387618 585342 387854
rect 585578 387618 585662 387854
rect 585898 387618 592650 387854
rect -8726 387586 592650 387618
rect -8726 384454 592650 384486
rect -8726 384218 -2934 384454
rect -2698 384218 -2614 384454
rect -2378 384218 586302 384454
rect 586538 384218 586622 384454
rect 586858 384218 592650 384454
rect -8726 384134 592650 384218
rect -8726 383898 -2934 384134
rect -2698 383898 -2614 384134
rect -2378 383898 586302 384134
rect 586538 383898 586622 384134
rect 586858 383898 592650 384134
rect -8726 383866 592650 383898
rect -8726 378174 592650 378206
rect -8726 377938 -1974 378174
rect -1738 377938 -1654 378174
rect -1418 377938 585342 378174
rect 585578 377938 585662 378174
rect 585898 377938 592650 378174
rect -8726 377854 592650 377938
rect -8726 377618 -1974 377854
rect -1738 377618 -1654 377854
rect -1418 377618 585342 377854
rect 585578 377618 585662 377854
rect 585898 377618 592650 377854
rect -8726 377586 592650 377618
rect -8726 374454 592650 374486
rect -8726 374218 -2934 374454
rect -2698 374218 -2614 374454
rect -2378 374218 586302 374454
rect 586538 374218 586622 374454
rect 586858 374218 592650 374454
rect -8726 374134 592650 374218
rect -8726 373898 -2934 374134
rect -2698 373898 -2614 374134
rect -2378 373898 586302 374134
rect 586538 373898 586622 374134
rect 586858 373898 592650 374134
rect -8726 373866 592650 373898
rect -8726 368174 592650 368206
rect -8726 367938 -1974 368174
rect -1738 367938 -1654 368174
rect -1418 367938 585342 368174
rect 585578 367938 585662 368174
rect 585898 367938 592650 368174
rect -8726 367854 592650 367938
rect -8726 367618 -1974 367854
rect -1738 367618 -1654 367854
rect -1418 367618 585342 367854
rect 585578 367618 585662 367854
rect 585898 367618 592650 367854
rect -8726 367586 592650 367618
rect -8726 364454 592650 364486
rect -8726 364218 -2934 364454
rect -2698 364218 -2614 364454
rect -2378 364218 586302 364454
rect 586538 364218 586622 364454
rect 586858 364218 592650 364454
rect -8726 364134 592650 364218
rect -8726 363898 -2934 364134
rect -2698 363898 -2614 364134
rect -2378 363898 586302 364134
rect 586538 363898 586622 364134
rect 586858 363898 592650 364134
rect -8726 363866 592650 363898
rect -8726 358174 592650 358206
rect -8726 357938 -1974 358174
rect -1738 357938 -1654 358174
rect -1418 357938 585342 358174
rect 585578 357938 585662 358174
rect 585898 357938 592650 358174
rect -8726 357854 592650 357938
rect -8726 357618 -1974 357854
rect -1738 357618 -1654 357854
rect -1418 357618 585342 357854
rect 585578 357618 585662 357854
rect 585898 357618 592650 357854
rect -8726 357586 592650 357618
rect -8726 354454 592650 354486
rect -8726 354218 -2934 354454
rect -2698 354218 -2614 354454
rect -2378 354218 586302 354454
rect 586538 354218 586622 354454
rect 586858 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -2934 354134
rect -2698 353898 -2614 354134
rect -2378 353898 586302 354134
rect 586538 353898 586622 354134
rect 586858 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 348174 592650 348206
rect -8726 347938 -1974 348174
rect -1738 347938 -1654 348174
rect -1418 347938 585342 348174
rect 585578 347938 585662 348174
rect 585898 347938 592650 348174
rect -8726 347854 592650 347938
rect -8726 347618 -1974 347854
rect -1738 347618 -1654 347854
rect -1418 347618 585342 347854
rect 585578 347618 585662 347854
rect 585898 347618 592650 347854
rect -8726 347586 592650 347618
rect -8726 344454 592650 344486
rect -8726 344218 -2934 344454
rect -2698 344218 -2614 344454
rect -2378 344218 586302 344454
rect 586538 344218 586622 344454
rect 586858 344218 592650 344454
rect -8726 344134 592650 344218
rect -8726 343898 -2934 344134
rect -2698 343898 -2614 344134
rect -2378 343898 586302 344134
rect 586538 343898 586622 344134
rect 586858 343898 592650 344134
rect -8726 343866 592650 343898
rect -8726 338174 592650 338206
rect -8726 337938 -1974 338174
rect -1738 337938 -1654 338174
rect -1418 337938 585342 338174
rect 585578 337938 585662 338174
rect 585898 337938 592650 338174
rect -8726 337854 592650 337938
rect -8726 337618 -1974 337854
rect -1738 337618 -1654 337854
rect -1418 337618 585342 337854
rect 585578 337618 585662 337854
rect 585898 337618 592650 337854
rect -8726 337586 592650 337618
rect -8726 334454 592650 334486
rect -8726 334218 -2934 334454
rect -2698 334218 -2614 334454
rect -2378 334218 586302 334454
rect 586538 334218 586622 334454
rect 586858 334218 592650 334454
rect -8726 334134 592650 334218
rect -8726 333898 -2934 334134
rect -2698 333898 -2614 334134
rect -2378 333898 586302 334134
rect 586538 333898 586622 334134
rect 586858 333898 592650 334134
rect -8726 333866 592650 333898
rect -8726 328174 592650 328206
rect -8726 327938 -1974 328174
rect -1738 327938 -1654 328174
rect -1418 327938 585342 328174
rect 585578 327938 585662 328174
rect 585898 327938 592650 328174
rect -8726 327854 592650 327938
rect -8726 327618 -1974 327854
rect -1738 327618 -1654 327854
rect -1418 327618 585342 327854
rect 585578 327618 585662 327854
rect 585898 327618 592650 327854
rect -8726 327586 592650 327618
rect -8726 324454 592650 324486
rect -8726 324218 -2934 324454
rect -2698 324218 -2614 324454
rect -2378 324218 586302 324454
rect 586538 324218 586622 324454
rect 586858 324218 592650 324454
rect -8726 324134 592650 324218
rect -8726 323898 -2934 324134
rect -2698 323898 -2614 324134
rect -2378 323898 586302 324134
rect 586538 323898 586622 324134
rect 586858 323898 592650 324134
rect -8726 323866 592650 323898
rect -8726 318174 592650 318206
rect -8726 317938 -1974 318174
rect -1738 317938 -1654 318174
rect -1418 317938 585342 318174
rect 585578 317938 585662 318174
rect 585898 317938 592650 318174
rect -8726 317854 592650 317938
rect -8726 317618 -1974 317854
rect -1738 317618 -1654 317854
rect -1418 317618 585342 317854
rect 585578 317618 585662 317854
rect 585898 317618 592650 317854
rect -8726 317586 592650 317618
rect -8726 314454 592650 314486
rect -8726 314218 -2934 314454
rect -2698 314218 -2614 314454
rect -2378 314218 586302 314454
rect 586538 314218 586622 314454
rect 586858 314218 592650 314454
rect -8726 314134 592650 314218
rect -8726 313898 -2934 314134
rect -2698 313898 -2614 314134
rect -2378 313898 586302 314134
rect 586538 313898 586622 314134
rect 586858 313898 592650 314134
rect -8726 313866 592650 313898
rect -8726 308174 592650 308206
rect -8726 307938 -1974 308174
rect -1738 307938 -1654 308174
rect -1418 307938 585342 308174
rect 585578 307938 585662 308174
rect 585898 307938 592650 308174
rect -8726 307854 592650 307938
rect -8726 307618 -1974 307854
rect -1738 307618 -1654 307854
rect -1418 307618 585342 307854
rect 585578 307618 585662 307854
rect 585898 307618 592650 307854
rect -8726 307586 592650 307618
rect -8726 304454 592650 304486
rect -8726 304218 -2934 304454
rect -2698 304218 -2614 304454
rect -2378 304218 586302 304454
rect 586538 304218 586622 304454
rect 586858 304218 592650 304454
rect -8726 304134 592650 304218
rect -8726 303898 -2934 304134
rect -2698 303898 -2614 304134
rect -2378 303898 586302 304134
rect 586538 303898 586622 304134
rect 586858 303898 592650 304134
rect -8726 303866 592650 303898
rect -8726 298174 592650 298206
rect -8726 297938 -1974 298174
rect -1738 297938 -1654 298174
rect -1418 297938 585342 298174
rect 585578 297938 585662 298174
rect 585898 297938 592650 298174
rect -8726 297854 592650 297938
rect -8726 297618 -1974 297854
rect -1738 297618 -1654 297854
rect -1418 297618 585342 297854
rect 585578 297618 585662 297854
rect 585898 297618 592650 297854
rect -8726 297586 592650 297618
rect -8726 294454 592650 294486
rect -8726 294218 -2934 294454
rect -2698 294218 -2614 294454
rect -2378 294218 586302 294454
rect 586538 294218 586622 294454
rect 586858 294218 592650 294454
rect -8726 294134 592650 294218
rect -8726 293898 -2934 294134
rect -2698 293898 -2614 294134
rect -2378 293898 586302 294134
rect 586538 293898 586622 294134
rect 586858 293898 592650 294134
rect -8726 293866 592650 293898
rect -8726 288174 592650 288206
rect -8726 287938 -1974 288174
rect -1738 287938 -1654 288174
rect -1418 287938 585342 288174
rect 585578 287938 585662 288174
rect 585898 287938 592650 288174
rect -8726 287854 592650 287938
rect -8726 287618 -1974 287854
rect -1738 287618 -1654 287854
rect -1418 287618 585342 287854
rect 585578 287618 585662 287854
rect 585898 287618 592650 287854
rect -8726 287586 592650 287618
rect -8726 284454 592650 284486
rect -8726 284218 -2934 284454
rect -2698 284218 -2614 284454
rect -2378 284218 586302 284454
rect 586538 284218 586622 284454
rect 586858 284218 592650 284454
rect -8726 284134 592650 284218
rect -8726 283898 -2934 284134
rect -2698 283898 -2614 284134
rect -2378 283898 586302 284134
rect 586538 283898 586622 284134
rect 586858 283898 592650 284134
rect -8726 283866 592650 283898
rect -8726 278174 592650 278206
rect -8726 277938 -1974 278174
rect -1738 277938 -1654 278174
rect -1418 277938 585342 278174
rect 585578 277938 585662 278174
rect 585898 277938 592650 278174
rect -8726 277854 592650 277938
rect -8726 277618 -1974 277854
rect -1738 277618 -1654 277854
rect -1418 277618 585342 277854
rect 585578 277618 585662 277854
rect 585898 277618 592650 277854
rect -8726 277586 592650 277618
rect -8726 274454 592650 274486
rect -8726 274218 -2934 274454
rect -2698 274218 -2614 274454
rect -2378 274218 586302 274454
rect 586538 274218 586622 274454
rect 586858 274218 592650 274454
rect -8726 274134 592650 274218
rect -8726 273898 -2934 274134
rect -2698 273898 -2614 274134
rect -2378 273898 586302 274134
rect 586538 273898 586622 274134
rect 586858 273898 592650 274134
rect -8726 273866 592650 273898
rect -8726 268174 592650 268206
rect -8726 267938 -1974 268174
rect -1738 267938 -1654 268174
rect -1418 267938 585342 268174
rect 585578 267938 585662 268174
rect 585898 267938 592650 268174
rect -8726 267854 592650 267938
rect -8726 267618 -1974 267854
rect -1738 267618 -1654 267854
rect -1418 267618 585342 267854
rect 585578 267618 585662 267854
rect 585898 267618 592650 267854
rect -8726 267586 592650 267618
rect -8726 264454 592650 264486
rect -8726 264218 -2934 264454
rect -2698 264218 -2614 264454
rect -2378 264218 586302 264454
rect 586538 264218 586622 264454
rect 586858 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -2934 264134
rect -2698 263898 -2614 264134
rect -2378 263898 586302 264134
rect 586538 263898 586622 264134
rect 586858 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 258174 592650 258206
rect -8726 257938 -1974 258174
rect -1738 257938 -1654 258174
rect -1418 257938 585342 258174
rect 585578 257938 585662 258174
rect 585898 257938 592650 258174
rect -8726 257854 592650 257938
rect -8726 257618 -1974 257854
rect -1738 257618 -1654 257854
rect -1418 257618 585342 257854
rect 585578 257618 585662 257854
rect 585898 257618 592650 257854
rect -8726 257586 592650 257618
rect -8726 254454 592650 254486
rect -8726 254218 -2934 254454
rect -2698 254218 -2614 254454
rect -2378 254218 586302 254454
rect 586538 254218 586622 254454
rect 586858 254218 592650 254454
rect -8726 254134 592650 254218
rect -8726 253898 -2934 254134
rect -2698 253898 -2614 254134
rect -2378 253898 586302 254134
rect 586538 253898 586622 254134
rect 586858 253898 592650 254134
rect -8726 253866 592650 253898
rect -8726 248174 592650 248206
rect -8726 247938 -1974 248174
rect -1738 247938 -1654 248174
rect -1418 247938 585342 248174
rect 585578 247938 585662 248174
rect 585898 247938 592650 248174
rect -8726 247854 592650 247938
rect -8726 247618 -1974 247854
rect -1738 247618 -1654 247854
rect -1418 247618 585342 247854
rect 585578 247618 585662 247854
rect 585898 247618 592650 247854
rect -8726 247586 592650 247618
rect -8726 244454 592650 244486
rect -8726 244218 -2934 244454
rect -2698 244218 -2614 244454
rect -2378 244218 586302 244454
rect 586538 244218 586622 244454
rect 586858 244218 592650 244454
rect -8726 244134 592650 244218
rect -8726 243898 -2934 244134
rect -2698 243898 -2614 244134
rect -2378 243898 586302 244134
rect 586538 243898 586622 244134
rect 586858 243898 592650 244134
rect -8726 243866 592650 243898
rect -8726 238174 592650 238206
rect -8726 237938 -1974 238174
rect -1738 237938 -1654 238174
rect -1418 237938 585342 238174
rect 585578 237938 585662 238174
rect 585898 237938 592650 238174
rect -8726 237854 592650 237938
rect -8726 237618 -1974 237854
rect -1738 237618 -1654 237854
rect -1418 237618 585342 237854
rect 585578 237618 585662 237854
rect 585898 237618 592650 237854
rect -8726 237586 592650 237618
rect -8726 234454 592650 234486
rect -8726 234218 -2934 234454
rect -2698 234218 -2614 234454
rect -2378 234218 586302 234454
rect 586538 234218 586622 234454
rect 586858 234218 592650 234454
rect -8726 234134 592650 234218
rect -8726 233898 -2934 234134
rect -2698 233898 -2614 234134
rect -2378 233898 586302 234134
rect 586538 233898 586622 234134
rect 586858 233898 592650 234134
rect -8726 233866 592650 233898
rect -8726 228174 592650 228206
rect -8726 227938 -1974 228174
rect -1738 227938 -1654 228174
rect -1418 227938 585342 228174
rect 585578 227938 585662 228174
rect 585898 227938 592650 228174
rect -8726 227854 592650 227938
rect -8726 227618 -1974 227854
rect -1738 227618 -1654 227854
rect -1418 227618 585342 227854
rect 585578 227618 585662 227854
rect 585898 227618 592650 227854
rect -8726 227586 592650 227618
rect -8726 224454 592650 224486
rect -8726 224218 -2934 224454
rect -2698 224218 -2614 224454
rect -2378 224218 586302 224454
rect 586538 224218 586622 224454
rect 586858 224218 592650 224454
rect -8726 224134 592650 224218
rect -8726 223898 -2934 224134
rect -2698 223898 -2614 224134
rect -2378 223898 586302 224134
rect 586538 223898 586622 224134
rect 586858 223898 592650 224134
rect -8726 223866 592650 223898
rect -8726 218174 592650 218206
rect -8726 217938 -1974 218174
rect -1738 217938 -1654 218174
rect -1418 217938 585342 218174
rect 585578 217938 585662 218174
rect 585898 217938 592650 218174
rect -8726 217854 592650 217938
rect -8726 217618 -1974 217854
rect -1738 217618 -1654 217854
rect -1418 217618 585342 217854
rect 585578 217618 585662 217854
rect 585898 217618 592650 217854
rect -8726 217586 592650 217618
rect -8726 214454 592650 214486
rect -8726 214218 -2934 214454
rect -2698 214218 -2614 214454
rect -2378 214218 586302 214454
rect 586538 214218 586622 214454
rect 586858 214218 592650 214454
rect -8726 214134 592650 214218
rect -8726 213898 -2934 214134
rect -2698 213898 -2614 214134
rect -2378 213898 586302 214134
rect 586538 213898 586622 214134
rect 586858 213898 592650 214134
rect -8726 213866 592650 213898
rect -8726 208174 592650 208206
rect -8726 207938 -1974 208174
rect -1738 207938 -1654 208174
rect -1418 207938 14107 208174
rect 14343 207938 21949 208174
rect 22185 207938 29791 208174
rect 30027 207938 37633 208174
rect 37869 207938 48239 208174
rect 48475 207938 56081 208174
rect 56317 207938 63923 208174
rect 64159 207938 71765 208174
rect 72001 207938 82371 208174
rect 82607 207938 90213 208174
rect 90449 207938 98055 208174
rect 98291 207938 105897 208174
rect 106133 207938 116503 208174
rect 116739 207938 124345 208174
rect 124581 207938 132187 208174
rect 132423 207938 140029 208174
rect 140265 207938 150635 208174
rect 150871 207938 158477 208174
rect 158713 207938 166319 208174
rect 166555 207938 174161 208174
rect 174397 207938 184767 208174
rect 185003 207938 192609 208174
rect 192845 207938 200451 208174
rect 200687 207938 208293 208174
rect 208529 207938 218899 208174
rect 219135 207938 226741 208174
rect 226977 207938 234583 208174
rect 234819 207938 242425 208174
rect 242661 207938 253031 208174
rect 253267 207938 260873 208174
rect 261109 207938 268715 208174
rect 268951 207938 276557 208174
rect 276793 207938 307407 208174
rect 307643 207938 315249 208174
rect 315485 207938 323091 208174
rect 323327 207938 330933 208174
rect 331169 207938 341539 208174
rect 341775 207938 349381 208174
rect 349617 207938 357223 208174
rect 357459 207938 365065 208174
rect 365301 207938 375671 208174
rect 375907 207938 383513 208174
rect 383749 207938 391355 208174
rect 391591 207938 399197 208174
rect 399433 207938 409803 208174
rect 410039 207938 417645 208174
rect 417881 207938 425487 208174
rect 425723 207938 433329 208174
rect 433565 207938 443935 208174
rect 444171 207938 451777 208174
rect 452013 207938 459619 208174
rect 459855 207938 467461 208174
rect 467697 207938 478067 208174
rect 478303 207938 485909 208174
rect 486145 207938 493751 208174
rect 493987 207938 501593 208174
rect 501829 207938 512199 208174
rect 512435 207938 520041 208174
rect 520277 207938 527883 208174
rect 528119 207938 535725 208174
rect 535961 207938 546331 208174
rect 546567 207938 554173 208174
rect 554409 207938 562015 208174
rect 562251 207938 569857 208174
rect 570093 207938 585342 208174
rect 585578 207938 585662 208174
rect 585898 207938 592650 208174
rect -8726 207854 592650 207938
rect -8726 207618 -1974 207854
rect -1738 207618 -1654 207854
rect -1418 207618 14107 207854
rect 14343 207618 21949 207854
rect 22185 207618 29791 207854
rect 30027 207618 37633 207854
rect 37869 207618 48239 207854
rect 48475 207618 56081 207854
rect 56317 207618 63923 207854
rect 64159 207618 71765 207854
rect 72001 207618 82371 207854
rect 82607 207618 90213 207854
rect 90449 207618 98055 207854
rect 98291 207618 105897 207854
rect 106133 207618 116503 207854
rect 116739 207618 124345 207854
rect 124581 207618 132187 207854
rect 132423 207618 140029 207854
rect 140265 207618 150635 207854
rect 150871 207618 158477 207854
rect 158713 207618 166319 207854
rect 166555 207618 174161 207854
rect 174397 207618 184767 207854
rect 185003 207618 192609 207854
rect 192845 207618 200451 207854
rect 200687 207618 208293 207854
rect 208529 207618 218899 207854
rect 219135 207618 226741 207854
rect 226977 207618 234583 207854
rect 234819 207618 242425 207854
rect 242661 207618 253031 207854
rect 253267 207618 260873 207854
rect 261109 207618 268715 207854
rect 268951 207618 276557 207854
rect 276793 207618 307407 207854
rect 307643 207618 315249 207854
rect 315485 207618 323091 207854
rect 323327 207618 330933 207854
rect 331169 207618 341539 207854
rect 341775 207618 349381 207854
rect 349617 207618 357223 207854
rect 357459 207618 365065 207854
rect 365301 207618 375671 207854
rect 375907 207618 383513 207854
rect 383749 207618 391355 207854
rect 391591 207618 399197 207854
rect 399433 207618 409803 207854
rect 410039 207618 417645 207854
rect 417881 207618 425487 207854
rect 425723 207618 433329 207854
rect 433565 207618 443935 207854
rect 444171 207618 451777 207854
rect 452013 207618 459619 207854
rect 459855 207618 467461 207854
rect 467697 207618 478067 207854
rect 478303 207618 485909 207854
rect 486145 207618 493751 207854
rect 493987 207618 501593 207854
rect 501829 207618 512199 207854
rect 512435 207618 520041 207854
rect 520277 207618 527883 207854
rect 528119 207618 535725 207854
rect 535961 207618 546331 207854
rect 546567 207618 554173 207854
rect 554409 207618 562015 207854
rect 562251 207618 569857 207854
rect 570093 207618 585342 207854
rect 585578 207618 585662 207854
rect 585898 207618 592650 207854
rect -8726 207586 592650 207618
rect -8726 204454 592650 204486
rect -8726 204218 -2934 204454
rect -2698 204218 -2614 204454
rect -2378 204218 18028 204454
rect 18264 204218 25870 204454
rect 26106 204218 33712 204454
rect 33948 204218 41554 204454
rect 41790 204218 52160 204454
rect 52396 204218 60002 204454
rect 60238 204218 67844 204454
rect 68080 204218 75686 204454
rect 75922 204218 86292 204454
rect 86528 204218 94134 204454
rect 94370 204218 101976 204454
rect 102212 204218 109818 204454
rect 110054 204218 120424 204454
rect 120660 204218 128266 204454
rect 128502 204218 136108 204454
rect 136344 204218 143950 204454
rect 144186 204218 154556 204454
rect 154792 204218 162398 204454
rect 162634 204218 170240 204454
rect 170476 204218 178082 204454
rect 178318 204218 188688 204454
rect 188924 204218 196530 204454
rect 196766 204218 204372 204454
rect 204608 204218 212214 204454
rect 212450 204218 222820 204454
rect 223056 204218 230662 204454
rect 230898 204218 238504 204454
rect 238740 204218 246346 204454
rect 246582 204218 256952 204454
rect 257188 204218 264794 204454
rect 265030 204218 272636 204454
rect 272872 204218 280478 204454
rect 280714 204218 303486 204454
rect 303722 204218 311328 204454
rect 311564 204218 319170 204454
rect 319406 204218 327012 204454
rect 327248 204218 337618 204454
rect 337854 204218 345460 204454
rect 345696 204218 353302 204454
rect 353538 204218 361144 204454
rect 361380 204218 371750 204454
rect 371986 204218 379592 204454
rect 379828 204218 387434 204454
rect 387670 204218 395276 204454
rect 395512 204218 405882 204454
rect 406118 204218 413724 204454
rect 413960 204218 421566 204454
rect 421802 204218 429408 204454
rect 429644 204218 440014 204454
rect 440250 204218 447856 204454
rect 448092 204218 455698 204454
rect 455934 204218 463540 204454
rect 463776 204218 474146 204454
rect 474382 204218 481988 204454
rect 482224 204218 489830 204454
rect 490066 204218 497672 204454
rect 497908 204218 508278 204454
rect 508514 204218 516120 204454
rect 516356 204218 523962 204454
rect 524198 204218 531804 204454
rect 532040 204218 542410 204454
rect 542646 204218 550252 204454
rect 550488 204218 558094 204454
rect 558330 204218 565936 204454
rect 566172 204218 586302 204454
rect 586538 204218 586622 204454
rect 586858 204218 592650 204454
rect -8726 204134 592650 204218
rect -8726 203898 -2934 204134
rect -2698 203898 -2614 204134
rect -2378 203898 18028 204134
rect 18264 203898 25870 204134
rect 26106 203898 33712 204134
rect 33948 203898 41554 204134
rect 41790 203898 52160 204134
rect 52396 203898 60002 204134
rect 60238 203898 67844 204134
rect 68080 203898 75686 204134
rect 75922 203898 86292 204134
rect 86528 203898 94134 204134
rect 94370 203898 101976 204134
rect 102212 203898 109818 204134
rect 110054 203898 120424 204134
rect 120660 203898 128266 204134
rect 128502 203898 136108 204134
rect 136344 203898 143950 204134
rect 144186 203898 154556 204134
rect 154792 203898 162398 204134
rect 162634 203898 170240 204134
rect 170476 203898 178082 204134
rect 178318 203898 188688 204134
rect 188924 203898 196530 204134
rect 196766 203898 204372 204134
rect 204608 203898 212214 204134
rect 212450 203898 222820 204134
rect 223056 203898 230662 204134
rect 230898 203898 238504 204134
rect 238740 203898 246346 204134
rect 246582 203898 256952 204134
rect 257188 203898 264794 204134
rect 265030 203898 272636 204134
rect 272872 203898 280478 204134
rect 280714 203898 303486 204134
rect 303722 203898 311328 204134
rect 311564 203898 319170 204134
rect 319406 203898 327012 204134
rect 327248 203898 337618 204134
rect 337854 203898 345460 204134
rect 345696 203898 353302 204134
rect 353538 203898 361144 204134
rect 361380 203898 371750 204134
rect 371986 203898 379592 204134
rect 379828 203898 387434 204134
rect 387670 203898 395276 204134
rect 395512 203898 405882 204134
rect 406118 203898 413724 204134
rect 413960 203898 421566 204134
rect 421802 203898 429408 204134
rect 429644 203898 440014 204134
rect 440250 203898 447856 204134
rect 448092 203898 455698 204134
rect 455934 203898 463540 204134
rect 463776 203898 474146 204134
rect 474382 203898 481988 204134
rect 482224 203898 489830 204134
rect 490066 203898 497672 204134
rect 497908 203898 508278 204134
rect 508514 203898 516120 204134
rect 516356 203898 523962 204134
rect 524198 203898 531804 204134
rect 532040 203898 542410 204134
rect 542646 203898 550252 204134
rect 550488 203898 558094 204134
rect 558330 203898 565936 204134
rect 566172 203898 586302 204134
rect 586538 203898 586622 204134
rect 586858 203898 592650 204134
rect -8726 203866 592650 203898
rect -8726 198174 592650 198206
rect -8726 197938 -1974 198174
rect -1738 197938 -1654 198174
rect -1418 197938 14107 198174
rect 14343 197938 21949 198174
rect 22185 197938 29791 198174
rect 30027 197938 37633 198174
rect 37869 197938 48239 198174
rect 48475 197938 56081 198174
rect 56317 197938 63923 198174
rect 64159 197938 71765 198174
rect 72001 197938 82371 198174
rect 82607 197938 90213 198174
rect 90449 197938 98055 198174
rect 98291 197938 105897 198174
rect 106133 197938 116503 198174
rect 116739 197938 124345 198174
rect 124581 197938 132187 198174
rect 132423 197938 140029 198174
rect 140265 197938 150635 198174
rect 150871 197938 158477 198174
rect 158713 197938 166319 198174
rect 166555 197938 174161 198174
rect 174397 197938 184767 198174
rect 185003 197938 192609 198174
rect 192845 197938 200451 198174
rect 200687 197938 208293 198174
rect 208529 197938 218899 198174
rect 219135 197938 226741 198174
rect 226977 197938 234583 198174
rect 234819 197938 242425 198174
rect 242661 197938 253031 198174
rect 253267 197938 260873 198174
rect 261109 197938 268715 198174
rect 268951 197938 276557 198174
rect 276793 197938 307407 198174
rect 307643 197938 315249 198174
rect 315485 197938 323091 198174
rect 323327 197938 330933 198174
rect 331169 197938 341539 198174
rect 341775 197938 349381 198174
rect 349617 197938 357223 198174
rect 357459 197938 365065 198174
rect 365301 197938 375671 198174
rect 375907 197938 383513 198174
rect 383749 197938 391355 198174
rect 391591 197938 399197 198174
rect 399433 197938 409803 198174
rect 410039 197938 417645 198174
rect 417881 197938 425487 198174
rect 425723 197938 433329 198174
rect 433565 197938 443935 198174
rect 444171 197938 451777 198174
rect 452013 197938 459619 198174
rect 459855 197938 467461 198174
rect 467697 197938 478067 198174
rect 478303 197938 485909 198174
rect 486145 197938 493751 198174
rect 493987 197938 501593 198174
rect 501829 197938 512199 198174
rect 512435 197938 520041 198174
rect 520277 197938 527883 198174
rect 528119 197938 535725 198174
rect 535961 197938 546331 198174
rect 546567 197938 554173 198174
rect 554409 197938 562015 198174
rect 562251 197938 569857 198174
rect 570093 197938 585342 198174
rect 585578 197938 585662 198174
rect 585898 197938 592650 198174
rect -8726 197854 592650 197938
rect -8726 197618 -1974 197854
rect -1738 197618 -1654 197854
rect -1418 197618 14107 197854
rect 14343 197618 21949 197854
rect 22185 197618 29791 197854
rect 30027 197618 37633 197854
rect 37869 197618 48239 197854
rect 48475 197618 56081 197854
rect 56317 197618 63923 197854
rect 64159 197618 71765 197854
rect 72001 197618 82371 197854
rect 82607 197618 90213 197854
rect 90449 197618 98055 197854
rect 98291 197618 105897 197854
rect 106133 197618 116503 197854
rect 116739 197618 124345 197854
rect 124581 197618 132187 197854
rect 132423 197618 140029 197854
rect 140265 197618 150635 197854
rect 150871 197618 158477 197854
rect 158713 197618 166319 197854
rect 166555 197618 174161 197854
rect 174397 197618 184767 197854
rect 185003 197618 192609 197854
rect 192845 197618 200451 197854
rect 200687 197618 208293 197854
rect 208529 197618 218899 197854
rect 219135 197618 226741 197854
rect 226977 197618 234583 197854
rect 234819 197618 242425 197854
rect 242661 197618 253031 197854
rect 253267 197618 260873 197854
rect 261109 197618 268715 197854
rect 268951 197618 276557 197854
rect 276793 197618 307407 197854
rect 307643 197618 315249 197854
rect 315485 197618 323091 197854
rect 323327 197618 330933 197854
rect 331169 197618 341539 197854
rect 341775 197618 349381 197854
rect 349617 197618 357223 197854
rect 357459 197618 365065 197854
rect 365301 197618 375671 197854
rect 375907 197618 383513 197854
rect 383749 197618 391355 197854
rect 391591 197618 399197 197854
rect 399433 197618 409803 197854
rect 410039 197618 417645 197854
rect 417881 197618 425487 197854
rect 425723 197618 433329 197854
rect 433565 197618 443935 197854
rect 444171 197618 451777 197854
rect 452013 197618 459619 197854
rect 459855 197618 467461 197854
rect 467697 197618 478067 197854
rect 478303 197618 485909 197854
rect 486145 197618 493751 197854
rect 493987 197618 501593 197854
rect 501829 197618 512199 197854
rect 512435 197618 520041 197854
rect 520277 197618 527883 197854
rect 528119 197618 535725 197854
rect 535961 197618 546331 197854
rect 546567 197618 554173 197854
rect 554409 197618 562015 197854
rect 562251 197618 569857 197854
rect 570093 197618 585342 197854
rect 585578 197618 585662 197854
rect 585898 197618 592650 197854
rect -8726 197586 592650 197618
rect -8726 194454 592650 194486
rect -8726 194218 -2934 194454
rect -2698 194218 -2614 194454
rect -2378 194218 18028 194454
rect 18264 194218 25870 194454
rect 26106 194218 33712 194454
rect 33948 194218 41554 194454
rect 41790 194218 52160 194454
rect 52396 194218 60002 194454
rect 60238 194218 67844 194454
rect 68080 194218 75686 194454
rect 75922 194218 86292 194454
rect 86528 194218 94134 194454
rect 94370 194218 101976 194454
rect 102212 194218 109818 194454
rect 110054 194218 120424 194454
rect 120660 194218 128266 194454
rect 128502 194218 136108 194454
rect 136344 194218 143950 194454
rect 144186 194218 154556 194454
rect 154792 194218 162398 194454
rect 162634 194218 170240 194454
rect 170476 194218 178082 194454
rect 178318 194218 188688 194454
rect 188924 194218 196530 194454
rect 196766 194218 204372 194454
rect 204608 194218 212214 194454
rect 212450 194218 222820 194454
rect 223056 194218 230662 194454
rect 230898 194218 238504 194454
rect 238740 194218 246346 194454
rect 246582 194218 256952 194454
rect 257188 194218 264794 194454
rect 265030 194218 272636 194454
rect 272872 194218 280478 194454
rect 280714 194218 303486 194454
rect 303722 194218 311328 194454
rect 311564 194218 319170 194454
rect 319406 194218 327012 194454
rect 327248 194218 337618 194454
rect 337854 194218 345460 194454
rect 345696 194218 353302 194454
rect 353538 194218 361144 194454
rect 361380 194218 371750 194454
rect 371986 194218 379592 194454
rect 379828 194218 387434 194454
rect 387670 194218 395276 194454
rect 395512 194218 405882 194454
rect 406118 194218 413724 194454
rect 413960 194218 421566 194454
rect 421802 194218 429408 194454
rect 429644 194218 440014 194454
rect 440250 194218 447856 194454
rect 448092 194218 455698 194454
rect 455934 194218 463540 194454
rect 463776 194218 474146 194454
rect 474382 194218 481988 194454
rect 482224 194218 489830 194454
rect 490066 194218 497672 194454
rect 497908 194218 508278 194454
rect 508514 194218 516120 194454
rect 516356 194218 523962 194454
rect 524198 194218 531804 194454
rect 532040 194218 542410 194454
rect 542646 194218 550252 194454
rect 550488 194218 558094 194454
rect 558330 194218 565936 194454
rect 566172 194218 586302 194454
rect 586538 194218 586622 194454
rect 586858 194218 592650 194454
rect -8726 194134 592650 194218
rect -8726 193898 -2934 194134
rect -2698 193898 -2614 194134
rect -2378 193898 18028 194134
rect 18264 193898 25870 194134
rect 26106 193898 33712 194134
rect 33948 193898 41554 194134
rect 41790 193898 52160 194134
rect 52396 193898 60002 194134
rect 60238 193898 67844 194134
rect 68080 193898 75686 194134
rect 75922 193898 86292 194134
rect 86528 193898 94134 194134
rect 94370 193898 101976 194134
rect 102212 193898 109818 194134
rect 110054 193898 120424 194134
rect 120660 193898 128266 194134
rect 128502 193898 136108 194134
rect 136344 193898 143950 194134
rect 144186 193898 154556 194134
rect 154792 193898 162398 194134
rect 162634 193898 170240 194134
rect 170476 193898 178082 194134
rect 178318 193898 188688 194134
rect 188924 193898 196530 194134
rect 196766 193898 204372 194134
rect 204608 193898 212214 194134
rect 212450 193898 222820 194134
rect 223056 193898 230662 194134
rect 230898 193898 238504 194134
rect 238740 193898 246346 194134
rect 246582 193898 256952 194134
rect 257188 193898 264794 194134
rect 265030 193898 272636 194134
rect 272872 193898 280478 194134
rect 280714 193898 303486 194134
rect 303722 193898 311328 194134
rect 311564 193898 319170 194134
rect 319406 193898 327012 194134
rect 327248 193898 337618 194134
rect 337854 193898 345460 194134
rect 345696 193898 353302 194134
rect 353538 193898 361144 194134
rect 361380 193898 371750 194134
rect 371986 193898 379592 194134
rect 379828 193898 387434 194134
rect 387670 193898 395276 194134
rect 395512 193898 405882 194134
rect 406118 193898 413724 194134
rect 413960 193898 421566 194134
rect 421802 193898 429408 194134
rect 429644 193898 440014 194134
rect 440250 193898 447856 194134
rect 448092 193898 455698 194134
rect 455934 193898 463540 194134
rect 463776 193898 474146 194134
rect 474382 193898 481988 194134
rect 482224 193898 489830 194134
rect 490066 193898 497672 194134
rect 497908 193898 508278 194134
rect 508514 193898 516120 194134
rect 516356 193898 523962 194134
rect 524198 193898 531804 194134
rect 532040 193898 542410 194134
rect 542646 193898 550252 194134
rect 550488 193898 558094 194134
rect 558330 193898 565936 194134
rect 566172 193898 586302 194134
rect 586538 193898 586622 194134
rect 586858 193898 592650 194134
rect -8726 193866 592650 193898
rect -8726 188174 592650 188206
rect -8726 187938 -1974 188174
rect -1738 187938 -1654 188174
rect -1418 187938 43984 188174
rect 44220 187938 111581 188174
rect 111817 187938 179178 188174
rect 179414 187938 246775 188174
rect 247011 187938 337189 188174
rect 337425 187938 404786 188174
rect 405022 187938 472383 188174
rect 472619 187938 539980 188174
rect 540216 187938 585342 188174
rect 585578 187938 585662 188174
rect 585898 187938 592650 188174
rect -8726 187854 592650 187938
rect -8726 187618 -1974 187854
rect -1738 187618 -1654 187854
rect -1418 187618 43984 187854
rect 44220 187618 111581 187854
rect 111817 187618 179178 187854
rect 179414 187618 246775 187854
rect 247011 187618 337189 187854
rect 337425 187618 404786 187854
rect 405022 187618 472383 187854
rect 472619 187618 539980 187854
rect 540216 187618 585342 187854
rect 585578 187618 585662 187854
rect 585898 187618 592650 187854
rect -8726 187586 592650 187618
rect -8726 184454 592650 184486
rect -8726 184218 -2934 184454
rect -2698 184218 -2614 184454
rect -2378 184218 77782 184454
rect 78018 184218 145379 184454
rect 145615 184218 212976 184454
rect 213212 184218 280573 184454
rect 280809 184218 303391 184454
rect 303627 184218 370988 184454
rect 371224 184218 438585 184454
rect 438821 184218 506182 184454
rect 506418 184218 586302 184454
rect 586538 184218 586622 184454
rect 586858 184218 592650 184454
rect -8726 184134 592650 184218
rect -8726 183898 -2934 184134
rect -2698 183898 -2614 184134
rect -2378 183898 77782 184134
rect 78018 183898 145379 184134
rect 145615 183898 212976 184134
rect 213212 183898 280573 184134
rect 280809 183898 303391 184134
rect 303627 183898 370988 184134
rect 371224 183898 438585 184134
rect 438821 183898 506182 184134
rect 506418 183898 586302 184134
rect 586538 183898 586622 184134
rect 586858 183898 592650 184134
rect -8726 183866 592650 183898
rect -8726 178174 592650 178206
rect -8726 177938 -1974 178174
rect -1738 177938 -1654 178174
rect -1418 177938 585342 178174
rect 585578 177938 585662 178174
rect 585898 177938 592650 178174
rect -8726 177879 592650 177938
rect -8726 177854 14107 177879
rect -8726 177618 -1974 177854
rect -1738 177618 -1654 177854
rect -1418 177643 14107 177854
rect 14343 177643 21949 177879
rect 22185 177643 29791 177879
rect 30027 177643 37633 177879
rect 37869 177643 48239 177879
rect 48475 177643 56081 177879
rect 56317 177643 63923 177879
rect 64159 177643 71765 177879
rect 72001 177643 82371 177879
rect 82607 177643 90213 177879
rect 90449 177643 98055 177879
rect 98291 177643 105897 177879
rect 106133 177643 116503 177879
rect 116739 177643 124345 177879
rect 124581 177643 132187 177879
rect 132423 177643 140029 177879
rect 140265 177643 150635 177879
rect 150871 177643 158477 177879
rect 158713 177643 166319 177879
rect 166555 177643 174161 177879
rect 174397 177643 184767 177879
rect 185003 177643 192609 177879
rect 192845 177643 200451 177879
rect 200687 177643 208293 177879
rect 208529 177643 218899 177879
rect 219135 177643 226741 177879
rect 226977 177643 234583 177879
rect 234819 177643 242425 177879
rect 242661 177643 253031 177879
rect 253267 177643 260873 177879
rect 261109 177643 268715 177879
rect 268951 177643 276557 177879
rect 276793 177643 307407 177879
rect 307643 177643 315249 177879
rect 315485 177643 323091 177879
rect 323327 177643 330933 177879
rect 331169 177643 341539 177879
rect 341775 177643 349381 177879
rect 349617 177643 357223 177879
rect 357459 177643 365065 177879
rect 365301 177643 375671 177879
rect 375907 177643 383513 177879
rect 383749 177643 391355 177879
rect 391591 177643 399197 177879
rect 399433 177643 409803 177879
rect 410039 177643 417645 177879
rect 417881 177643 425487 177879
rect 425723 177643 433329 177879
rect 433565 177643 443935 177879
rect 444171 177643 451777 177879
rect 452013 177643 459619 177879
rect 459855 177643 467461 177879
rect 467697 177643 478067 177879
rect 478303 177643 485909 177879
rect 486145 177643 493751 177879
rect 493987 177643 501593 177879
rect 501829 177643 512199 177879
rect 512435 177643 520041 177879
rect 520277 177643 527883 177879
rect 528119 177643 535725 177879
rect 535961 177643 546331 177879
rect 546567 177643 554173 177879
rect 554409 177643 562015 177879
rect 562251 177643 569857 177879
rect 570093 177854 592650 177879
rect 570093 177643 585342 177854
rect -1418 177618 585342 177643
rect 585578 177618 585662 177854
rect 585898 177618 592650 177854
rect -8726 177586 592650 177618
rect -8726 174454 592650 174486
rect -8726 174218 -2934 174454
rect -2698 174218 -2614 174454
rect -2378 174218 18028 174454
rect 18264 174218 25870 174454
rect 26106 174218 33712 174454
rect 33948 174218 41554 174454
rect 41790 174218 52160 174454
rect 52396 174218 60002 174454
rect 60238 174218 67844 174454
rect 68080 174218 75686 174454
rect 75922 174218 86292 174454
rect 86528 174218 94134 174454
rect 94370 174218 101976 174454
rect 102212 174218 109818 174454
rect 110054 174218 120424 174454
rect 120660 174218 128266 174454
rect 128502 174218 136108 174454
rect 136344 174218 143950 174454
rect 144186 174218 154556 174454
rect 154792 174218 162398 174454
rect 162634 174218 170240 174454
rect 170476 174218 178082 174454
rect 178318 174218 188688 174454
rect 188924 174218 196530 174454
rect 196766 174218 204372 174454
rect 204608 174218 212214 174454
rect 212450 174218 222820 174454
rect 223056 174218 230662 174454
rect 230898 174218 238504 174454
rect 238740 174218 246346 174454
rect 246582 174218 256952 174454
rect 257188 174218 264794 174454
rect 265030 174218 272636 174454
rect 272872 174218 280478 174454
rect 280714 174218 303486 174454
rect 303722 174218 311328 174454
rect 311564 174218 319170 174454
rect 319406 174218 327012 174454
rect 327248 174218 337618 174454
rect 337854 174218 345460 174454
rect 345696 174218 353302 174454
rect 353538 174218 361144 174454
rect 361380 174218 371750 174454
rect 371986 174218 379592 174454
rect 379828 174218 387434 174454
rect 387670 174218 395276 174454
rect 395512 174218 405882 174454
rect 406118 174218 413724 174454
rect 413960 174218 421566 174454
rect 421802 174218 429408 174454
rect 429644 174218 440014 174454
rect 440250 174218 447856 174454
rect 448092 174218 455698 174454
rect 455934 174218 463540 174454
rect 463776 174218 474146 174454
rect 474382 174218 481988 174454
rect 482224 174218 489830 174454
rect 490066 174218 497672 174454
rect 497908 174218 508278 174454
rect 508514 174218 516120 174454
rect 516356 174218 523962 174454
rect 524198 174218 531804 174454
rect 532040 174218 542410 174454
rect 542646 174218 550252 174454
rect 550488 174218 558094 174454
rect 558330 174218 565936 174454
rect 566172 174218 586302 174454
rect 586538 174218 586622 174454
rect 586858 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -2934 174134
rect -2698 173898 -2614 174134
rect -2378 173898 18028 174134
rect 18264 173898 25870 174134
rect 26106 173898 33712 174134
rect 33948 173898 41554 174134
rect 41790 173898 52160 174134
rect 52396 173898 60002 174134
rect 60238 173898 67844 174134
rect 68080 173898 75686 174134
rect 75922 173898 86292 174134
rect 86528 173898 94134 174134
rect 94370 173898 101976 174134
rect 102212 173898 109818 174134
rect 110054 173898 120424 174134
rect 120660 173898 128266 174134
rect 128502 173898 136108 174134
rect 136344 173898 143950 174134
rect 144186 173898 154556 174134
rect 154792 173898 162398 174134
rect 162634 173898 170240 174134
rect 170476 173898 178082 174134
rect 178318 173898 188688 174134
rect 188924 173898 196530 174134
rect 196766 173898 204372 174134
rect 204608 173898 212214 174134
rect 212450 173898 222820 174134
rect 223056 173898 230662 174134
rect 230898 173898 238504 174134
rect 238740 173898 246346 174134
rect 246582 173898 256952 174134
rect 257188 173898 264794 174134
rect 265030 173898 272636 174134
rect 272872 173898 280478 174134
rect 280714 173898 303486 174134
rect 303722 173898 311328 174134
rect 311564 173898 319170 174134
rect 319406 173898 327012 174134
rect 327248 173898 337618 174134
rect 337854 173898 345460 174134
rect 345696 173898 353302 174134
rect 353538 173898 361144 174134
rect 361380 173898 371750 174134
rect 371986 173898 379592 174134
rect 379828 173898 387434 174134
rect 387670 173898 395276 174134
rect 395512 173898 405882 174134
rect 406118 173898 413724 174134
rect 413960 173898 421566 174134
rect 421802 173898 429408 174134
rect 429644 173898 440014 174134
rect 440250 173898 447856 174134
rect 448092 173898 455698 174134
rect 455934 173898 463540 174134
rect 463776 173898 474146 174134
rect 474382 173898 481988 174134
rect 482224 173898 489830 174134
rect 490066 173898 497672 174134
rect 497908 173898 508278 174134
rect 508514 173898 516120 174134
rect 516356 173898 523962 174134
rect 524198 173898 531804 174134
rect 532040 173898 542410 174134
rect 542646 173898 550252 174134
rect 550488 173898 558094 174134
rect 558330 173898 565936 174134
rect 566172 173898 586302 174134
rect 586538 173898 586622 174134
rect 586858 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 168174 592650 168206
rect -8726 167938 -1974 168174
rect -1738 167938 -1654 168174
rect -1418 167938 14107 168174
rect 14343 167938 21949 168174
rect 22185 167938 29791 168174
rect 30027 167938 37633 168174
rect 37869 167938 48239 168174
rect 48475 167938 56081 168174
rect 56317 167938 63923 168174
rect 64159 167938 71765 168174
rect 72001 167938 82371 168174
rect 82607 167938 90213 168174
rect 90449 167938 98055 168174
rect 98291 167938 105897 168174
rect 106133 167938 116503 168174
rect 116739 167938 124345 168174
rect 124581 167938 132187 168174
rect 132423 167938 140029 168174
rect 140265 167938 150635 168174
rect 150871 167938 158477 168174
rect 158713 167938 166319 168174
rect 166555 167938 174161 168174
rect 174397 167938 184767 168174
rect 185003 167938 192609 168174
rect 192845 167938 200451 168174
rect 200687 167938 208293 168174
rect 208529 167938 218899 168174
rect 219135 167938 226741 168174
rect 226977 167938 234583 168174
rect 234819 167938 242425 168174
rect 242661 167938 253031 168174
rect 253267 167938 260873 168174
rect 261109 167938 268715 168174
rect 268951 167938 276557 168174
rect 276793 167938 307407 168174
rect 307643 167938 315249 168174
rect 315485 167938 323091 168174
rect 323327 167938 330933 168174
rect 331169 167938 341539 168174
rect 341775 167938 349381 168174
rect 349617 167938 357223 168174
rect 357459 167938 365065 168174
rect 365301 167938 375671 168174
rect 375907 167938 383513 168174
rect 383749 167938 391355 168174
rect 391591 167938 399197 168174
rect 399433 167938 409803 168174
rect 410039 167938 417645 168174
rect 417881 167938 425487 168174
rect 425723 167938 433329 168174
rect 433565 167938 443935 168174
rect 444171 167938 451777 168174
rect 452013 167938 459619 168174
rect 459855 167938 467461 168174
rect 467697 167938 478067 168174
rect 478303 167938 485909 168174
rect 486145 167938 493751 168174
rect 493987 167938 501593 168174
rect 501829 167938 512199 168174
rect 512435 167938 520041 168174
rect 520277 167938 527883 168174
rect 528119 167938 535725 168174
rect 535961 167938 546331 168174
rect 546567 167938 554173 168174
rect 554409 167938 562015 168174
rect 562251 167938 569857 168174
rect 570093 167938 585342 168174
rect 585578 167938 585662 168174
rect 585898 167938 592650 168174
rect -8726 167854 592650 167938
rect -8726 167618 -1974 167854
rect -1738 167618 -1654 167854
rect -1418 167618 14107 167854
rect 14343 167618 21949 167854
rect 22185 167618 29791 167854
rect 30027 167618 37633 167854
rect 37869 167618 48239 167854
rect 48475 167618 56081 167854
rect 56317 167618 63923 167854
rect 64159 167618 71765 167854
rect 72001 167618 82371 167854
rect 82607 167618 90213 167854
rect 90449 167618 98055 167854
rect 98291 167618 105897 167854
rect 106133 167618 116503 167854
rect 116739 167618 124345 167854
rect 124581 167618 132187 167854
rect 132423 167618 140029 167854
rect 140265 167618 150635 167854
rect 150871 167618 158477 167854
rect 158713 167618 166319 167854
rect 166555 167618 174161 167854
rect 174397 167618 184767 167854
rect 185003 167618 192609 167854
rect 192845 167618 200451 167854
rect 200687 167618 208293 167854
rect 208529 167618 218899 167854
rect 219135 167618 226741 167854
rect 226977 167618 234583 167854
rect 234819 167618 242425 167854
rect 242661 167618 253031 167854
rect 253267 167618 260873 167854
rect 261109 167618 268715 167854
rect 268951 167618 276557 167854
rect 276793 167618 307407 167854
rect 307643 167618 315249 167854
rect 315485 167618 323091 167854
rect 323327 167618 330933 167854
rect 331169 167618 341539 167854
rect 341775 167618 349381 167854
rect 349617 167618 357223 167854
rect 357459 167618 365065 167854
rect 365301 167618 375671 167854
rect 375907 167618 383513 167854
rect 383749 167618 391355 167854
rect 391591 167618 399197 167854
rect 399433 167618 409803 167854
rect 410039 167618 417645 167854
rect 417881 167618 425487 167854
rect 425723 167618 433329 167854
rect 433565 167618 443935 167854
rect 444171 167618 451777 167854
rect 452013 167618 459619 167854
rect 459855 167618 467461 167854
rect 467697 167618 478067 167854
rect 478303 167618 485909 167854
rect 486145 167618 493751 167854
rect 493987 167618 501593 167854
rect 501829 167618 512199 167854
rect 512435 167618 520041 167854
rect 520277 167618 527883 167854
rect 528119 167618 535725 167854
rect 535961 167618 546331 167854
rect 546567 167618 554173 167854
rect 554409 167618 562015 167854
rect 562251 167618 569857 167854
rect 570093 167618 585342 167854
rect 585578 167618 585662 167854
rect 585898 167618 592650 167854
rect -8726 167586 592650 167618
rect -8726 164454 592650 164486
rect -8726 164218 -2934 164454
rect -2698 164218 -2614 164454
rect -2378 164218 18028 164454
rect 18264 164218 25870 164454
rect 26106 164218 33712 164454
rect 33948 164218 41554 164454
rect 41790 164218 52160 164454
rect 52396 164218 60002 164454
rect 60238 164218 67844 164454
rect 68080 164218 75686 164454
rect 75922 164218 86292 164454
rect 86528 164218 94134 164454
rect 94370 164218 101976 164454
rect 102212 164218 109818 164454
rect 110054 164218 120424 164454
rect 120660 164218 128266 164454
rect 128502 164218 136108 164454
rect 136344 164218 143950 164454
rect 144186 164218 154556 164454
rect 154792 164218 162398 164454
rect 162634 164218 170240 164454
rect 170476 164218 178082 164454
rect 178318 164218 188688 164454
rect 188924 164218 196530 164454
rect 196766 164218 204372 164454
rect 204608 164218 212214 164454
rect 212450 164218 222820 164454
rect 223056 164218 230662 164454
rect 230898 164218 238504 164454
rect 238740 164218 246346 164454
rect 246582 164218 256952 164454
rect 257188 164218 264794 164454
rect 265030 164218 272636 164454
rect 272872 164218 280478 164454
rect 280714 164218 303486 164454
rect 303722 164218 311328 164454
rect 311564 164218 319170 164454
rect 319406 164218 327012 164454
rect 327248 164218 337618 164454
rect 337854 164218 345460 164454
rect 345696 164218 353302 164454
rect 353538 164218 361144 164454
rect 361380 164218 371750 164454
rect 371986 164218 379592 164454
rect 379828 164218 387434 164454
rect 387670 164218 395276 164454
rect 395512 164218 405882 164454
rect 406118 164218 413724 164454
rect 413960 164218 421566 164454
rect 421802 164218 429408 164454
rect 429644 164218 440014 164454
rect 440250 164218 447856 164454
rect 448092 164218 455698 164454
rect 455934 164218 463540 164454
rect 463776 164218 474146 164454
rect 474382 164218 481988 164454
rect 482224 164218 489830 164454
rect 490066 164218 497672 164454
rect 497908 164218 508278 164454
rect 508514 164218 516120 164454
rect 516356 164218 523962 164454
rect 524198 164218 531804 164454
rect 532040 164218 542410 164454
rect 542646 164218 550252 164454
rect 550488 164218 558094 164454
rect 558330 164218 565936 164454
rect 566172 164218 586302 164454
rect 586538 164218 586622 164454
rect 586858 164218 592650 164454
rect -8726 164134 592650 164218
rect -8726 163898 -2934 164134
rect -2698 163898 -2614 164134
rect -2378 163898 18028 164134
rect 18264 163898 25870 164134
rect 26106 163898 33712 164134
rect 33948 163898 41554 164134
rect 41790 163898 52160 164134
rect 52396 163898 60002 164134
rect 60238 163898 67844 164134
rect 68080 163898 75686 164134
rect 75922 163898 86292 164134
rect 86528 163898 94134 164134
rect 94370 163898 101976 164134
rect 102212 163898 109818 164134
rect 110054 163898 120424 164134
rect 120660 163898 128266 164134
rect 128502 163898 136108 164134
rect 136344 163898 143950 164134
rect 144186 163898 154556 164134
rect 154792 163898 162398 164134
rect 162634 163898 170240 164134
rect 170476 163898 178082 164134
rect 178318 163898 188688 164134
rect 188924 163898 196530 164134
rect 196766 163898 204372 164134
rect 204608 163898 212214 164134
rect 212450 163898 222820 164134
rect 223056 163898 230662 164134
rect 230898 163898 238504 164134
rect 238740 163898 246346 164134
rect 246582 163898 256952 164134
rect 257188 163898 264794 164134
rect 265030 163898 272636 164134
rect 272872 163898 280478 164134
rect 280714 163898 303486 164134
rect 303722 163898 311328 164134
rect 311564 163898 319170 164134
rect 319406 163898 327012 164134
rect 327248 163898 337618 164134
rect 337854 163898 345460 164134
rect 345696 163898 353302 164134
rect 353538 163898 361144 164134
rect 361380 163898 371750 164134
rect 371986 163898 379592 164134
rect 379828 163898 387434 164134
rect 387670 163898 395276 164134
rect 395512 163898 405882 164134
rect 406118 163898 413724 164134
rect 413960 163898 421566 164134
rect 421802 163898 429408 164134
rect 429644 163898 440014 164134
rect 440250 163898 447856 164134
rect 448092 163898 455698 164134
rect 455934 163898 463540 164134
rect 463776 163898 474146 164134
rect 474382 163898 481988 164134
rect 482224 163898 489830 164134
rect 490066 163898 497672 164134
rect 497908 163898 508278 164134
rect 508514 163898 516120 164134
rect 516356 163898 523962 164134
rect 524198 163898 531804 164134
rect 532040 163898 542410 164134
rect 542646 163898 550252 164134
rect 550488 163898 558094 164134
rect 558330 163898 565936 164134
rect 566172 163898 586302 164134
rect 586538 163898 586622 164134
rect 586858 163898 592650 164134
rect -8726 163866 592650 163898
rect -8726 158174 592650 158206
rect -8726 157938 -1974 158174
rect -1738 157938 -1654 158174
rect -1418 157938 585342 158174
rect 585578 157938 585662 158174
rect 585898 157938 592650 158174
rect -8726 157854 592650 157938
rect -8726 157618 -1974 157854
rect -1738 157618 -1654 157854
rect -1418 157618 585342 157854
rect 585578 157618 585662 157854
rect 585898 157618 592650 157854
rect -8726 157586 592650 157618
rect -8726 154454 592650 154486
rect -8726 154218 -2934 154454
rect -2698 154218 -2614 154454
rect -2378 154218 586302 154454
rect 586538 154218 586622 154454
rect 586858 154218 592650 154454
rect -8726 154134 592650 154218
rect -8726 153898 -2934 154134
rect -2698 153898 -2614 154134
rect -2378 153898 586302 154134
rect 586538 153898 586622 154134
rect 586858 153898 592650 154134
rect -8726 153866 592650 153898
rect -8726 148174 592650 148206
rect -8726 147938 -1974 148174
rect -1738 147938 -1654 148174
rect -1418 147938 585342 148174
rect 585578 147938 585662 148174
rect 585898 147938 592650 148174
rect -8726 147854 592650 147938
rect -8726 147618 -1974 147854
rect -1738 147618 -1654 147854
rect -1418 147618 585342 147854
rect 585578 147618 585662 147854
rect 585898 147618 592650 147854
rect -8726 147586 592650 147618
rect -8726 144454 592650 144486
rect -8726 144218 -2934 144454
rect -2698 144218 -2614 144454
rect -2378 144218 586302 144454
rect 586538 144218 586622 144454
rect 586858 144218 592650 144454
rect -8726 144134 592650 144218
rect -8726 143898 -2934 144134
rect -2698 143898 -2614 144134
rect -2378 143898 586302 144134
rect 586538 143898 586622 144134
rect 586858 143898 592650 144134
rect -8726 143866 592650 143898
rect -8726 138174 592650 138206
rect -8726 137938 -1974 138174
rect -1738 137938 -1654 138174
rect -1418 137938 585342 138174
rect 585578 137938 585662 138174
rect 585898 137938 592650 138174
rect -8726 137854 592650 137938
rect -8726 137618 -1974 137854
rect -1738 137618 -1654 137854
rect -1418 137618 585342 137854
rect 585578 137618 585662 137854
rect 585898 137618 592650 137854
rect -8726 137586 592650 137618
rect -8726 134454 592650 134486
rect -8726 134218 -2934 134454
rect -2698 134218 -2614 134454
rect -2378 134218 586302 134454
rect 586538 134218 586622 134454
rect 586858 134218 592650 134454
rect -8726 134134 592650 134218
rect -8726 133898 -2934 134134
rect -2698 133898 -2614 134134
rect -2378 133898 586302 134134
rect 586538 133898 586622 134134
rect 586858 133898 592650 134134
rect -8726 133866 592650 133898
rect -8726 128174 592650 128206
rect -8726 127938 -1974 128174
rect -1738 127938 -1654 128174
rect -1418 127938 585342 128174
rect 585578 127938 585662 128174
rect 585898 127938 592650 128174
rect -8726 127854 592650 127938
rect -8726 127618 -1974 127854
rect -1738 127618 -1654 127854
rect -1418 127618 585342 127854
rect 585578 127618 585662 127854
rect 585898 127618 592650 127854
rect -8726 127586 592650 127618
rect -8726 124454 592650 124486
rect -8726 124218 -2934 124454
rect -2698 124218 -2614 124454
rect -2378 124218 586302 124454
rect 586538 124218 586622 124454
rect 586858 124218 592650 124454
rect -8726 124134 592650 124218
rect -8726 123898 -2934 124134
rect -2698 123898 -2614 124134
rect -2378 123898 586302 124134
rect 586538 123898 586622 124134
rect 586858 123898 592650 124134
rect -8726 123866 592650 123898
rect -8726 118174 592650 118206
rect -8726 117938 -1974 118174
rect -1738 117938 -1654 118174
rect -1418 117938 585342 118174
rect 585578 117938 585662 118174
rect 585898 117938 592650 118174
rect -8726 117854 592650 117938
rect -8726 117618 -1974 117854
rect -1738 117618 -1654 117854
rect -1418 117618 585342 117854
rect 585578 117618 585662 117854
rect 585898 117618 592650 117854
rect -8726 117586 592650 117618
rect -8726 114454 592650 114486
rect -8726 114218 -2934 114454
rect -2698 114218 -2614 114454
rect -2378 114218 586302 114454
rect 586538 114218 586622 114454
rect 586858 114218 592650 114454
rect -8726 114134 592650 114218
rect -8726 113898 -2934 114134
rect -2698 113898 -2614 114134
rect -2378 113898 586302 114134
rect 586538 113898 586622 114134
rect 586858 113898 592650 114134
rect -8726 113866 592650 113898
rect -8726 108174 592650 108206
rect -8726 107938 -1974 108174
rect -1738 107938 -1654 108174
rect -1418 107938 585342 108174
rect 585578 107938 585662 108174
rect 585898 107938 592650 108174
rect -8726 107854 592650 107938
rect -8726 107618 -1974 107854
rect -1738 107618 -1654 107854
rect -1418 107618 585342 107854
rect 585578 107618 585662 107854
rect 585898 107618 592650 107854
rect -8726 107586 592650 107618
rect -8726 104454 592650 104486
rect -8726 104218 -2934 104454
rect -2698 104218 -2614 104454
rect -2378 104218 586302 104454
rect 586538 104218 586622 104454
rect 586858 104218 592650 104454
rect -8726 104134 592650 104218
rect -8726 103898 -2934 104134
rect -2698 103898 -2614 104134
rect -2378 103898 586302 104134
rect 586538 103898 586622 104134
rect 586858 103898 592650 104134
rect -8726 103866 592650 103898
rect -8726 98174 592650 98206
rect -8726 97938 -1974 98174
rect -1738 97938 -1654 98174
rect -1418 97938 585342 98174
rect 585578 97938 585662 98174
rect 585898 97938 592650 98174
rect -8726 97854 592650 97938
rect -8726 97618 -1974 97854
rect -1738 97618 -1654 97854
rect -1418 97618 585342 97854
rect 585578 97618 585662 97854
rect 585898 97618 592650 97854
rect -8726 97586 592650 97618
rect -8726 94454 592650 94486
rect -8726 94218 -2934 94454
rect -2698 94218 -2614 94454
rect -2378 94218 586302 94454
rect 586538 94218 586622 94454
rect 586858 94218 592650 94454
rect -8726 94134 592650 94218
rect -8726 93898 -2934 94134
rect -2698 93898 -2614 94134
rect -2378 93898 586302 94134
rect 586538 93898 586622 94134
rect 586858 93898 592650 94134
rect -8726 93866 592650 93898
rect -8726 88174 592650 88206
rect -8726 87938 -1974 88174
rect -1738 87938 -1654 88174
rect -1418 87938 585342 88174
rect 585578 87938 585662 88174
rect 585898 87938 592650 88174
rect -8726 87854 592650 87938
rect -8726 87618 -1974 87854
rect -1738 87618 -1654 87854
rect -1418 87618 585342 87854
rect 585578 87618 585662 87854
rect 585898 87618 592650 87854
rect -8726 87586 592650 87618
rect -8726 84454 592650 84486
rect -8726 84218 -2934 84454
rect -2698 84218 -2614 84454
rect -2378 84218 586302 84454
rect 586538 84218 586622 84454
rect 586858 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -2934 84134
rect -2698 83898 -2614 84134
rect -2378 83898 586302 84134
rect 586538 83898 586622 84134
rect 586858 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 78174 592650 78206
rect -8726 77938 -1974 78174
rect -1738 77938 -1654 78174
rect -1418 77938 585342 78174
rect 585578 77938 585662 78174
rect 585898 77938 592650 78174
rect -8726 77854 592650 77938
rect -8726 77618 -1974 77854
rect -1738 77618 -1654 77854
rect -1418 77618 585342 77854
rect 585578 77618 585662 77854
rect 585898 77618 592650 77854
rect -8726 77586 592650 77618
rect -8726 74454 592650 74486
rect -8726 74218 -2934 74454
rect -2698 74218 -2614 74454
rect -2378 74218 586302 74454
rect 586538 74218 586622 74454
rect 586858 74218 592650 74454
rect -8726 74134 592650 74218
rect -8726 73898 -2934 74134
rect -2698 73898 -2614 74134
rect -2378 73898 586302 74134
rect 586538 73898 586622 74134
rect 586858 73898 592650 74134
rect -8726 73866 592650 73898
rect -8726 68174 592650 68206
rect -8726 67938 -1974 68174
rect -1738 67938 -1654 68174
rect -1418 67938 585342 68174
rect 585578 67938 585662 68174
rect 585898 67938 592650 68174
rect -8726 67854 592650 67938
rect -8726 67618 -1974 67854
rect -1738 67618 -1654 67854
rect -1418 67618 585342 67854
rect 585578 67618 585662 67854
rect 585898 67618 592650 67854
rect -8726 67586 592650 67618
rect -8726 64454 592650 64486
rect -8726 64218 -2934 64454
rect -2698 64218 -2614 64454
rect -2378 64218 586302 64454
rect 586538 64218 586622 64454
rect 586858 64218 592650 64454
rect -8726 64171 592650 64218
rect -8726 64134 293034 64171
rect -8726 63898 -2934 64134
rect -2698 63898 -2614 64134
rect -2378 63935 293034 64134
rect 293270 64134 592650 64171
rect 293270 63935 586302 64134
rect -2378 63898 586302 63935
rect 586538 63898 586622 64134
rect 586858 63898 592650 64134
rect -8726 63866 592650 63898
rect -8726 58174 592650 58206
rect -8726 57938 -1974 58174
rect -1738 57938 -1654 58174
rect -1418 57938 277674 58174
rect 277910 57938 308394 58174
rect 308630 57938 585342 58174
rect 585578 57938 585662 58174
rect 585898 57938 592650 58174
rect -8726 57854 592650 57938
rect -8726 57618 -1974 57854
rect -1738 57618 -1654 57854
rect -1418 57618 277674 57854
rect 277910 57618 308394 57854
rect 308630 57618 585342 57854
rect 585578 57618 585662 57854
rect 585898 57618 592650 57854
rect -8726 57586 592650 57618
rect -8726 54454 592650 54486
rect -8726 54218 -2934 54454
rect -2698 54218 -2614 54454
rect -2378 54218 293034 54454
rect 293270 54218 586302 54454
rect 586538 54218 586622 54454
rect 586858 54218 592650 54454
rect -8726 54134 592650 54218
rect -8726 53898 -2934 54134
rect -2698 53898 -2614 54134
rect -2378 53898 293034 54134
rect 293270 53898 586302 54134
rect 586538 53898 586622 54134
rect 586858 53898 592650 54134
rect -8726 53866 592650 53898
rect -8726 48174 592650 48206
rect -8726 47938 -1974 48174
rect -1738 47938 -1654 48174
rect -1418 47938 277674 48174
rect 277910 47938 308394 48174
rect 308630 47938 585342 48174
rect 585578 47938 585662 48174
rect 585898 47938 592650 48174
rect -8726 47854 592650 47938
rect -8726 47618 -1974 47854
rect -1738 47618 -1654 47854
rect -1418 47618 277674 47854
rect 277910 47618 308394 47854
rect 308630 47618 585342 47854
rect 585578 47618 585662 47854
rect 585898 47618 592650 47854
rect -8726 47586 592650 47618
rect -8726 44454 592650 44486
rect -8726 44218 -2934 44454
rect -2698 44218 -2614 44454
rect -2378 44218 293034 44454
rect 293270 44218 586302 44454
rect 586538 44218 586622 44454
rect 586858 44218 592650 44454
rect -8726 44134 592650 44218
rect -8726 43898 -2934 44134
rect -2698 43898 -2614 44134
rect -2378 43898 293034 44134
rect 293270 43898 586302 44134
rect 586538 43898 586622 44134
rect 586858 43898 592650 44134
rect -8726 43866 592650 43898
rect -8726 38174 592650 38206
rect -8726 37938 -1974 38174
rect -1738 37938 -1654 38174
rect -1418 37938 277674 38174
rect 277910 37938 308394 38174
rect 308630 37938 585342 38174
rect 585578 37938 585662 38174
rect 585898 37938 592650 38174
rect -8726 37854 592650 37938
rect -8726 37618 -1974 37854
rect -1738 37618 -1654 37854
rect -1418 37618 277674 37854
rect 277910 37618 308394 37854
rect 308630 37618 585342 37854
rect 585578 37618 585662 37854
rect 585898 37618 592650 37854
rect -8726 37586 592650 37618
rect -8726 34454 592650 34486
rect -8726 34218 -2934 34454
rect -2698 34218 -2614 34454
rect -2378 34218 293034 34454
rect 293270 34218 586302 34454
rect 586538 34218 586622 34454
rect 586858 34218 592650 34454
rect -8726 34134 592650 34218
rect -8726 33898 -2934 34134
rect -2698 33898 -2614 34134
rect -2378 33898 293034 34134
rect 293270 33898 586302 34134
rect 586538 33898 586622 34134
rect 586858 33898 592650 34134
rect -8726 33866 592650 33898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use tt_um_test  tt_top1.branch\[0\].col_um\[0\].um_bot_I.block_0_0.tt_um_I
timestamp 0
transform 1 0 9200 0 1 157216
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[0\].col_um\[0\].um_top_I.block_1_0.tt_um_I
timestamp 0
transform 1 0 9200 0 -1 212704
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[0\].col_um\[1\].um_bot_I.block_0_1.tt_um_I
timestamp 0
transform 1 0 43332 0 1 157216
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[0\].col_um\[1\].um_top_I.block_1_1.tt_um_I
timestamp 0
transform 1 0 43332 0 -1 212704
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[0\].col_um\[2\].um_bot_I.block_0_2.tt_um_I
timestamp 0
transform 1 0 77464 0 1 157216
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[0\].col_um\[2\].um_top_I.block_1_2.tt_um_I
timestamp 0
transform 1 0 77464 0 -1 212704
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[0\].col_um\[3\].um_bot_I.block_0_3.tt_um_I
timestamp 0
transform 1 0 111596 0 1 157216
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[0\].col_um\[3\].um_top_I.block_1_3.tt_um_I
timestamp 0
transform 1 0 111596 0 -1 212704
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[0\].col_um\[4\].um_bot_I.block_0_4.tt_um_I
timestamp 0
transform 1 0 145728 0 1 157216
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[0\].col_um\[4\].um_top_I.block_1_4.tt_um_I
timestamp 0
transform 1 0 145728 0 -1 212704
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[0\].col_um\[5\].um_bot_I.block_0_5.tt_um_I
timestamp 0
transform 1 0 179860 0 1 157216
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[0\].col_um\[5\].um_top_I.block_1_5.tt_um_I
timestamp 0
transform 1 0 179860 0 -1 212704
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[0\].col_um\[6\].um_bot_I.block_0_6.tt_um_I
timestamp 0
transform 1 0 213992 0 1 157216
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[0\].col_um\[6\].um_top_I.block_1_6.tt_um_I
timestamp 0
transform 1 0 213992 0 -1 212704
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[0\].col_um\[7\].um_bot_I.block_0_7.tt_um_I
timestamp 0
transform 1 0 248124 0 1 157216
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[0\].col_um\[7\].um_top_I.block_1_7.tt_um_I
timestamp 0
transform 1 0 248124 0 -1 212704
box 1066 1040 32632 21760
use tt_mux  tt_top1.branch\[0\].mux_I
timestamp 0
transform 1 0 9200 0 1 179520
box 750 0 272504 10880
use tt_um_test  tt_top1.branch\[1\].col_um\[0\].um_bot_I.block_0_16.tt_um_I
timestamp 0
transform -1 0 575000 0 1 157216
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[1\].col_um\[0\].um_top_I.block_1_16.tt_um_I
timestamp 0
transform -1 0 575000 0 -1 212704
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[1\].col_um\[1\].um_bot_I.block_0_17.tt_um_I
timestamp 0
transform -1 0 540868 0 1 157216
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[1\].col_um\[1\].um_top_I.block_1_17.tt_um_I
timestamp 0
transform -1 0 540868 0 -1 212704
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[1\].col_um\[2\].um_bot_I.block_0_18.tt_um_I
timestamp 0
transform -1 0 506736 0 1 157216
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[1\].col_um\[2\].um_top_I.block_1_18.tt_um_I
timestamp 0
transform -1 0 506736 0 -1 212704
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[1\].col_um\[3\].um_bot_I.block_0_19.tt_um_I
timestamp 0
transform -1 0 472604 0 1 157216
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[1\].col_um\[3\].um_top_I.block_1_19.tt_um_I
timestamp 0
transform -1 0 472604 0 -1 212704
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[1\].col_um\[4\].um_bot_I.block_0_20.tt_um_I
timestamp 0
transform -1 0 438472 0 1 157216
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[1\].col_um\[4\].um_top_I.block_1_20.tt_um_I
timestamp 0
transform -1 0 438472 0 -1 212704
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[1\].col_um\[5\].um_bot_I.block_0_21.tt_um_I
timestamp 0
transform -1 0 404340 0 1 157216
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[1\].col_um\[5\].um_top_I.block_1_21.tt_um_I
timestamp 0
transform -1 0 404340 0 -1 212704
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[1\].col_um\[6\].um_bot_I.block_0_22.tt_um_I
timestamp 0
transform -1 0 370208 0 1 157216
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[1\].col_um\[6\].um_top_I.block_1_22.tt_um_I
timestamp 0
transform -1 0 370208 0 -1 212704
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[1\].col_um\[7\].um_bot_I.block_0_23.tt_um_I
timestamp 0
transform -1 0 336076 0 1 157216
box 1066 1040 32632 21760
use tt_um_test  tt_top1.branch\[1\].col_um\[7\].um_top_I.block_1_23.tt_um_I
timestamp 0
transform -1 0 336076 0 -1 212704
box 1066 1040 32632 21760
use tt_mux  tt_top1.branch\[1\].mux_I
timestamp 0
transform -1 0 575000 0 1 179520
box 750 0 272504 10880
use tt_ctrl  tt_top1.ctrl_I
timestamp 0
transform 1 0 273424 0 1 21760
box 790 0 36010 44064
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 37586 592650 38206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 47586 592650 48206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 57586 592650 58206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 67586 592650 68206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 77586 592650 78206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 87586 592650 88206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 97586 592650 98206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 107586 592650 108206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 117586 592650 118206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 127586 592650 128206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 137586 592650 138206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 147586 592650 148206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 157586 592650 158206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 167586 592650 168206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 177586 592650 178206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 187586 592650 188206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 197586 592650 198206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 207586 592650 208206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 217586 592650 218206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 227586 592650 228206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 237586 592650 238206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 247586 592650 248206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 257586 592650 258206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 267586 592650 268206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 277586 592650 278206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 287586 592650 288206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 297586 592650 298206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 307586 592650 308206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 317586 592650 318206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 327586 592650 328206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 337586 592650 338206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 347586 592650 348206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 357586 592650 358206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 367586 592650 368206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 377586 592650 378206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 387586 592650 388206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 397586 592650 398206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 407586 592650 408206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 417586 592650 418206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 427586 592650 428206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 437586 592650 438206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 447586 592650 448206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 457586 592650 458206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 467586 592650 468206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 477586 592650 478206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 487586 592650 488206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 497586 592650 498206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 507586 592650 508206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 517586 592650 518206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 527586 592650 528206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 537586 592650 538206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 547586 592650 548206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 557586 592650 558206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 567586 592650 568206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 577586 592650 578206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 587586 592650 588206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 597586 592650 598206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 607586 592650 608206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 617586 592650 618206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 627586 592650 628206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 637586 592650 638206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 647586 592650 648206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 657586 592650 658206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 667586 592650 668206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 677586 592650 678206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 687586 592650 688206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 697586 592650 698206 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 33866 592650 34486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43866 592650 44486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 53866 592650 54486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 63866 592650 64486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 73866 592650 74486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 93866 592650 94486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 103866 592650 104486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 113866 592650 114486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 123866 592650 124486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 133866 592650 134486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 143866 592650 144486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 153866 592650 154486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 163866 592650 164486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 183866 592650 184486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 193866 592650 194486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 203866 592650 204486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 213866 592650 214486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223866 592650 224486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 233866 592650 234486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 243866 592650 244486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 253866 592650 254486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 273866 592650 274486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 283866 592650 284486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 293866 592650 294486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 303866 592650 304486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 313866 592650 314486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 323866 592650 324486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 333866 592650 334486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 343866 592650 344486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 363866 592650 364486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 373866 592650 374486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 383866 592650 384486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 393866 592650 394486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403866 592650 404486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 413866 592650 414486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 423866 592650 424486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 433866 592650 434486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 453866 592650 454486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 463866 592650 464486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 473866 592650 474486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 483866 592650 484486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 493866 592650 494486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 503866 592650 504486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 513866 592650 514486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 523866 592650 524486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 543866 592650 544486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 553866 592650 554486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 563866 592650 564486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 573866 592650 574486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583866 592650 584486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 593866 592650 594486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 603866 592650 604486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 613866 592650 614486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 633866 592650 634486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 643866 592650 644486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 653866 592650 654486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 663866 592650 664486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 673866 592650 674486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 683866 592650 684486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 693866 592650 694486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
