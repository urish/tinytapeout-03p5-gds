VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_as1802
  CLASS BLOCK ;
  FOREIGN tt_um_as1802 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1362.520 BY 220.320 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 215.750 158.850 220.320 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 162.230 219.320 162.530 220.320 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 216.740 155.170 220.320 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 218.780 151.490 220.320 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 215.380 147.810 220.320 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 214.020 144.130 220.320 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 216.740 140.450 220.320 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 217.420 136.770 220.320 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 218.780 133.090 220.320 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 215.380 129.410 220.320 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 219.320 125.730 220.320 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 217.420 122.050 220.320 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 218.780 118.370 220.320 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 217.420 114.690 220.320 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 214.020 111.010 220.320 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 218.780 107.330 220.320 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 215.380 103.650 220.320 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 216.740 99.970 220.320 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 216.740 96.290 220.320 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 218.780 33.730 220.320 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 218.780 30.050 220.320 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 214.700 26.370 220.320 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 218.780 22.690 220.320 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 219.150 19.010 220.320 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 218.780 15.330 220.320 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 218.780 11.650 220.320 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 218.780 7.970 220.320 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 218.780 63.170 220.320 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 218.780 59.490 220.320 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 193.620 55.810 220.320 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 218.780 52.130 220.320 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 193.620 48.450 220.320 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 218.780 44.770 220.320 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 218.780 41.090 220.320 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 218.780 37.410 220.320 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 218.780 92.610 220.320 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 218.780 88.930 220.320 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 218.780 85.250 220.320 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 211.980 81.570 220.320 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 218.780 77.890 220.320 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 214.700 74.210 220.320 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 218.780 70.530 220.320 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 218.780 66.850 220.320 ;
    END
  END uo_out[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 5.200 22.640 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 5.200 176.240 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 5.200 329.840 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 5.200 483.440 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 5.200 637.040 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 5.200 790.640 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 5.200 944.240 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 5.200 1097.840 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 5.200 1251.440 215.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 5.200 99.440 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 5.200 253.040 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 5.200 406.640 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 5.200 560.240 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 5.200 713.840 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 5.200 867.440 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 5.200 1021.040 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 5.200 1174.640 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 5.200 1328.240 215.120 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 213.465 1357.190 215.070 ;
        RECT 5.330 208.025 1357.190 210.855 ;
        RECT 5.330 202.585 1357.190 205.415 ;
        RECT 5.330 197.145 1357.190 199.975 ;
        RECT 5.330 191.705 1357.190 194.535 ;
        RECT 5.330 186.265 1357.190 189.095 ;
        RECT 5.330 180.825 1357.190 183.655 ;
        RECT 5.330 175.385 1357.190 178.215 ;
        RECT 5.330 169.945 1357.190 172.775 ;
        RECT 5.330 164.505 1357.190 167.335 ;
        RECT 5.330 159.065 1357.190 161.895 ;
        RECT 5.330 153.625 1357.190 156.455 ;
        RECT 5.330 148.185 1357.190 151.015 ;
        RECT 5.330 142.745 1357.190 145.575 ;
        RECT 5.330 137.305 1357.190 140.135 ;
        RECT 5.330 131.865 1357.190 134.695 ;
        RECT 5.330 126.425 1357.190 129.255 ;
        RECT 5.330 120.985 1357.190 123.815 ;
        RECT 5.330 115.545 1357.190 118.375 ;
        RECT 5.330 110.105 1357.190 112.935 ;
        RECT 5.330 104.665 1357.190 107.495 ;
        RECT 5.330 99.225 1357.190 102.055 ;
        RECT 5.330 93.785 1357.190 96.615 ;
        RECT 5.330 88.345 1357.190 91.175 ;
        RECT 5.330 82.905 1357.190 85.735 ;
        RECT 5.330 77.465 1357.190 80.295 ;
        RECT 5.330 72.025 1357.190 74.855 ;
        RECT 5.330 66.585 1357.190 69.415 ;
        RECT 5.330 61.145 1357.190 63.975 ;
        RECT 5.330 55.705 1357.190 58.535 ;
        RECT 5.330 50.265 1357.190 53.095 ;
        RECT 5.330 44.825 1357.190 47.655 ;
        RECT 5.330 39.385 1357.190 42.215 ;
        RECT 5.330 33.945 1357.190 36.775 ;
        RECT 5.330 28.505 1357.190 31.335 ;
        RECT 5.330 23.065 1357.190 25.895 ;
        RECT 5.330 17.625 1357.190 20.455 ;
        RECT 5.330 12.185 1357.190 15.015 ;
        RECT 5.330 6.745 1357.190 9.575 ;
      LAYER li1 ;
        RECT 5.520 5.355 1357.000 214.965 ;
      LAYER met1 ;
        RECT 5.520 0.720 1357.000 220.280 ;
      LAYER met2 ;
        RECT 10.670 0.155 1353.680 220.310 ;
      LAYER met3 ;
        RECT 7.630 0.175 1349.575 219.465 ;
      LAYER met4 ;
        RECT 8.370 218.380 10.950 219.465 ;
        RECT 12.050 218.380 14.630 219.465 ;
        RECT 15.730 218.750 18.310 219.465 ;
        RECT 19.410 218.750 21.990 219.465 ;
        RECT 15.730 218.380 21.990 218.750 ;
        RECT 23.090 218.380 25.670 219.465 ;
        RECT 7.655 215.520 25.670 218.380 ;
        RECT 7.655 4.800 20.640 215.520 ;
        RECT 23.040 214.300 25.670 215.520 ;
        RECT 26.770 218.380 29.350 219.465 ;
        RECT 30.450 218.380 33.030 219.465 ;
        RECT 34.130 218.380 36.710 219.465 ;
        RECT 37.810 218.380 40.390 219.465 ;
        RECT 41.490 218.380 44.070 219.465 ;
        RECT 45.170 218.380 47.750 219.465 ;
        RECT 26.770 214.300 47.750 218.380 ;
        RECT 23.040 193.220 47.750 214.300 ;
        RECT 48.850 218.380 51.430 219.465 ;
        RECT 52.530 218.380 55.110 219.465 ;
        RECT 48.850 193.220 55.110 218.380 ;
        RECT 56.210 218.380 58.790 219.465 ;
        RECT 59.890 218.380 62.470 219.465 ;
        RECT 63.570 218.380 66.150 219.465 ;
        RECT 67.250 218.380 69.830 219.465 ;
        RECT 70.930 218.380 73.510 219.465 ;
        RECT 56.210 214.300 73.510 218.380 ;
        RECT 74.610 218.380 77.190 219.465 ;
        RECT 78.290 218.380 80.870 219.465 ;
        RECT 74.610 214.300 80.870 218.380 ;
        RECT 56.210 211.580 80.870 214.300 ;
        RECT 81.970 218.380 84.550 219.465 ;
        RECT 85.650 218.380 88.230 219.465 ;
        RECT 89.330 218.380 91.910 219.465 ;
        RECT 93.010 218.380 95.590 219.465 ;
        RECT 81.970 216.340 95.590 218.380 ;
        RECT 96.690 216.340 99.270 219.465 ;
        RECT 100.370 216.340 102.950 219.465 ;
        RECT 81.970 215.520 102.950 216.340 ;
        RECT 81.970 211.580 97.440 215.520 ;
        RECT 56.210 193.220 97.440 211.580 ;
        RECT 23.040 4.800 97.440 193.220 ;
        RECT 99.840 214.980 102.950 215.520 ;
        RECT 104.050 218.380 106.630 219.465 ;
        RECT 107.730 218.380 110.310 219.465 ;
        RECT 104.050 214.980 110.310 218.380 ;
        RECT 99.840 213.620 110.310 214.980 ;
        RECT 111.410 217.020 113.990 219.465 ;
        RECT 115.090 218.380 117.670 219.465 ;
        RECT 118.770 218.380 121.350 219.465 ;
        RECT 115.090 217.020 121.350 218.380 ;
        RECT 122.450 218.920 125.030 219.465 ;
        RECT 126.130 218.920 128.710 219.465 ;
        RECT 122.450 217.020 128.710 218.920 ;
        RECT 111.410 214.980 128.710 217.020 ;
        RECT 129.810 218.380 132.390 219.465 ;
        RECT 133.490 218.380 136.070 219.465 ;
        RECT 129.810 217.020 136.070 218.380 ;
        RECT 137.170 217.020 139.750 219.465 ;
        RECT 129.810 216.340 139.750 217.020 ;
        RECT 140.850 216.340 143.430 219.465 ;
        RECT 129.810 214.980 143.430 216.340 ;
        RECT 111.410 213.620 143.430 214.980 ;
        RECT 144.530 214.980 147.110 219.465 ;
        RECT 148.210 218.380 150.790 219.465 ;
        RECT 151.890 218.380 154.470 219.465 ;
        RECT 148.210 216.340 154.470 218.380 ;
        RECT 155.570 216.340 158.150 219.465 ;
        RECT 148.210 215.350 158.150 216.340 ;
        RECT 159.250 218.920 161.830 219.465 ;
        RECT 162.930 218.920 1170.865 219.465 ;
        RECT 159.250 215.520 1170.865 218.920 ;
        RECT 159.250 215.350 174.240 215.520 ;
        RECT 148.210 214.980 174.240 215.350 ;
        RECT 144.530 213.620 174.240 214.980 ;
        RECT 99.840 4.800 174.240 213.620 ;
        RECT 176.640 4.800 251.040 215.520 ;
        RECT 253.440 4.800 327.840 215.520 ;
        RECT 330.240 4.800 404.640 215.520 ;
        RECT 407.040 4.800 481.440 215.520 ;
        RECT 483.840 4.800 558.240 215.520 ;
        RECT 560.640 4.800 635.040 215.520 ;
        RECT 637.440 4.800 711.840 215.520 ;
        RECT 714.240 4.800 788.640 215.520 ;
        RECT 791.040 4.800 865.440 215.520 ;
        RECT 867.840 4.800 942.240 215.520 ;
        RECT 944.640 4.800 1019.040 215.520 ;
        RECT 1021.440 4.800 1095.840 215.520 ;
        RECT 1098.240 4.800 1170.865 215.520 ;
        RECT 7.655 0.175 1170.865 4.800 ;
  END
END tt_um_as1802
END LIBRARY

