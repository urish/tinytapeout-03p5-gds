* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for tt_um_TrainLED2_top abstract view
.subckt tt_um_TrainLED2_top clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4]
+ ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5]
+ uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5]
+ uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5]
+ uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5]
+ uo_out[6] uo_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tt_um_as1802 abstract view
.subckt tt_um_as1802 clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5]
+ ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6]
+ uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6]
+ uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6]
+ uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6]
+ uo_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tt_um_test abstract view
.subckt tt_um_test clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5]
+ ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6]
+ uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6]
+ uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6]
+ uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6]
+ uo_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tt_mux abstract view
.subckt tt_mux addr[0] addr[1] addr[2] addr[3] addr[4] k_one k_zero spine_iw[0] spine_iw[10]
+ spine_iw[11] spine_iw[12] spine_iw[13] spine_iw[14] spine_iw[15] spine_iw[16] spine_iw[17]
+ spine_iw[18] spine_iw[19] spine_iw[1] spine_iw[20] spine_iw[21] spine_iw[22] spine_iw[23]
+ spine_iw[24] spine_iw[25] spine_iw[26] spine_iw[27] spine_iw[28] spine_iw[29] spine_iw[2]
+ spine_iw[30] spine_iw[3] spine_iw[4] spine_iw[5] spine_iw[6] spine_iw[7] spine_iw[8]
+ spine_iw[9] spine_ow[0] spine_ow[10] spine_ow[11] spine_ow[12] spine_ow[13] spine_ow[14]
+ spine_ow[15] spine_ow[16] spine_ow[17] spine_ow[18] spine_ow[19] spine_ow[1] spine_ow[20]
+ spine_ow[21] spine_ow[22] spine_ow[23] spine_ow[24] spine_ow[25] spine_ow[2] spine_ow[3]
+ spine_ow[4] spine_ow[5] spine_ow[6] spine_ow[7] spine_ow[8] spine_ow[9] um_ena[0]
+ um_ena[10] um_ena[11] um_ena[12] um_ena[13] um_ena[14] um_ena[15] um_ena[1] um_ena[2]
+ um_ena[3] um_ena[4] um_ena[5] um_ena[6] um_ena[7] um_ena[8] um_ena[9] um_iw[0] um_iw[100]
+ um_iw[101] um_iw[102] um_iw[103] um_iw[104] um_iw[105] um_iw[106] um_iw[107] um_iw[108]
+ um_iw[109] um_iw[10] um_iw[110] um_iw[111] um_iw[112] um_iw[113] um_iw[114] um_iw[115]
+ um_iw[116] um_iw[117] um_iw[118] um_iw[119] um_iw[11] um_iw[120] um_iw[121] um_iw[122]
+ um_iw[123] um_iw[124] um_iw[125] um_iw[126] um_iw[127] um_iw[128] um_iw[129] um_iw[12]
+ um_iw[130] um_iw[131] um_iw[132] um_iw[133] um_iw[134] um_iw[135] um_iw[136] um_iw[137]
+ um_iw[138] um_iw[139] um_iw[13] um_iw[140] um_iw[141] um_iw[142] um_iw[143] um_iw[144]
+ um_iw[145] um_iw[146] um_iw[147] um_iw[148] um_iw[149] um_iw[14] um_iw[150] um_iw[151]
+ um_iw[152] um_iw[153] um_iw[154] um_iw[155] um_iw[156] um_iw[157] um_iw[158] um_iw[159]
+ um_iw[15] um_iw[160] um_iw[161] um_iw[162] um_iw[163] um_iw[164] um_iw[165] um_iw[166]
+ um_iw[167] um_iw[168] um_iw[169] um_iw[16] um_iw[170] um_iw[171] um_iw[172] um_iw[173]
+ um_iw[174] um_iw[175] um_iw[176] um_iw[177] um_iw[178] um_iw[179] um_iw[17] um_iw[180]
+ um_iw[181] um_iw[182] um_iw[183] um_iw[184] um_iw[185] um_iw[186] um_iw[187] um_iw[188]
+ um_iw[189] um_iw[18] um_iw[190] um_iw[191] um_iw[192] um_iw[193] um_iw[194] um_iw[195]
+ um_iw[196] um_iw[197] um_iw[198] um_iw[199] um_iw[19] um_iw[1] um_iw[200] um_iw[201]
+ um_iw[202] um_iw[203] um_iw[204] um_iw[205] um_iw[206] um_iw[207] um_iw[208] um_iw[209]
+ um_iw[20] um_iw[210] um_iw[211] um_iw[212] um_iw[213] um_iw[214] um_iw[215] um_iw[216]
+ um_iw[217] um_iw[218] um_iw[219] um_iw[21] um_iw[220] um_iw[221] um_iw[222] um_iw[223]
+ um_iw[224] um_iw[225] um_iw[226] um_iw[227] um_iw[228] um_iw[229] um_iw[22] um_iw[230]
+ um_iw[231] um_iw[232] um_iw[233] um_iw[234] um_iw[235] um_iw[236] um_iw[237] um_iw[238]
+ um_iw[239] um_iw[23] um_iw[240] um_iw[241] um_iw[242] um_iw[243] um_iw[244] um_iw[245]
+ um_iw[246] um_iw[247] um_iw[248] um_iw[249] um_iw[24] um_iw[250] um_iw[251] um_iw[252]
+ um_iw[253] um_iw[254] um_iw[255] um_iw[256] um_iw[257] um_iw[258] um_iw[259] um_iw[25]
+ um_iw[260] um_iw[261] um_iw[262] um_iw[263] um_iw[264] um_iw[265] um_iw[266] um_iw[267]
+ um_iw[268] um_iw[269] um_iw[26] um_iw[270] um_iw[271] um_iw[272] um_iw[273] um_iw[274]
+ um_iw[275] um_iw[276] um_iw[277] um_iw[278] um_iw[279] um_iw[27] um_iw[280] um_iw[281]
+ um_iw[282] um_iw[283] um_iw[284] um_iw[285] um_iw[286] um_iw[287] um_iw[28] um_iw[29]
+ um_iw[2] um_iw[30] um_iw[31] um_iw[32] um_iw[33] um_iw[34] um_iw[35] um_iw[36] um_iw[37]
+ um_iw[38] um_iw[39] um_iw[3] um_iw[40] um_iw[41] um_iw[42] um_iw[43] um_iw[44] um_iw[45]
+ um_iw[46] um_iw[47] um_iw[48] um_iw[49] um_iw[4] um_iw[50] um_iw[51] um_iw[52] um_iw[53]
+ um_iw[54] um_iw[55] um_iw[56] um_iw[57] um_iw[58] um_iw[59] um_iw[5] um_iw[60] um_iw[61]
+ um_iw[62] um_iw[63] um_iw[64] um_iw[65] um_iw[66] um_iw[67] um_iw[68] um_iw[69]
+ um_iw[6] um_iw[70] um_iw[71] um_iw[72] um_iw[73] um_iw[74] um_iw[75] um_iw[76] um_iw[77]
+ um_iw[78] um_iw[79] um_iw[7] um_iw[80] um_iw[81] um_iw[82] um_iw[83] um_iw[84] um_iw[85]
+ um_iw[86] um_iw[87] um_iw[88] um_iw[89] um_iw[8] um_iw[90] um_iw[91] um_iw[92] um_iw[93]
+ um_iw[94] um_iw[95] um_iw[96] um_iw[97] um_iw[98] um_iw[99] um_iw[9] um_k_zero[0]
+ um_k_zero[10] um_k_zero[11] um_k_zero[12] um_k_zero[13] um_k_zero[14] um_k_zero[15]
+ um_k_zero[1] um_k_zero[2] um_k_zero[3] um_k_zero[4] um_k_zero[5] um_k_zero[6] um_k_zero[7]
+ um_k_zero[8] um_k_zero[9] um_ow[0] um_ow[100] um_ow[101] um_ow[102] um_ow[103] um_ow[104]
+ um_ow[105] um_ow[106] um_ow[107] um_ow[108] um_ow[109] um_ow[10] um_ow[110] um_ow[111]
+ um_ow[112] um_ow[113] um_ow[114] um_ow[115] um_ow[116] um_ow[117] um_ow[118] um_ow[119]
+ um_ow[11] um_ow[120] um_ow[121] um_ow[122] um_ow[123] um_ow[124] um_ow[125] um_ow[126]
+ um_ow[127] um_ow[128] um_ow[129] um_ow[12] um_ow[130] um_ow[131] um_ow[132] um_ow[133]
+ um_ow[134] um_ow[135] um_ow[136] um_ow[137] um_ow[138] um_ow[139] um_ow[13] um_ow[140]
+ um_ow[141] um_ow[142] um_ow[143] um_ow[144] um_ow[145] um_ow[146] um_ow[147] um_ow[148]
+ um_ow[149] um_ow[14] um_ow[150] um_ow[151] um_ow[152] um_ow[153] um_ow[154] um_ow[155]
+ um_ow[156] um_ow[157] um_ow[158] um_ow[159] um_ow[15] um_ow[160] um_ow[161] um_ow[162]
+ um_ow[163] um_ow[164] um_ow[165] um_ow[166] um_ow[167] um_ow[168] um_ow[169] um_ow[16]
+ um_ow[170] um_ow[171] um_ow[172] um_ow[173] um_ow[174] um_ow[175] um_ow[176] um_ow[177]
+ um_ow[178] um_ow[179] um_ow[17] um_ow[180] um_ow[181] um_ow[182] um_ow[183] um_ow[184]
+ um_ow[185] um_ow[186] um_ow[187] um_ow[188] um_ow[189] um_ow[18] um_ow[190] um_ow[191]
+ um_ow[192] um_ow[193] um_ow[194] um_ow[195] um_ow[196] um_ow[197] um_ow[198] um_ow[199]
+ um_ow[19] um_ow[1] um_ow[200] um_ow[201] um_ow[202] um_ow[203] um_ow[204] um_ow[205]
+ um_ow[206] um_ow[207] um_ow[208] um_ow[209] um_ow[20] um_ow[210] um_ow[211] um_ow[212]
+ um_ow[213] um_ow[214] um_ow[215] um_ow[216] um_ow[217] um_ow[218] um_ow[219] um_ow[21]
+ um_ow[220] um_ow[221] um_ow[222] um_ow[223] um_ow[224] um_ow[225] um_ow[226] um_ow[227]
+ um_ow[228] um_ow[229] um_ow[22] um_ow[230] um_ow[231] um_ow[232] um_ow[233] um_ow[234]
+ um_ow[235] um_ow[236] um_ow[237] um_ow[238] um_ow[239] um_ow[23] um_ow[240] um_ow[241]
+ um_ow[242] um_ow[243] um_ow[244] um_ow[245] um_ow[246] um_ow[247] um_ow[248] um_ow[249]
+ um_ow[24] um_ow[250] um_ow[251] um_ow[252] um_ow[253] um_ow[254] um_ow[255] um_ow[256]
+ um_ow[257] um_ow[258] um_ow[259] um_ow[25] um_ow[260] um_ow[261] um_ow[262] um_ow[263]
+ um_ow[264] um_ow[265] um_ow[266] um_ow[267] um_ow[268] um_ow[269] um_ow[26] um_ow[270]
+ um_ow[271] um_ow[272] um_ow[273] um_ow[274] um_ow[275] um_ow[276] um_ow[277] um_ow[278]
+ um_ow[279] um_ow[27] um_ow[280] um_ow[281] um_ow[282] um_ow[283] um_ow[284] um_ow[285]
+ um_ow[286] um_ow[287] um_ow[288] um_ow[289] um_ow[28] um_ow[290] um_ow[291] um_ow[292]
+ um_ow[293] um_ow[294] um_ow[295] um_ow[296] um_ow[297] um_ow[298] um_ow[299] um_ow[29]
+ um_ow[2] um_ow[300] um_ow[301] um_ow[302] um_ow[303] um_ow[304] um_ow[305] um_ow[306]
+ um_ow[307] um_ow[308] um_ow[309] um_ow[30] um_ow[310] um_ow[311] um_ow[312] um_ow[313]
+ um_ow[314] um_ow[315] um_ow[316] um_ow[317] um_ow[318] um_ow[319] um_ow[31] um_ow[320]
+ um_ow[321] um_ow[322] um_ow[323] um_ow[324] um_ow[325] um_ow[326] um_ow[327] um_ow[328]
+ um_ow[329] um_ow[32] um_ow[330] um_ow[331] um_ow[332] um_ow[333] um_ow[334] um_ow[335]
+ um_ow[336] um_ow[337] um_ow[338] um_ow[339] um_ow[33] um_ow[340] um_ow[341] um_ow[342]
+ um_ow[343] um_ow[344] um_ow[345] um_ow[346] um_ow[347] um_ow[348] um_ow[349] um_ow[34]
+ um_ow[350] um_ow[351] um_ow[352] um_ow[353] um_ow[354] um_ow[355] um_ow[356] um_ow[357]
+ um_ow[358] um_ow[359] um_ow[35] um_ow[360] um_ow[361] um_ow[362] um_ow[363] um_ow[364]
+ um_ow[365] um_ow[366] um_ow[367] um_ow[368] um_ow[369] um_ow[36] um_ow[370] um_ow[371]
+ um_ow[372] um_ow[373] um_ow[374] um_ow[375] um_ow[376] um_ow[377] um_ow[378] um_ow[379]
+ um_ow[37] um_ow[380] um_ow[381] um_ow[382] um_ow[383] um_ow[38] um_ow[39] um_ow[3]
+ um_ow[40] um_ow[41] um_ow[42] um_ow[43] um_ow[44] um_ow[45] um_ow[46] um_ow[47]
+ um_ow[48] um_ow[49] um_ow[4] um_ow[50] um_ow[51] um_ow[52] um_ow[53] um_ow[54] um_ow[55]
+ um_ow[56] um_ow[57] um_ow[58] um_ow[59] um_ow[5] um_ow[60] um_ow[61] um_ow[62] um_ow[63]
+ um_ow[64] um_ow[65] um_ow[66] um_ow[67] um_ow[68] um_ow[69] um_ow[6] um_ow[70] um_ow[71]
+ um_ow[72] um_ow[73] um_ow[74] um_ow[75] um_ow[76] um_ow[77] um_ow[78] um_ow[79]
+ um_ow[7] um_ow[80] um_ow[81] um_ow[82] um_ow[83] um_ow[84] um_ow[85] um_ow[86] um_ow[87]
+ um_ow[88] um_ow[89] um_ow[8] um_ow[90] um_ow[91] um_ow[92] um_ow[93] um_ow[94] um_ow[95]
+ um_ow[96] um_ow[97] um_ow[98] um_ow[99] um_ow[9] vccd1 vssd1
.ends

* Black-box entry subcircuit for tt_ctrl abstract view
.subckt tt_ctrl ctrl_ena ctrl_sel_inc ctrl_sel_rst_n k_one k_zero pad_ui_in[0] pad_ui_in[1]
+ pad_ui_in[2] pad_ui_in[3] pad_ui_in[4] pad_ui_in[5] pad_ui_in[6] pad_ui_in[7] pad_ui_in[8]
+ pad_ui_in[9] pad_uio_in[0] pad_uio_in[1] pad_uio_in[2] pad_uio_in[3] pad_uio_in[4]
+ pad_uio_in[5] pad_uio_in[6] pad_uio_in[7] pad_uio_oe_n[0] pad_uio_oe_n[1] pad_uio_oe_n[2]
+ pad_uio_oe_n[3] pad_uio_oe_n[4] pad_uio_oe_n[5] pad_uio_oe_n[6] pad_uio_oe_n[7]
+ pad_uio_out[0] pad_uio_out[1] pad_uio_out[2] pad_uio_out[3] pad_uio_out[4] pad_uio_out[5]
+ pad_uio_out[6] pad_uio_out[7] pad_uo_out[0] pad_uo_out[1] pad_uo_out[2] pad_uo_out[3]
+ pad_uo_out[4] pad_uo_out[5] pad_uo_out[6] pad_uo_out[7] spine_iw[0] spine_iw[10]
+ spine_iw[11] spine_iw[12] spine_iw[13] spine_iw[14] spine_iw[15] spine_iw[16] spine_iw[17]
+ spine_iw[18] spine_iw[19] spine_iw[1] spine_iw[20] spine_iw[21] spine_iw[22] spine_iw[23]
+ spine_iw[24] spine_iw[25] spine_iw[26] spine_iw[27] spine_iw[28] spine_iw[29] spine_iw[2]
+ spine_iw[30] spine_iw[3] spine_iw[4] spine_iw[5] spine_iw[6] spine_iw[7] spine_iw[8]
+ spine_iw[9] spine_ow[0] spine_ow[10] spine_ow[11] spine_ow[12] spine_ow[13] spine_ow[14]
+ spine_ow[15] spine_ow[16] spine_ow[17] spine_ow[18] spine_ow[19] spine_ow[1] spine_ow[20]
+ spine_ow[21] spine_ow[22] spine_ow[23] spine_ow[24] spine_ow[25] spine_ow[2] spine_ow[3]
+ spine_ow[4] spine_ow[5] spine_ow[6] spine_ow[7] spine_ow[8] spine_ow[9] vccd1 vssd1
.ends

* Black-box entry subcircuit for tt_um_moyes0_top_module abstract view
.subckt tt_um_moyes0_top_module clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tt_um_urish_dffram abstract view
.subckt tt_um_urish_dffram clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4]
+ ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5]
+ uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5]
+ uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5]
+ uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5]
+ uo_out[6] uo_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tt_um_cam abstract view
.subckt tt_um_cam clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5]
+ ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6]
+ uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6]
+ uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6]
+ uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6]
+ uo_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tt_um_MichaelBell_hovalaag abstract view
.subckt tt_um_MichaelBell_hovalaag clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tt_um_urish_simon abstract view
.subckt tt_um_urish_simon clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4]
+ ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5]
+ uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5]
+ uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5]
+ uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5]
+ uo_out[6] uo_out[7] vccd1 vssd1
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[30] io_oeb[31] io_out[16] io_out[17] io_out[18] io_out[19] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[30] io_out[31] io_out[4] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
Xtt_top1.branch\[1\].col_um\[0\].um_bot_I.block_0_16.tt_um_I tt_top1.branch\[1\].mux_I/um_iw[0]
+ tt_top1.branch\[1\].mux_I/um_ena[0] tt_top1.branch\[1\].mux_I/um_iw[1] tt_top1.branch\[1\].mux_I/um_iw[2]
+ tt_top1.branch\[1\].mux_I/um_iw[3] tt_top1.branch\[1\].mux_I/um_iw[4] tt_top1.branch\[1\].mux_I/um_iw[5]
+ tt_top1.branch\[1\].mux_I/um_iw[6] tt_top1.branch\[1\].mux_I/um_iw[7] tt_top1.branch\[1\].mux_I/um_iw[8]
+ tt_top1.branch\[1\].mux_I/um_iw[9] tt_top1.branch\[1\].mux_I/um_iw[10] tt_top1.branch\[1\].mux_I/um_iw[11]
+ tt_top1.branch\[1\].mux_I/um_iw[12] tt_top1.branch\[1\].mux_I/um_iw[13] tt_top1.branch\[1\].mux_I/um_iw[14]
+ tt_top1.branch\[1\].mux_I/um_iw[15] tt_top1.branch\[1\].mux_I/um_iw[16] tt_top1.branch\[1\].mux_I/um_iw[17]
+ tt_top1.branch\[1\].mux_I/um_ow[16] tt_top1.branch\[1\].mux_I/um_ow[17] tt_top1.branch\[1\].mux_I/um_ow[18]
+ tt_top1.branch\[1\].mux_I/um_ow[19] tt_top1.branch\[1\].mux_I/um_ow[20] tt_top1.branch\[1\].mux_I/um_ow[21]
+ tt_top1.branch\[1\].mux_I/um_ow[22] tt_top1.branch\[1\].mux_I/um_ow[23] tt_top1.branch\[1\].mux_I/um_ow[8]
+ tt_top1.branch\[1\].mux_I/um_ow[9] tt_top1.branch\[1\].mux_I/um_ow[10] tt_top1.branch\[1\].mux_I/um_ow[11]
+ tt_top1.branch\[1\].mux_I/um_ow[12] tt_top1.branch\[1\].mux_I/um_ow[13] tt_top1.branch\[1\].mux_I/um_ow[14]
+ tt_top1.branch\[1\].mux_I/um_ow[15] tt_top1.branch\[1\].mux_I/um_ow[0] tt_top1.branch\[1\].mux_I/um_ow[1]
+ tt_top1.branch\[1\].mux_I/um_ow[2] tt_top1.branch\[1\].mux_I/um_ow[3] tt_top1.branch\[1\].mux_I/um_ow[4]
+ tt_top1.branch\[1\].mux_I/um_ow[5] tt_top1.branch\[1\].mux_I/um_ow[6] tt_top1.branch\[1\].mux_I/um_ow[7]
+ vccd1 vssd1 tt_um_TrainLED2_top
Xtt_top1.branch\[0\].col_um\[0\].um_bot_I.block_0_0.tt_um_I tt_top1.branch\[0\].mux_I/um_iw[0]
+ tt_top1.branch\[0\].mux_I/um_ena[0] tt_top1.branch\[0\].mux_I/um_iw[1] tt_top1.branch\[0\].mux_I/um_iw[2]
+ tt_top1.branch\[0\].mux_I/um_iw[3] tt_top1.branch\[0\].mux_I/um_iw[4] tt_top1.branch\[0\].mux_I/um_iw[5]
+ tt_top1.branch\[0\].mux_I/um_iw[6] tt_top1.branch\[0\].mux_I/um_iw[7] tt_top1.branch\[0\].mux_I/um_iw[8]
+ tt_top1.branch\[0\].mux_I/um_iw[9] tt_top1.branch\[0\].mux_I/um_iw[10] tt_top1.branch\[0\].mux_I/um_iw[11]
+ tt_top1.branch\[0\].mux_I/um_iw[12] tt_top1.branch\[0\].mux_I/um_iw[13] tt_top1.branch\[0\].mux_I/um_iw[14]
+ tt_top1.branch\[0\].mux_I/um_iw[15] tt_top1.branch\[0\].mux_I/um_iw[16] tt_top1.branch\[0\].mux_I/um_iw[17]
+ tt_top1.branch\[0\].mux_I/um_ow[16] tt_top1.branch\[0\].mux_I/um_ow[17] tt_top1.branch\[0\].mux_I/um_ow[18]
+ tt_top1.branch\[0\].mux_I/um_ow[19] tt_top1.branch\[0\].mux_I/um_ow[20] tt_top1.branch\[0\].mux_I/um_ow[21]
+ tt_top1.branch\[0\].mux_I/um_ow[22] tt_top1.branch\[0\].mux_I/um_ow[23] tt_top1.branch\[0\].mux_I/um_ow[8]
+ tt_top1.branch\[0\].mux_I/um_ow[9] tt_top1.branch\[0\].mux_I/um_ow[10] tt_top1.branch\[0\].mux_I/um_ow[11]
+ tt_top1.branch\[0\].mux_I/um_ow[12] tt_top1.branch\[0\].mux_I/um_ow[13] tt_top1.branch\[0\].mux_I/um_ow[14]
+ tt_top1.branch\[0\].mux_I/um_ow[15] tt_top1.branch\[0\].mux_I/um_ow[0] tt_top1.branch\[0\].mux_I/um_ow[1]
+ tt_top1.branch\[0\].mux_I/um_ow[2] tt_top1.branch\[0\].mux_I/um_ow[3] tt_top1.branch\[0\].mux_I/um_ow[4]
+ tt_top1.branch\[0\].mux_I/um_ow[5] tt_top1.branch\[0\].mux_I/um_ow[6] tt_top1.branch\[0\].mux_I/um_ow[7]
+ vccd1 vssd1 tt_um_as1802
Xtt_top1.branch\[1\].col_um\[7\].um_top_I.block_1_23.tt_um_I tt_top1.branch\[1\].mux_I/um_iw[270]
+ tt_top1.branch\[1\].mux_I/um_ena[15] tt_top1.branch\[1\].mux_I/um_iw[271] tt_top1.branch\[1\].mux_I/um_iw[272]
+ tt_top1.branch\[1\].mux_I/um_iw[273] tt_top1.branch\[1\].mux_I/um_iw[274] tt_top1.branch\[1\].mux_I/um_iw[275]
+ tt_top1.branch\[1\].mux_I/um_iw[276] tt_top1.branch\[1\].mux_I/um_iw[277] tt_top1.branch\[1\].mux_I/um_iw[278]
+ tt_top1.branch\[1\].mux_I/um_iw[279] tt_top1.branch\[1\].mux_I/um_iw[280] tt_top1.branch\[1\].mux_I/um_iw[281]
+ tt_top1.branch\[1\].mux_I/um_iw[282] tt_top1.branch\[1\].mux_I/um_iw[283] tt_top1.branch\[1\].mux_I/um_iw[284]
+ tt_top1.branch\[1\].mux_I/um_iw[285] tt_top1.branch\[1\].mux_I/um_iw[286] tt_top1.branch\[1\].mux_I/um_iw[287]
+ tt_top1.branch\[1\].mux_I/um_ow[376] tt_top1.branch\[1\].mux_I/um_ow[377] tt_top1.branch\[1\].mux_I/um_ow[378]
+ tt_top1.branch\[1\].mux_I/um_ow[379] tt_top1.branch\[1\].mux_I/um_ow[380] tt_top1.branch\[1\].mux_I/um_ow[381]
+ tt_top1.branch\[1\].mux_I/um_ow[382] tt_top1.branch\[1\].mux_I/um_ow[383] tt_top1.branch\[1\].mux_I/um_ow[368]
+ tt_top1.branch\[1\].mux_I/um_ow[369] tt_top1.branch\[1\].mux_I/um_ow[370] tt_top1.branch\[1\].mux_I/um_ow[371]
+ tt_top1.branch\[1\].mux_I/um_ow[372] tt_top1.branch\[1\].mux_I/um_ow[373] tt_top1.branch\[1\].mux_I/um_ow[374]
+ tt_top1.branch\[1\].mux_I/um_ow[375] tt_top1.branch\[1\].mux_I/um_ow[360] tt_top1.branch\[1\].mux_I/um_ow[361]
+ tt_top1.branch\[1\].mux_I/um_ow[362] tt_top1.branch\[1\].mux_I/um_ow[363] tt_top1.branch\[1\].mux_I/um_ow[364]
+ tt_top1.branch\[1\].mux_I/um_ow[365] tt_top1.branch\[1\].mux_I/um_ow[366] tt_top1.branch\[1\].mux_I/um_ow[367]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[1\].col_um\[1\].um_top_I.block_1_17.tt_um_I tt_top1.branch\[1\].mux_I/um_iw[54]
+ tt_top1.branch\[1\].mux_I/um_ena[3] tt_top1.branch\[1\].mux_I/um_iw[55] tt_top1.branch\[1\].mux_I/um_iw[56]
+ tt_top1.branch\[1\].mux_I/um_iw[57] tt_top1.branch\[1\].mux_I/um_iw[58] tt_top1.branch\[1\].mux_I/um_iw[59]
+ tt_top1.branch\[1\].mux_I/um_iw[60] tt_top1.branch\[1\].mux_I/um_iw[61] tt_top1.branch\[1\].mux_I/um_iw[62]
+ tt_top1.branch\[1\].mux_I/um_iw[63] tt_top1.branch\[1\].mux_I/um_iw[64] tt_top1.branch\[1\].mux_I/um_iw[65]
+ tt_top1.branch\[1\].mux_I/um_iw[66] tt_top1.branch\[1\].mux_I/um_iw[67] tt_top1.branch\[1\].mux_I/um_iw[68]
+ tt_top1.branch\[1\].mux_I/um_iw[69] tt_top1.branch\[1\].mux_I/um_iw[70] tt_top1.branch\[1\].mux_I/um_iw[71]
+ tt_top1.branch\[1\].mux_I/um_ow[88] tt_top1.branch\[1\].mux_I/um_ow[89] tt_top1.branch\[1\].mux_I/um_ow[90]
+ tt_top1.branch\[1\].mux_I/um_ow[91] tt_top1.branch\[1\].mux_I/um_ow[92] tt_top1.branch\[1\].mux_I/um_ow[93]
+ tt_top1.branch\[1\].mux_I/um_ow[94] tt_top1.branch\[1\].mux_I/um_ow[95] tt_top1.branch\[1\].mux_I/um_ow[80]
+ tt_top1.branch\[1\].mux_I/um_ow[81] tt_top1.branch\[1\].mux_I/um_ow[82] tt_top1.branch\[1\].mux_I/um_ow[83]
+ tt_top1.branch\[1\].mux_I/um_ow[84] tt_top1.branch\[1\].mux_I/um_ow[85] tt_top1.branch\[1\].mux_I/um_ow[86]
+ tt_top1.branch\[1\].mux_I/um_ow[87] tt_top1.branch\[1\].mux_I/um_ow[72] tt_top1.branch\[1\].mux_I/um_ow[73]
+ tt_top1.branch\[1\].mux_I/um_ow[74] tt_top1.branch\[1\].mux_I/um_ow[75] tt_top1.branch\[1\].mux_I/um_ow[76]
+ tt_top1.branch\[1\].mux_I/um_ow[77] tt_top1.branch\[1\].mux_I/um_ow[78] tt_top1.branch\[1\].mux_I/um_ow[79]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[1\].col_um\[2\].um_bot_I.block_0_18.tt_um_I tt_top1.branch\[1\].mux_I/um_iw[72]
+ tt_top1.branch\[1\].mux_I/um_ena[4] tt_top1.branch\[1\].mux_I/um_iw[73] tt_top1.branch\[1\].mux_I/um_iw[74]
+ tt_top1.branch\[1\].mux_I/um_iw[75] tt_top1.branch\[1\].mux_I/um_iw[76] tt_top1.branch\[1\].mux_I/um_iw[77]
+ tt_top1.branch\[1\].mux_I/um_iw[78] tt_top1.branch\[1\].mux_I/um_iw[79] tt_top1.branch\[1\].mux_I/um_iw[80]
+ tt_top1.branch\[1\].mux_I/um_iw[81] tt_top1.branch\[1\].mux_I/um_iw[82] tt_top1.branch\[1\].mux_I/um_iw[83]
+ tt_top1.branch\[1\].mux_I/um_iw[84] tt_top1.branch\[1\].mux_I/um_iw[85] tt_top1.branch\[1\].mux_I/um_iw[86]
+ tt_top1.branch\[1\].mux_I/um_iw[87] tt_top1.branch\[1\].mux_I/um_iw[88] tt_top1.branch\[1\].mux_I/um_iw[89]
+ tt_top1.branch\[1\].mux_I/um_ow[112] tt_top1.branch\[1\].mux_I/um_ow[113] tt_top1.branch\[1\].mux_I/um_ow[114]
+ tt_top1.branch\[1\].mux_I/um_ow[115] tt_top1.branch\[1\].mux_I/um_ow[116] tt_top1.branch\[1\].mux_I/um_ow[117]
+ tt_top1.branch\[1\].mux_I/um_ow[118] tt_top1.branch\[1\].mux_I/um_ow[119] tt_top1.branch\[1\].mux_I/um_ow[104]
+ tt_top1.branch\[1\].mux_I/um_ow[105] tt_top1.branch\[1\].mux_I/um_ow[106] tt_top1.branch\[1\].mux_I/um_ow[107]
+ tt_top1.branch\[1\].mux_I/um_ow[108] tt_top1.branch\[1\].mux_I/um_ow[109] tt_top1.branch\[1\].mux_I/um_ow[110]
+ tt_top1.branch\[1\].mux_I/um_ow[111] tt_top1.branch\[1\].mux_I/um_ow[96] tt_top1.branch\[1\].mux_I/um_ow[97]
+ tt_top1.branch\[1\].mux_I/um_ow[98] tt_top1.branch\[1\].mux_I/um_ow[99] tt_top1.branch\[1\].mux_I/um_ow[100]
+ tt_top1.branch\[1\].mux_I/um_ow[101] tt_top1.branch\[1\].mux_I/um_ow[102] tt_top1.branch\[1\].mux_I/um_ow[103]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[0\].col_um\[7\].um_top_I.block_1_7.tt_um_I tt_top1.branch\[0\].mux_I/um_iw[270]
+ tt_top1.branch\[0\].mux_I/um_ena[15] tt_top1.branch\[0\].mux_I/um_iw[271] tt_top1.branch\[0\].mux_I/um_iw[272]
+ tt_top1.branch\[0\].mux_I/um_iw[273] tt_top1.branch\[0\].mux_I/um_iw[274] tt_top1.branch\[0\].mux_I/um_iw[275]
+ tt_top1.branch\[0\].mux_I/um_iw[276] tt_top1.branch\[0\].mux_I/um_iw[277] tt_top1.branch\[0\].mux_I/um_iw[278]
+ tt_top1.branch\[0\].mux_I/um_iw[279] tt_top1.branch\[0\].mux_I/um_iw[280] tt_top1.branch\[0\].mux_I/um_iw[281]
+ tt_top1.branch\[0\].mux_I/um_iw[282] tt_top1.branch\[0\].mux_I/um_iw[283] tt_top1.branch\[0\].mux_I/um_iw[284]
+ tt_top1.branch\[0\].mux_I/um_iw[285] tt_top1.branch\[0\].mux_I/um_iw[286] tt_top1.branch\[0\].mux_I/um_iw[287]
+ tt_top1.branch\[0\].mux_I/um_ow[376] tt_top1.branch\[0\].mux_I/um_ow[377] tt_top1.branch\[0\].mux_I/um_ow[378]
+ tt_top1.branch\[0\].mux_I/um_ow[379] tt_top1.branch\[0\].mux_I/um_ow[380] tt_top1.branch\[0\].mux_I/um_ow[381]
+ tt_top1.branch\[0\].mux_I/um_ow[382] tt_top1.branch\[0\].mux_I/um_ow[383] tt_top1.branch\[0\].mux_I/um_ow[368]
+ tt_top1.branch\[0\].mux_I/um_ow[369] tt_top1.branch\[0\].mux_I/um_ow[370] tt_top1.branch\[0\].mux_I/um_ow[371]
+ tt_top1.branch\[0\].mux_I/um_ow[372] tt_top1.branch\[0\].mux_I/um_ow[373] tt_top1.branch\[0\].mux_I/um_ow[374]
+ tt_top1.branch\[0\].mux_I/um_ow[375] tt_top1.branch\[0\].mux_I/um_ow[360] tt_top1.branch\[0\].mux_I/um_ow[361]
+ tt_top1.branch\[0\].mux_I/um_ow[362] tt_top1.branch\[0\].mux_I/um_ow[363] tt_top1.branch\[0\].mux_I/um_ow[364]
+ tt_top1.branch\[0\].mux_I/um_ow[365] tt_top1.branch\[0\].mux_I/um_ow[366] tt_top1.branch\[0\].mux_I/um_ow[367]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[1\].col_um\[4\].um_top_I.block_1_20.tt_um_I tt_top1.branch\[1\].mux_I/um_iw[162]
+ tt_top1.branch\[1\].mux_I/um_ena[9] tt_top1.branch\[1\].mux_I/um_iw[163] tt_top1.branch\[1\].mux_I/um_iw[164]
+ tt_top1.branch\[1\].mux_I/um_iw[165] tt_top1.branch\[1\].mux_I/um_iw[166] tt_top1.branch\[1\].mux_I/um_iw[167]
+ tt_top1.branch\[1\].mux_I/um_iw[168] tt_top1.branch\[1\].mux_I/um_iw[169] tt_top1.branch\[1\].mux_I/um_iw[170]
+ tt_top1.branch\[1\].mux_I/um_iw[171] tt_top1.branch\[1\].mux_I/um_iw[172] tt_top1.branch\[1\].mux_I/um_iw[173]
+ tt_top1.branch\[1\].mux_I/um_iw[174] tt_top1.branch\[1\].mux_I/um_iw[175] tt_top1.branch\[1\].mux_I/um_iw[176]
+ tt_top1.branch\[1\].mux_I/um_iw[177] tt_top1.branch\[1\].mux_I/um_iw[178] tt_top1.branch\[1\].mux_I/um_iw[179]
+ tt_top1.branch\[1\].mux_I/um_ow[232] tt_top1.branch\[1\].mux_I/um_ow[233] tt_top1.branch\[1\].mux_I/um_ow[234]
+ tt_top1.branch\[1\].mux_I/um_ow[235] tt_top1.branch\[1\].mux_I/um_ow[236] tt_top1.branch\[1\].mux_I/um_ow[237]
+ tt_top1.branch\[1\].mux_I/um_ow[238] tt_top1.branch\[1\].mux_I/um_ow[239] tt_top1.branch\[1\].mux_I/um_ow[224]
+ tt_top1.branch\[1\].mux_I/um_ow[225] tt_top1.branch\[1\].mux_I/um_ow[226] tt_top1.branch\[1\].mux_I/um_ow[227]
+ tt_top1.branch\[1\].mux_I/um_ow[228] tt_top1.branch\[1\].mux_I/um_ow[229] tt_top1.branch\[1\].mux_I/um_ow[230]
+ tt_top1.branch\[1\].mux_I/um_ow[231] tt_top1.branch\[1\].mux_I/um_ow[216] tt_top1.branch\[1\].mux_I/um_ow[217]
+ tt_top1.branch\[1\].mux_I/um_ow[218] tt_top1.branch\[1\].mux_I/um_ow[219] tt_top1.branch\[1\].mux_I/um_ow[220]
+ tt_top1.branch\[1\].mux_I/um_ow[221] tt_top1.branch\[1\].mux_I/um_ow[222] tt_top1.branch\[1\].mux_I/um_ow[223]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[0\].col_um\[6\].um_top_I.block_1_6.tt_um_I tt_top1.branch\[0\].mux_I/um_iw[234]
+ tt_top1.branch\[0\].mux_I/um_ena[13] tt_top1.branch\[0\].mux_I/um_iw[235] tt_top1.branch\[0\].mux_I/um_iw[236]
+ tt_top1.branch\[0\].mux_I/um_iw[237] tt_top1.branch\[0\].mux_I/um_iw[238] tt_top1.branch\[0\].mux_I/um_iw[239]
+ tt_top1.branch\[0\].mux_I/um_iw[240] tt_top1.branch\[0\].mux_I/um_iw[241] tt_top1.branch\[0\].mux_I/um_iw[242]
+ tt_top1.branch\[0\].mux_I/um_iw[243] tt_top1.branch\[0\].mux_I/um_iw[244] tt_top1.branch\[0\].mux_I/um_iw[245]
+ tt_top1.branch\[0\].mux_I/um_iw[246] tt_top1.branch\[0\].mux_I/um_iw[247] tt_top1.branch\[0\].mux_I/um_iw[248]
+ tt_top1.branch\[0\].mux_I/um_iw[249] tt_top1.branch\[0\].mux_I/um_iw[250] tt_top1.branch\[0\].mux_I/um_iw[251]
+ tt_top1.branch\[0\].mux_I/um_ow[328] tt_top1.branch\[0\].mux_I/um_ow[329] tt_top1.branch\[0\].mux_I/um_ow[330]
+ tt_top1.branch\[0\].mux_I/um_ow[331] tt_top1.branch\[0\].mux_I/um_ow[332] tt_top1.branch\[0\].mux_I/um_ow[333]
+ tt_top1.branch\[0\].mux_I/um_ow[334] tt_top1.branch\[0\].mux_I/um_ow[335] tt_top1.branch\[0\].mux_I/um_ow[320]
+ tt_top1.branch\[0\].mux_I/um_ow[321] tt_top1.branch\[0\].mux_I/um_ow[322] tt_top1.branch\[0\].mux_I/um_ow[323]
+ tt_top1.branch\[0\].mux_I/um_ow[324] tt_top1.branch\[0\].mux_I/um_ow[325] tt_top1.branch\[0\].mux_I/um_ow[326]
+ tt_top1.branch\[0\].mux_I/um_ow[327] tt_top1.branch\[0\].mux_I/um_ow[312] tt_top1.branch\[0\].mux_I/um_ow[313]
+ tt_top1.branch\[0\].mux_I/um_ow[314] tt_top1.branch\[0\].mux_I/um_ow[315] tt_top1.branch\[0\].mux_I/um_ow[316]
+ tt_top1.branch\[0\].mux_I/um_ow[317] tt_top1.branch\[0\].mux_I/um_ow[318] tt_top1.branch\[0\].mux_I/um_ow[319]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[1\].col_um\[5\].um_bot_I.block_0_21.tt_um_I tt_top1.branch\[1\].mux_I/um_iw[180]
+ tt_top1.branch\[1\].mux_I/um_ena[10] tt_top1.branch\[1\].mux_I/um_iw[181] tt_top1.branch\[1\].mux_I/um_iw[182]
+ tt_top1.branch\[1\].mux_I/um_iw[183] tt_top1.branch\[1\].mux_I/um_iw[184] tt_top1.branch\[1\].mux_I/um_iw[185]
+ tt_top1.branch\[1\].mux_I/um_iw[186] tt_top1.branch\[1\].mux_I/um_iw[187] tt_top1.branch\[1\].mux_I/um_iw[188]
+ tt_top1.branch\[1\].mux_I/um_iw[189] tt_top1.branch\[1\].mux_I/um_iw[190] tt_top1.branch\[1\].mux_I/um_iw[191]
+ tt_top1.branch\[1\].mux_I/um_iw[192] tt_top1.branch\[1\].mux_I/um_iw[193] tt_top1.branch\[1\].mux_I/um_iw[194]
+ tt_top1.branch\[1\].mux_I/um_iw[195] tt_top1.branch\[1\].mux_I/um_iw[196] tt_top1.branch\[1\].mux_I/um_iw[197]
+ tt_top1.branch\[1\].mux_I/um_ow[256] tt_top1.branch\[1\].mux_I/um_ow[257] tt_top1.branch\[1\].mux_I/um_ow[258]
+ tt_top1.branch\[1\].mux_I/um_ow[259] tt_top1.branch\[1\].mux_I/um_ow[260] tt_top1.branch\[1\].mux_I/um_ow[261]
+ tt_top1.branch\[1\].mux_I/um_ow[262] tt_top1.branch\[1\].mux_I/um_ow[263] tt_top1.branch\[1\].mux_I/um_ow[248]
+ tt_top1.branch\[1\].mux_I/um_ow[249] tt_top1.branch\[1\].mux_I/um_ow[250] tt_top1.branch\[1\].mux_I/um_ow[251]
+ tt_top1.branch\[1\].mux_I/um_ow[252] tt_top1.branch\[1\].mux_I/um_ow[253] tt_top1.branch\[1\].mux_I/um_ow[254]
+ tt_top1.branch\[1\].mux_I/um_ow[255] tt_top1.branch\[1\].mux_I/um_ow[240] tt_top1.branch\[1\].mux_I/um_ow[241]
+ tt_top1.branch\[1\].mux_I/um_ow[242] tt_top1.branch\[1\].mux_I/um_ow[243] tt_top1.branch\[1\].mux_I/um_ow[244]
+ tt_top1.branch\[1\].mux_I/um_ow[245] tt_top1.branch\[1\].mux_I/um_ow[246] tt_top1.branch\[1\].mux_I/um_ow[247]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[0\].col_um\[5\].um_top_I.block_1_5.tt_um_I tt_top1.branch\[0\].mux_I/um_iw[198]
+ tt_top1.branch\[0\].mux_I/um_ena[11] tt_top1.branch\[0\].mux_I/um_iw[199] tt_top1.branch\[0\].mux_I/um_iw[200]
+ tt_top1.branch\[0\].mux_I/um_iw[201] tt_top1.branch\[0\].mux_I/um_iw[202] tt_top1.branch\[0\].mux_I/um_iw[203]
+ tt_top1.branch\[0\].mux_I/um_iw[204] tt_top1.branch\[0\].mux_I/um_iw[205] tt_top1.branch\[0\].mux_I/um_iw[206]
+ tt_top1.branch\[0\].mux_I/um_iw[207] tt_top1.branch\[0\].mux_I/um_iw[208] tt_top1.branch\[0\].mux_I/um_iw[209]
+ tt_top1.branch\[0\].mux_I/um_iw[210] tt_top1.branch\[0\].mux_I/um_iw[211] tt_top1.branch\[0\].mux_I/um_iw[212]
+ tt_top1.branch\[0\].mux_I/um_iw[213] tt_top1.branch\[0\].mux_I/um_iw[214] tt_top1.branch\[0\].mux_I/um_iw[215]
+ tt_top1.branch\[0\].mux_I/um_ow[280] tt_top1.branch\[0\].mux_I/um_ow[281] tt_top1.branch\[0\].mux_I/um_ow[282]
+ tt_top1.branch\[0\].mux_I/um_ow[283] tt_top1.branch\[0\].mux_I/um_ow[284] tt_top1.branch\[0\].mux_I/um_ow[285]
+ tt_top1.branch\[0\].mux_I/um_ow[286] tt_top1.branch\[0\].mux_I/um_ow[287] tt_top1.branch\[0\].mux_I/um_ow[272]
+ tt_top1.branch\[0\].mux_I/um_ow[273] tt_top1.branch\[0\].mux_I/um_ow[274] tt_top1.branch\[0\].mux_I/um_ow[275]
+ tt_top1.branch\[0\].mux_I/um_ow[276] tt_top1.branch\[0\].mux_I/um_ow[277] tt_top1.branch\[0\].mux_I/um_ow[278]
+ tt_top1.branch\[0\].mux_I/um_ow[279] tt_top1.branch\[0\].mux_I/um_ow[264] tt_top1.branch\[0\].mux_I/um_ow[265]
+ tt_top1.branch\[0\].mux_I/um_ow[266] tt_top1.branch\[0\].mux_I/um_ow[267] tt_top1.branch\[0\].mux_I/um_ow[268]
+ tt_top1.branch\[0\].mux_I/um_ow[269] tt_top1.branch\[0\].mux_I/um_ow[270] tt_top1.branch\[0\].mux_I/um_ow[271]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[0\].col_um\[4\].um_top_I.block_1_4.tt_um_I tt_top1.branch\[0\].mux_I/um_iw[162]
+ tt_top1.branch\[0\].mux_I/um_ena[9] tt_top1.branch\[0\].mux_I/um_iw[163] tt_top1.branch\[0\].mux_I/um_iw[164]
+ tt_top1.branch\[0\].mux_I/um_iw[165] tt_top1.branch\[0\].mux_I/um_iw[166] tt_top1.branch\[0\].mux_I/um_iw[167]
+ tt_top1.branch\[0\].mux_I/um_iw[168] tt_top1.branch\[0\].mux_I/um_iw[169] tt_top1.branch\[0\].mux_I/um_iw[170]
+ tt_top1.branch\[0\].mux_I/um_iw[171] tt_top1.branch\[0\].mux_I/um_iw[172] tt_top1.branch\[0\].mux_I/um_iw[173]
+ tt_top1.branch\[0\].mux_I/um_iw[174] tt_top1.branch\[0\].mux_I/um_iw[175] tt_top1.branch\[0\].mux_I/um_iw[176]
+ tt_top1.branch\[0\].mux_I/um_iw[177] tt_top1.branch\[0\].mux_I/um_iw[178] tt_top1.branch\[0\].mux_I/um_iw[179]
+ tt_top1.branch\[0\].mux_I/um_ow[232] tt_top1.branch\[0\].mux_I/um_ow[233] tt_top1.branch\[0\].mux_I/um_ow[234]
+ tt_top1.branch\[0\].mux_I/um_ow[235] tt_top1.branch\[0\].mux_I/um_ow[236] tt_top1.branch\[0\].mux_I/um_ow[237]
+ tt_top1.branch\[0\].mux_I/um_ow[238] tt_top1.branch\[0\].mux_I/um_ow[239] tt_top1.branch\[0\].mux_I/um_ow[224]
+ tt_top1.branch\[0\].mux_I/um_ow[225] tt_top1.branch\[0\].mux_I/um_ow[226] tt_top1.branch\[0\].mux_I/um_ow[227]
+ tt_top1.branch\[0\].mux_I/um_ow[228] tt_top1.branch\[0\].mux_I/um_ow[229] tt_top1.branch\[0\].mux_I/um_ow[230]
+ tt_top1.branch\[0\].mux_I/um_ow[231] tt_top1.branch\[0\].mux_I/um_ow[216] tt_top1.branch\[0\].mux_I/um_ow[217]
+ tt_top1.branch\[0\].mux_I/um_ow[218] tt_top1.branch\[0\].mux_I/um_ow[219] tt_top1.branch\[0\].mux_I/um_ow[220]
+ tt_top1.branch\[0\].mux_I/um_ow[221] tt_top1.branch\[0\].mux_I/um_ow[222] tt_top1.branch\[0\].mux_I/um_ow[223]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[1\].col_um\[3\].um_top_I.block_1_19.tt_um_I tt_top1.branch\[1\].mux_I/um_iw[126]
+ tt_top1.branch\[1\].mux_I/um_ena[7] tt_top1.branch\[1\].mux_I/um_iw[127] tt_top1.branch\[1\].mux_I/um_iw[128]
+ tt_top1.branch\[1\].mux_I/um_iw[129] tt_top1.branch\[1\].mux_I/um_iw[130] tt_top1.branch\[1\].mux_I/um_iw[131]
+ tt_top1.branch\[1\].mux_I/um_iw[132] tt_top1.branch\[1\].mux_I/um_iw[133] tt_top1.branch\[1\].mux_I/um_iw[134]
+ tt_top1.branch\[1\].mux_I/um_iw[135] tt_top1.branch\[1\].mux_I/um_iw[136] tt_top1.branch\[1\].mux_I/um_iw[137]
+ tt_top1.branch\[1\].mux_I/um_iw[138] tt_top1.branch\[1\].mux_I/um_iw[139] tt_top1.branch\[1\].mux_I/um_iw[140]
+ tt_top1.branch\[1\].mux_I/um_iw[141] tt_top1.branch\[1\].mux_I/um_iw[142] tt_top1.branch\[1\].mux_I/um_iw[143]
+ tt_top1.branch\[1\].mux_I/um_ow[184] tt_top1.branch\[1\].mux_I/um_ow[185] tt_top1.branch\[1\].mux_I/um_ow[186]
+ tt_top1.branch\[1\].mux_I/um_ow[187] tt_top1.branch\[1\].mux_I/um_ow[188] tt_top1.branch\[1\].mux_I/um_ow[189]
+ tt_top1.branch\[1\].mux_I/um_ow[190] tt_top1.branch\[1\].mux_I/um_ow[191] tt_top1.branch\[1\].mux_I/um_ow[176]
+ tt_top1.branch\[1\].mux_I/um_ow[177] tt_top1.branch\[1\].mux_I/um_ow[178] tt_top1.branch\[1\].mux_I/um_ow[179]
+ tt_top1.branch\[1\].mux_I/um_ow[180] tt_top1.branch\[1\].mux_I/um_ow[181] tt_top1.branch\[1\].mux_I/um_ow[182]
+ tt_top1.branch\[1\].mux_I/um_ow[183] tt_top1.branch\[1\].mux_I/um_ow[168] tt_top1.branch\[1\].mux_I/um_ow[169]
+ tt_top1.branch\[1\].mux_I/um_ow[170] tt_top1.branch\[1\].mux_I/um_ow[171] tt_top1.branch\[1\].mux_I/um_ow[172]
+ tt_top1.branch\[1\].mux_I/um_ow[173] tt_top1.branch\[1\].mux_I/um_ow[174] tt_top1.branch\[1\].mux_I/um_ow[175]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[0\].col_um\[3\].um_top_I.block_1_3.tt_um_I tt_top1.branch\[0\].mux_I/um_iw[126]
+ tt_top1.branch\[0\].mux_I/um_ena[7] tt_top1.branch\[0\].mux_I/um_iw[127] tt_top1.branch\[0\].mux_I/um_iw[128]
+ tt_top1.branch\[0\].mux_I/um_iw[129] tt_top1.branch\[0\].mux_I/um_iw[130] tt_top1.branch\[0\].mux_I/um_iw[131]
+ tt_top1.branch\[0\].mux_I/um_iw[132] tt_top1.branch\[0\].mux_I/um_iw[133] tt_top1.branch\[0\].mux_I/um_iw[134]
+ tt_top1.branch\[0\].mux_I/um_iw[135] tt_top1.branch\[0\].mux_I/um_iw[136] tt_top1.branch\[0\].mux_I/um_iw[137]
+ tt_top1.branch\[0\].mux_I/um_iw[138] tt_top1.branch\[0\].mux_I/um_iw[139] tt_top1.branch\[0\].mux_I/um_iw[140]
+ tt_top1.branch\[0\].mux_I/um_iw[141] tt_top1.branch\[0\].mux_I/um_iw[142] tt_top1.branch\[0\].mux_I/um_iw[143]
+ tt_top1.branch\[0\].mux_I/um_ow[184] tt_top1.branch\[0\].mux_I/um_ow[185] tt_top1.branch\[0\].mux_I/um_ow[186]
+ tt_top1.branch\[0\].mux_I/um_ow[187] tt_top1.branch\[0\].mux_I/um_ow[188] tt_top1.branch\[0\].mux_I/um_ow[189]
+ tt_top1.branch\[0\].mux_I/um_ow[190] tt_top1.branch\[0\].mux_I/um_ow[191] tt_top1.branch\[0\].mux_I/um_ow[176]
+ tt_top1.branch\[0\].mux_I/um_ow[177] tt_top1.branch\[0\].mux_I/um_ow[178] tt_top1.branch\[0\].mux_I/um_ow[179]
+ tt_top1.branch\[0\].mux_I/um_ow[180] tt_top1.branch\[0\].mux_I/um_ow[181] tt_top1.branch\[0\].mux_I/um_ow[182]
+ tt_top1.branch\[0\].mux_I/um_ow[183] tt_top1.branch\[0\].mux_I/um_ow[168] tt_top1.branch\[0\].mux_I/um_ow[169]
+ tt_top1.branch\[0\].mux_I/um_ow[170] tt_top1.branch\[0\].mux_I/um_ow[171] tt_top1.branch\[0\].mux_I/um_ow[172]
+ tt_top1.branch\[0\].mux_I/um_ow[173] tt_top1.branch\[0\].mux_I/um_ow[174] tt_top1.branch\[0\].mux_I/um_ow[175]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[0\].col_um\[2\].um_top_I.block_1_2.tt_um_I tt_top1.branch\[0\].mux_I/um_iw[90]
+ tt_top1.branch\[0\].mux_I/um_ena[5] tt_top1.branch\[0\].mux_I/um_iw[91] tt_top1.branch\[0\].mux_I/um_iw[92]
+ tt_top1.branch\[0\].mux_I/um_iw[93] tt_top1.branch\[0\].mux_I/um_iw[94] tt_top1.branch\[0\].mux_I/um_iw[95]
+ tt_top1.branch\[0\].mux_I/um_iw[96] tt_top1.branch\[0\].mux_I/um_iw[97] tt_top1.branch\[0\].mux_I/um_iw[98]
+ tt_top1.branch\[0\].mux_I/um_iw[99] tt_top1.branch\[0\].mux_I/um_iw[100] tt_top1.branch\[0\].mux_I/um_iw[101]
+ tt_top1.branch\[0\].mux_I/um_iw[102] tt_top1.branch\[0\].mux_I/um_iw[103] tt_top1.branch\[0\].mux_I/um_iw[104]
+ tt_top1.branch\[0\].mux_I/um_iw[105] tt_top1.branch\[0\].mux_I/um_iw[106] tt_top1.branch\[0\].mux_I/um_iw[107]
+ tt_top1.branch\[0\].mux_I/um_ow[136] tt_top1.branch\[0\].mux_I/um_ow[137] tt_top1.branch\[0\].mux_I/um_ow[138]
+ tt_top1.branch\[0\].mux_I/um_ow[139] tt_top1.branch\[0\].mux_I/um_ow[140] tt_top1.branch\[0\].mux_I/um_ow[141]
+ tt_top1.branch\[0\].mux_I/um_ow[142] tt_top1.branch\[0\].mux_I/um_ow[143] tt_top1.branch\[0\].mux_I/um_ow[128]
+ tt_top1.branch\[0\].mux_I/um_ow[129] tt_top1.branch\[0\].mux_I/um_ow[130] tt_top1.branch\[0\].mux_I/um_ow[131]
+ tt_top1.branch\[0\].mux_I/um_ow[132] tt_top1.branch\[0\].mux_I/um_ow[133] tt_top1.branch\[0\].mux_I/um_ow[134]
+ tt_top1.branch\[0\].mux_I/um_ow[135] tt_top1.branch\[0\].mux_I/um_ow[120] tt_top1.branch\[0\].mux_I/um_ow[121]
+ tt_top1.branch\[0\].mux_I/um_ow[122] tt_top1.branch\[0\].mux_I/um_ow[123] tt_top1.branch\[0\].mux_I/um_ow[124]
+ tt_top1.branch\[0\].mux_I/um_ow[125] tt_top1.branch\[0\].mux_I/um_ow[126] tt_top1.branch\[0\].mux_I/um_ow[127]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[1\].mux_I tt_top1.branch\[1\].mux_I/k_one tt_top1.branch\[1\].mux_I/k_zero
+ tt_top1.branch\[1\].mux_I/k_zero tt_top1.branch\[1\].mux_I/k_zero tt_top1.branch\[1\].mux_I/k_zero
+ tt_top1.branch\[1\].mux_I/k_one tt_top1.branch\[1\].mux_I/k_zero tt_top1.ctrl_I/spine_iw[0]
+ tt_top1.ctrl_I/spine_iw[10] tt_top1.ctrl_I/spine_iw[11] tt_top1.ctrl_I/spine_iw[12]
+ tt_top1.ctrl_I/spine_iw[13] tt_top1.ctrl_I/spine_iw[14] tt_top1.ctrl_I/spine_iw[15]
+ tt_top1.ctrl_I/spine_iw[16] tt_top1.ctrl_I/spine_iw[17] tt_top1.ctrl_I/spine_iw[18]
+ tt_top1.ctrl_I/spine_iw[19] tt_top1.ctrl_I/spine_iw[1] tt_top1.ctrl_I/spine_iw[20]
+ tt_top1.ctrl_I/spine_iw[21] tt_top1.ctrl_I/spine_iw[22] tt_top1.ctrl_I/spine_iw[23]
+ tt_top1.ctrl_I/spine_iw[24] tt_top1.ctrl_I/spine_iw[25] tt_top1.ctrl_I/spine_iw[26]
+ tt_top1.ctrl_I/spine_iw[27] tt_top1.ctrl_I/spine_iw[28] tt_top1.ctrl_I/spine_iw[29]
+ tt_top1.ctrl_I/spine_iw[2] tt_top1.ctrl_I/spine_iw[30] tt_top1.ctrl_I/spine_iw[3]
+ tt_top1.ctrl_I/spine_iw[4] tt_top1.ctrl_I/spine_iw[5] tt_top1.ctrl_I/spine_iw[6]
+ tt_top1.ctrl_I/spine_iw[7] tt_top1.ctrl_I/spine_iw[8] tt_top1.ctrl_I/spine_iw[9]
+ tt_top1.ctrl_I/spine_ow[0] tt_top1.ctrl_I/spine_ow[10] tt_top1.ctrl_I/spine_ow[11]
+ tt_top1.ctrl_I/spine_ow[12] tt_top1.ctrl_I/spine_ow[13] tt_top1.ctrl_I/spine_ow[14]
+ tt_top1.ctrl_I/spine_ow[15] tt_top1.ctrl_I/spine_ow[16] tt_top1.ctrl_I/spine_ow[17]
+ tt_top1.ctrl_I/spine_ow[18] tt_top1.ctrl_I/spine_ow[19] tt_top1.ctrl_I/spine_ow[1]
+ tt_top1.ctrl_I/spine_ow[20] tt_top1.ctrl_I/spine_ow[21] tt_top1.ctrl_I/spine_ow[22]
+ tt_top1.ctrl_I/spine_ow[23] tt_top1.ctrl_I/spine_ow[24] tt_top1.ctrl_I/spine_ow[25]
+ tt_top1.ctrl_I/spine_ow[2] tt_top1.ctrl_I/spine_ow[3] tt_top1.ctrl_I/spine_ow[4]
+ tt_top1.ctrl_I/spine_ow[5] tt_top1.ctrl_I/spine_ow[6] tt_top1.ctrl_I/spine_ow[7]
+ tt_top1.ctrl_I/spine_ow[8] tt_top1.ctrl_I/spine_ow[9] tt_top1.branch\[1\].mux_I/um_ena[0]
+ tt_top1.branch\[1\].mux_I/um_ena[10] tt_top1.branch\[1\].mux_I/um_ena[11] tt_top1.branch\[1\].mux_I/um_ena[12]
+ tt_top1.branch\[1\].mux_I/um_ena[13] tt_top1.branch\[1\].mux_I/um_ena[14] tt_top1.branch\[1\].mux_I/um_ena[15]
+ tt_top1.branch\[1\].mux_I/um_ena[1] tt_top1.branch\[1\].mux_I/um_ena[2] tt_top1.branch\[1\].mux_I/um_ena[3]
+ tt_top1.branch\[1\].mux_I/um_ena[4] tt_top1.branch\[1\].mux_I/um_ena[5] tt_top1.branch\[1\].mux_I/um_ena[6]
+ tt_top1.branch\[1\].mux_I/um_ena[7] tt_top1.branch\[1\].mux_I/um_ena[8] tt_top1.branch\[1\].mux_I/um_ena[9]
+ tt_top1.branch\[1\].mux_I/um_iw[0] tt_top1.branch\[1\].mux_I/um_iw[100] tt_top1.branch\[1\].mux_I/um_iw[101]
+ tt_top1.branch\[1\].mux_I/um_iw[102] tt_top1.branch\[1\].mux_I/um_iw[103] tt_top1.branch\[1\].mux_I/um_iw[104]
+ tt_top1.branch\[1\].mux_I/um_iw[105] tt_top1.branch\[1\].mux_I/um_iw[106] tt_top1.branch\[1\].mux_I/um_iw[107]
+ tt_top1.branch\[1\].mux_I/um_iw[108] tt_top1.branch\[1\].mux_I/um_iw[109] tt_top1.branch\[1\].mux_I/um_iw[10]
+ tt_top1.branch\[1\].mux_I/um_iw[110] tt_top1.branch\[1\].mux_I/um_iw[111] tt_top1.branch\[1\].mux_I/um_iw[112]
+ tt_top1.branch\[1\].mux_I/um_iw[113] tt_top1.branch\[1\].mux_I/um_iw[114] tt_top1.branch\[1\].mux_I/um_iw[115]
+ tt_top1.branch\[1\].mux_I/um_iw[116] tt_top1.branch\[1\].mux_I/um_iw[117] tt_top1.branch\[1\].mux_I/um_iw[118]
+ tt_top1.branch\[1\].mux_I/um_iw[119] tt_top1.branch\[1\].mux_I/um_iw[11] tt_top1.branch\[1\].mux_I/um_iw[120]
+ tt_top1.branch\[1\].mux_I/um_iw[121] tt_top1.branch\[1\].mux_I/um_iw[122] tt_top1.branch\[1\].mux_I/um_iw[123]
+ tt_top1.branch\[1\].mux_I/um_iw[124] tt_top1.branch\[1\].mux_I/um_iw[125] tt_top1.branch\[1\].mux_I/um_iw[126]
+ tt_top1.branch\[1\].mux_I/um_iw[127] tt_top1.branch\[1\].mux_I/um_iw[128] tt_top1.branch\[1\].mux_I/um_iw[129]
+ tt_top1.branch\[1\].mux_I/um_iw[12] tt_top1.branch\[1\].mux_I/um_iw[130] tt_top1.branch\[1\].mux_I/um_iw[131]
+ tt_top1.branch\[1\].mux_I/um_iw[132] tt_top1.branch\[1\].mux_I/um_iw[133] tt_top1.branch\[1\].mux_I/um_iw[134]
+ tt_top1.branch\[1\].mux_I/um_iw[135] tt_top1.branch\[1\].mux_I/um_iw[136] tt_top1.branch\[1\].mux_I/um_iw[137]
+ tt_top1.branch\[1\].mux_I/um_iw[138] tt_top1.branch\[1\].mux_I/um_iw[139] tt_top1.branch\[1\].mux_I/um_iw[13]
+ tt_top1.branch\[1\].mux_I/um_iw[140] tt_top1.branch\[1\].mux_I/um_iw[141] tt_top1.branch\[1\].mux_I/um_iw[142]
+ tt_top1.branch\[1\].mux_I/um_iw[143] tt_top1.branch\[1\].mux_I/um_iw[144] tt_top1.branch\[1\].mux_I/um_iw[145]
+ tt_top1.branch\[1\].mux_I/um_iw[146] tt_top1.branch\[1\].mux_I/um_iw[147] tt_top1.branch\[1\].mux_I/um_iw[148]
+ tt_top1.branch\[1\].mux_I/um_iw[149] tt_top1.branch\[1\].mux_I/um_iw[14] tt_top1.branch\[1\].mux_I/um_iw[150]
+ tt_top1.branch\[1\].mux_I/um_iw[151] tt_top1.branch\[1\].mux_I/um_iw[152] tt_top1.branch\[1\].mux_I/um_iw[153]
+ tt_top1.branch\[1\].mux_I/um_iw[154] tt_top1.branch\[1\].mux_I/um_iw[155] tt_top1.branch\[1\].mux_I/um_iw[156]
+ tt_top1.branch\[1\].mux_I/um_iw[157] tt_top1.branch\[1\].mux_I/um_iw[158] tt_top1.branch\[1\].mux_I/um_iw[159]
+ tt_top1.branch\[1\].mux_I/um_iw[15] tt_top1.branch\[1\].mux_I/um_iw[160] tt_top1.branch\[1\].mux_I/um_iw[161]
+ tt_top1.branch\[1\].mux_I/um_iw[162] tt_top1.branch\[1\].mux_I/um_iw[163] tt_top1.branch\[1\].mux_I/um_iw[164]
+ tt_top1.branch\[1\].mux_I/um_iw[165] tt_top1.branch\[1\].mux_I/um_iw[166] tt_top1.branch\[1\].mux_I/um_iw[167]
+ tt_top1.branch\[1\].mux_I/um_iw[168] tt_top1.branch\[1\].mux_I/um_iw[169] tt_top1.branch\[1\].mux_I/um_iw[16]
+ tt_top1.branch\[1\].mux_I/um_iw[170] tt_top1.branch\[1\].mux_I/um_iw[171] tt_top1.branch\[1\].mux_I/um_iw[172]
+ tt_top1.branch\[1\].mux_I/um_iw[173] tt_top1.branch\[1\].mux_I/um_iw[174] tt_top1.branch\[1\].mux_I/um_iw[175]
+ tt_top1.branch\[1\].mux_I/um_iw[176] tt_top1.branch\[1\].mux_I/um_iw[177] tt_top1.branch\[1\].mux_I/um_iw[178]
+ tt_top1.branch\[1\].mux_I/um_iw[179] tt_top1.branch\[1\].mux_I/um_iw[17] tt_top1.branch\[1\].mux_I/um_iw[180]
+ tt_top1.branch\[1\].mux_I/um_iw[181] tt_top1.branch\[1\].mux_I/um_iw[182] tt_top1.branch\[1\].mux_I/um_iw[183]
+ tt_top1.branch\[1\].mux_I/um_iw[184] tt_top1.branch\[1\].mux_I/um_iw[185] tt_top1.branch\[1\].mux_I/um_iw[186]
+ tt_top1.branch\[1\].mux_I/um_iw[187] tt_top1.branch\[1\].mux_I/um_iw[188] tt_top1.branch\[1\].mux_I/um_iw[189]
+ tt_top1.branch\[1\].mux_I/um_iw[18] tt_top1.branch\[1\].mux_I/um_iw[190] tt_top1.branch\[1\].mux_I/um_iw[191]
+ tt_top1.branch\[1\].mux_I/um_iw[192] tt_top1.branch\[1\].mux_I/um_iw[193] tt_top1.branch\[1\].mux_I/um_iw[194]
+ tt_top1.branch\[1\].mux_I/um_iw[195] tt_top1.branch\[1\].mux_I/um_iw[196] tt_top1.branch\[1\].mux_I/um_iw[197]
+ tt_top1.branch\[1\].mux_I/um_iw[198] tt_top1.branch\[1\].mux_I/um_iw[199] tt_top1.branch\[1\].mux_I/um_iw[19]
+ tt_top1.branch\[1\].mux_I/um_iw[1] tt_top1.branch\[1\].mux_I/um_iw[200] tt_top1.branch\[1\].mux_I/um_iw[201]
+ tt_top1.branch\[1\].mux_I/um_iw[202] tt_top1.branch\[1\].mux_I/um_iw[203] tt_top1.branch\[1\].mux_I/um_iw[204]
+ tt_top1.branch\[1\].mux_I/um_iw[205] tt_top1.branch\[1\].mux_I/um_iw[206] tt_top1.branch\[1\].mux_I/um_iw[207]
+ tt_top1.branch\[1\].mux_I/um_iw[208] tt_top1.branch\[1\].mux_I/um_iw[209] tt_top1.branch\[1\].mux_I/um_iw[20]
+ tt_top1.branch\[1\].mux_I/um_iw[210] tt_top1.branch\[1\].mux_I/um_iw[211] tt_top1.branch\[1\].mux_I/um_iw[212]
+ tt_top1.branch\[1\].mux_I/um_iw[213] tt_top1.branch\[1\].mux_I/um_iw[214] tt_top1.branch\[1\].mux_I/um_iw[215]
+ tt_top1.branch\[1\].mux_I/um_iw[216] tt_top1.branch\[1\].mux_I/um_iw[217] tt_top1.branch\[1\].mux_I/um_iw[218]
+ tt_top1.branch\[1\].mux_I/um_iw[219] tt_top1.branch\[1\].mux_I/um_iw[21] tt_top1.branch\[1\].mux_I/um_iw[220]
+ tt_top1.branch\[1\].mux_I/um_iw[221] tt_top1.branch\[1\].mux_I/um_iw[222] tt_top1.branch\[1\].mux_I/um_iw[223]
+ tt_top1.branch\[1\].mux_I/um_iw[224] tt_top1.branch\[1\].mux_I/um_iw[225] tt_top1.branch\[1\].mux_I/um_iw[226]
+ tt_top1.branch\[1\].mux_I/um_iw[227] tt_top1.branch\[1\].mux_I/um_iw[228] tt_top1.branch\[1\].mux_I/um_iw[229]
+ tt_top1.branch\[1\].mux_I/um_iw[22] tt_top1.branch\[1\].mux_I/um_iw[230] tt_top1.branch\[1\].mux_I/um_iw[231]
+ tt_top1.branch\[1\].mux_I/um_iw[232] tt_top1.branch\[1\].mux_I/um_iw[233] tt_top1.branch\[1\].mux_I/um_iw[234]
+ tt_top1.branch\[1\].mux_I/um_iw[235] tt_top1.branch\[1\].mux_I/um_iw[236] tt_top1.branch\[1\].mux_I/um_iw[237]
+ tt_top1.branch\[1\].mux_I/um_iw[238] tt_top1.branch\[1\].mux_I/um_iw[239] tt_top1.branch\[1\].mux_I/um_iw[23]
+ tt_top1.branch\[1\].mux_I/um_iw[240] tt_top1.branch\[1\].mux_I/um_iw[241] tt_top1.branch\[1\].mux_I/um_iw[242]
+ tt_top1.branch\[1\].mux_I/um_iw[243] tt_top1.branch\[1\].mux_I/um_iw[244] tt_top1.branch\[1\].mux_I/um_iw[245]
+ tt_top1.branch\[1\].mux_I/um_iw[246] tt_top1.branch\[1\].mux_I/um_iw[247] tt_top1.branch\[1\].mux_I/um_iw[248]
+ tt_top1.branch\[1\].mux_I/um_iw[249] tt_top1.branch\[1\].mux_I/um_iw[24] tt_top1.branch\[1\].mux_I/um_iw[250]
+ tt_top1.branch\[1\].mux_I/um_iw[251] tt_top1.branch\[1\].mux_I/um_iw[252] tt_top1.branch\[1\].mux_I/um_iw[253]
+ tt_top1.branch\[1\].mux_I/um_iw[254] tt_top1.branch\[1\].mux_I/um_iw[255] tt_top1.branch\[1\].mux_I/um_iw[256]
+ tt_top1.branch\[1\].mux_I/um_iw[257] tt_top1.branch\[1\].mux_I/um_iw[258] tt_top1.branch\[1\].mux_I/um_iw[259]
+ tt_top1.branch\[1\].mux_I/um_iw[25] tt_top1.branch\[1\].mux_I/um_iw[260] tt_top1.branch\[1\].mux_I/um_iw[261]
+ tt_top1.branch\[1\].mux_I/um_iw[262] tt_top1.branch\[1\].mux_I/um_iw[263] tt_top1.branch\[1\].mux_I/um_iw[264]
+ tt_top1.branch\[1\].mux_I/um_iw[265] tt_top1.branch\[1\].mux_I/um_iw[266] tt_top1.branch\[1\].mux_I/um_iw[267]
+ tt_top1.branch\[1\].mux_I/um_iw[268] tt_top1.branch\[1\].mux_I/um_iw[269] tt_top1.branch\[1\].mux_I/um_iw[26]
+ tt_top1.branch\[1\].mux_I/um_iw[270] tt_top1.branch\[1\].mux_I/um_iw[271] tt_top1.branch\[1\].mux_I/um_iw[272]
+ tt_top1.branch\[1\].mux_I/um_iw[273] tt_top1.branch\[1\].mux_I/um_iw[274] tt_top1.branch\[1\].mux_I/um_iw[275]
+ tt_top1.branch\[1\].mux_I/um_iw[276] tt_top1.branch\[1\].mux_I/um_iw[277] tt_top1.branch\[1\].mux_I/um_iw[278]
+ tt_top1.branch\[1\].mux_I/um_iw[279] tt_top1.branch\[1\].mux_I/um_iw[27] tt_top1.branch\[1\].mux_I/um_iw[280]
+ tt_top1.branch\[1\].mux_I/um_iw[281] tt_top1.branch\[1\].mux_I/um_iw[282] tt_top1.branch\[1\].mux_I/um_iw[283]
+ tt_top1.branch\[1\].mux_I/um_iw[284] tt_top1.branch\[1\].mux_I/um_iw[285] tt_top1.branch\[1\].mux_I/um_iw[286]
+ tt_top1.branch\[1\].mux_I/um_iw[287] tt_top1.branch\[1\].mux_I/um_iw[28] tt_top1.branch\[1\].mux_I/um_iw[29]
+ tt_top1.branch\[1\].mux_I/um_iw[2] tt_top1.branch\[1\].mux_I/um_iw[30] tt_top1.branch\[1\].mux_I/um_iw[31]
+ tt_top1.branch\[1\].mux_I/um_iw[32] tt_top1.branch\[1\].mux_I/um_iw[33] tt_top1.branch\[1\].mux_I/um_iw[34]
+ tt_top1.branch\[1\].mux_I/um_iw[35] tt_top1.branch\[1\].mux_I/um_iw[36] tt_top1.branch\[1\].mux_I/um_iw[37]
+ tt_top1.branch\[1\].mux_I/um_iw[38] tt_top1.branch\[1\].mux_I/um_iw[39] tt_top1.branch\[1\].mux_I/um_iw[3]
+ tt_top1.branch\[1\].mux_I/um_iw[40] tt_top1.branch\[1\].mux_I/um_iw[41] tt_top1.branch\[1\].mux_I/um_iw[42]
+ tt_top1.branch\[1\].mux_I/um_iw[43] tt_top1.branch\[1\].mux_I/um_iw[44] tt_top1.branch\[1\].mux_I/um_iw[45]
+ tt_top1.branch\[1\].mux_I/um_iw[46] tt_top1.branch\[1\].mux_I/um_iw[47] tt_top1.branch\[1\].mux_I/um_iw[48]
+ tt_top1.branch\[1\].mux_I/um_iw[49] tt_top1.branch\[1\].mux_I/um_iw[4] tt_top1.branch\[1\].mux_I/um_iw[50]
+ tt_top1.branch\[1\].mux_I/um_iw[51] tt_top1.branch\[1\].mux_I/um_iw[52] tt_top1.branch\[1\].mux_I/um_iw[53]
+ tt_top1.branch\[1\].mux_I/um_iw[54] tt_top1.branch\[1\].mux_I/um_iw[55] tt_top1.branch\[1\].mux_I/um_iw[56]
+ tt_top1.branch\[1\].mux_I/um_iw[57] tt_top1.branch\[1\].mux_I/um_iw[58] tt_top1.branch\[1\].mux_I/um_iw[59]
+ tt_top1.branch\[1\].mux_I/um_iw[5] tt_top1.branch\[1\].mux_I/um_iw[60] tt_top1.branch\[1\].mux_I/um_iw[61]
+ tt_top1.branch\[1\].mux_I/um_iw[62] tt_top1.branch\[1\].mux_I/um_iw[63] tt_top1.branch\[1\].mux_I/um_iw[64]
+ tt_top1.branch\[1\].mux_I/um_iw[65] tt_top1.branch\[1\].mux_I/um_iw[66] tt_top1.branch\[1\].mux_I/um_iw[67]
+ tt_top1.branch\[1\].mux_I/um_iw[68] tt_top1.branch\[1\].mux_I/um_iw[69] tt_top1.branch\[1\].mux_I/um_iw[6]
+ tt_top1.branch\[1\].mux_I/um_iw[70] tt_top1.branch\[1\].mux_I/um_iw[71] tt_top1.branch\[1\].mux_I/um_iw[72]
+ tt_top1.branch\[1\].mux_I/um_iw[73] tt_top1.branch\[1\].mux_I/um_iw[74] tt_top1.branch\[1\].mux_I/um_iw[75]
+ tt_top1.branch\[1\].mux_I/um_iw[76] tt_top1.branch\[1\].mux_I/um_iw[77] tt_top1.branch\[1\].mux_I/um_iw[78]
+ tt_top1.branch\[1\].mux_I/um_iw[79] tt_top1.branch\[1\].mux_I/um_iw[7] tt_top1.branch\[1\].mux_I/um_iw[80]
+ tt_top1.branch\[1\].mux_I/um_iw[81] tt_top1.branch\[1\].mux_I/um_iw[82] tt_top1.branch\[1\].mux_I/um_iw[83]
+ tt_top1.branch\[1\].mux_I/um_iw[84] tt_top1.branch\[1\].mux_I/um_iw[85] tt_top1.branch\[1\].mux_I/um_iw[86]
+ tt_top1.branch\[1\].mux_I/um_iw[87] tt_top1.branch\[1\].mux_I/um_iw[88] tt_top1.branch\[1\].mux_I/um_iw[89]
+ tt_top1.branch\[1\].mux_I/um_iw[8] tt_top1.branch\[1\].mux_I/um_iw[90] tt_top1.branch\[1\].mux_I/um_iw[91]
+ tt_top1.branch\[1\].mux_I/um_iw[92] tt_top1.branch\[1\].mux_I/um_iw[93] tt_top1.branch\[1\].mux_I/um_iw[94]
+ tt_top1.branch\[1\].mux_I/um_iw[95] tt_top1.branch\[1\].mux_I/um_iw[96] tt_top1.branch\[1\].mux_I/um_iw[97]
+ tt_top1.branch\[1\].mux_I/um_iw[98] tt_top1.branch\[1\].mux_I/um_iw[99] tt_top1.branch\[1\].mux_I/um_iw[9]
+ tt_top1.branch\[1\].mux_I/um_k_zero[0] tt_top1.branch\[1\].mux_I/um_k_zero[10] tt_top1.branch\[1\].mux_I/um_k_zero[11]
+ tt_top1.branch\[1\].mux_I/um_k_zero[12] tt_top1.branch\[1\].mux_I/um_k_zero[13]
+ tt_top1.branch\[1\].mux_I/um_k_zero[14] tt_top1.branch\[1\].mux_I/um_k_zero[15]
+ tt_top1.branch\[1\].mux_I/um_k_zero[1] tt_top1.branch\[1\].mux_I/um_k_zero[2] tt_top1.branch\[1\].mux_I/um_k_zero[3]
+ tt_top1.branch\[1\].mux_I/um_k_zero[4] tt_top1.branch\[1\].mux_I/um_k_zero[5] tt_top1.branch\[1\].mux_I/um_k_zero[6]
+ tt_top1.branch\[1\].mux_I/um_k_zero[7] tt_top1.branch\[1\].mux_I/um_k_zero[8] tt_top1.branch\[1\].mux_I/um_k_zero[9]
+ tt_top1.branch\[1\].mux_I/um_ow[0] tt_top1.branch\[1\].mux_I/um_ow[100] tt_top1.branch\[1\].mux_I/um_ow[101]
+ tt_top1.branch\[1\].mux_I/um_ow[102] tt_top1.branch\[1\].mux_I/um_ow[103] tt_top1.branch\[1\].mux_I/um_ow[104]
+ tt_top1.branch\[1\].mux_I/um_ow[105] tt_top1.branch\[1\].mux_I/um_ow[106] tt_top1.branch\[1\].mux_I/um_ow[107]
+ tt_top1.branch\[1\].mux_I/um_ow[108] tt_top1.branch\[1\].mux_I/um_ow[109] tt_top1.branch\[1\].mux_I/um_ow[10]
+ tt_top1.branch\[1\].mux_I/um_ow[110] tt_top1.branch\[1\].mux_I/um_ow[111] tt_top1.branch\[1\].mux_I/um_ow[112]
+ tt_top1.branch\[1\].mux_I/um_ow[113] tt_top1.branch\[1\].mux_I/um_ow[114] tt_top1.branch\[1\].mux_I/um_ow[115]
+ tt_top1.branch\[1\].mux_I/um_ow[116] tt_top1.branch\[1\].mux_I/um_ow[117] tt_top1.branch\[1\].mux_I/um_ow[118]
+ tt_top1.branch\[1\].mux_I/um_ow[119] tt_top1.branch\[1\].mux_I/um_ow[11] tt_top1.branch\[1\].mux_I/um_ow[120]
+ tt_top1.branch\[1\].mux_I/um_ow[121] tt_top1.branch\[1\].mux_I/um_ow[122] tt_top1.branch\[1\].mux_I/um_ow[123]
+ tt_top1.branch\[1\].mux_I/um_ow[124] tt_top1.branch\[1\].mux_I/um_ow[125] tt_top1.branch\[1\].mux_I/um_ow[126]
+ tt_top1.branch\[1\].mux_I/um_ow[127] tt_top1.branch\[1\].mux_I/um_ow[128] tt_top1.branch\[1\].mux_I/um_ow[129]
+ tt_top1.branch\[1\].mux_I/um_ow[12] tt_top1.branch\[1\].mux_I/um_ow[130] tt_top1.branch\[1\].mux_I/um_ow[131]
+ tt_top1.branch\[1\].mux_I/um_ow[132] tt_top1.branch\[1\].mux_I/um_ow[133] tt_top1.branch\[1\].mux_I/um_ow[134]
+ tt_top1.branch\[1\].mux_I/um_ow[135] tt_top1.branch\[1\].mux_I/um_ow[136] tt_top1.branch\[1\].mux_I/um_ow[137]
+ tt_top1.branch\[1\].mux_I/um_ow[138] tt_top1.branch\[1\].mux_I/um_ow[139] tt_top1.branch\[1\].mux_I/um_ow[13]
+ tt_top1.branch\[1\].mux_I/um_ow[140] tt_top1.branch\[1\].mux_I/um_ow[141] tt_top1.branch\[1\].mux_I/um_ow[142]
+ tt_top1.branch\[1\].mux_I/um_ow[143] tt_top1.branch\[1\].mux_I/um_ow[144] tt_top1.branch\[1\].mux_I/um_ow[145]
+ tt_top1.branch\[1\].mux_I/um_ow[146] tt_top1.branch\[1\].mux_I/um_ow[147] tt_top1.branch\[1\].mux_I/um_ow[148]
+ tt_top1.branch\[1\].mux_I/um_ow[149] tt_top1.branch\[1\].mux_I/um_ow[14] tt_top1.branch\[1\].mux_I/um_ow[150]
+ tt_top1.branch\[1\].mux_I/um_ow[151] tt_top1.branch\[1\].mux_I/um_ow[152] tt_top1.branch\[1\].mux_I/um_ow[153]
+ tt_top1.branch\[1\].mux_I/um_ow[154] tt_top1.branch\[1\].mux_I/um_ow[155] tt_top1.branch\[1\].mux_I/um_ow[156]
+ tt_top1.branch\[1\].mux_I/um_ow[157] tt_top1.branch\[1\].mux_I/um_ow[158] tt_top1.branch\[1\].mux_I/um_ow[159]
+ tt_top1.branch\[1\].mux_I/um_ow[15] tt_top1.branch\[1\].mux_I/um_ow[160] tt_top1.branch\[1\].mux_I/um_ow[161]
+ tt_top1.branch\[1\].mux_I/um_ow[162] tt_top1.branch\[1\].mux_I/um_ow[163] tt_top1.branch\[1\].mux_I/um_ow[164]
+ tt_top1.branch\[1\].mux_I/um_ow[165] tt_top1.branch\[1\].mux_I/um_ow[166] tt_top1.branch\[1\].mux_I/um_ow[167]
+ tt_top1.branch\[1\].mux_I/um_ow[168] tt_top1.branch\[1\].mux_I/um_ow[169] tt_top1.branch\[1\].mux_I/um_ow[16]
+ tt_top1.branch\[1\].mux_I/um_ow[170] tt_top1.branch\[1\].mux_I/um_ow[171] tt_top1.branch\[1\].mux_I/um_ow[172]
+ tt_top1.branch\[1\].mux_I/um_ow[173] tt_top1.branch\[1\].mux_I/um_ow[174] tt_top1.branch\[1\].mux_I/um_ow[175]
+ tt_top1.branch\[1\].mux_I/um_ow[176] tt_top1.branch\[1\].mux_I/um_ow[177] tt_top1.branch\[1\].mux_I/um_ow[178]
+ tt_top1.branch\[1\].mux_I/um_ow[179] tt_top1.branch\[1\].mux_I/um_ow[17] tt_top1.branch\[1\].mux_I/um_ow[180]
+ tt_top1.branch\[1\].mux_I/um_ow[181] tt_top1.branch\[1\].mux_I/um_ow[182] tt_top1.branch\[1\].mux_I/um_ow[183]
+ tt_top1.branch\[1\].mux_I/um_ow[184] tt_top1.branch\[1\].mux_I/um_ow[185] tt_top1.branch\[1\].mux_I/um_ow[186]
+ tt_top1.branch\[1\].mux_I/um_ow[187] tt_top1.branch\[1\].mux_I/um_ow[188] tt_top1.branch\[1\].mux_I/um_ow[189]
+ tt_top1.branch\[1\].mux_I/um_ow[18] tt_top1.branch\[1\].mux_I/um_ow[190] tt_top1.branch\[1\].mux_I/um_ow[191]
+ tt_top1.branch\[1\].mux_I/um_ow[192] tt_top1.branch\[1\].mux_I/um_ow[193] tt_top1.branch\[1\].mux_I/um_ow[194]
+ tt_top1.branch\[1\].mux_I/um_ow[195] tt_top1.branch\[1\].mux_I/um_ow[196] tt_top1.branch\[1\].mux_I/um_ow[197]
+ tt_top1.branch\[1\].mux_I/um_ow[198] tt_top1.branch\[1\].mux_I/um_ow[199] tt_top1.branch\[1\].mux_I/um_ow[19]
+ tt_top1.branch\[1\].mux_I/um_ow[1] tt_top1.branch\[1\].mux_I/um_ow[200] tt_top1.branch\[1\].mux_I/um_ow[201]
+ tt_top1.branch\[1\].mux_I/um_ow[202] tt_top1.branch\[1\].mux_I/um_ow[203] tt_top1.branch\[1\].mux_I/um_ow[204]
+ tt_top1.branch\[1\].mux_I/um_ow[205] tt_top1.branch\[1\].mux_I/um_ow[206] tt_top1.branch\[1\].mux_I/um_ow[207]
+ tt_top1.branch\[1\].mux_I/um_ow[208] tt_top1.branch\[1\].mux_I/um_ow[209] tt_top1.branch\[1\].mux_I/um_ow[20]
+ tt_top1.branch\[1\].mux_I/um_ow[210] tt_top1.branch\[1\].mux_I/um_ow[211] tt_top1.branch\[1\].mux_I/um_ow[212]
+ tt_top1.branch\[1\].mux_I/um_ow[213] tt_top1.branch\[1\].mux_I/um_ow[214] tt_top1.branch\[1\].mux_I/um_ow[215]
+ tt_top1.branch\[1\].mux_I/um_ow[216] tt_top1.branch\[1\].mux_I/um_ow[217] tt_top1.branch\[1\].mux_I/um_ow[218]
+ tt_top1.branch\[1\].mux_I/um_ow[219] tt_top1.branch\[1\].mux_I/um_ow[21] tt_top1.branch\[1\].mux_I/um_ow[220]
+ tt_top1.branch\[1\].mux_I/um_ow[221] tt_top1.branch\[1\].mux_I/um_ow[222] tt_top1.branch\[1\].mux_I/um_ow[223]
+ tt_top1.branch\[1\].mux_I/um_ow[224] tt_top1.branch\[1\].mux_I/um_ow[225] tt_top1.branch\[1\].mux_I/um_ow[226]
+ tt_top1.branch\[1\].mux_I/um_ow[227] tt_top1.branch\[1\].mux_I/um_ow[228] tt_top1.branch\[1\].mux_I/um_ow[229]
+ tt_top1.branch\[1\].mux_I/um_ow[22] tt_top1.branch\[1\].mux_I/um_ow[230] tt_top1.branch\[1\].mux_I/um_ow[231]
+ tt_top1.branch\[1\].mux_I/um_ow[232] tt_top1.branch\[1\].mux_I/um_ow[233] tt_top1.branch\[1\].mux_I/um_ow[234]
+ tt_top1.branch\[1\].mux_I/um_ow[235] tt_top1.branch\[1\].mux_I/um_ow[236] tt_top1.branch\[1\].mux_I/um_ow[237]
+ tt_top1.branch\[1\].mux_I/um_ow[238] tt_top1.branch\[1\].mux_I/um_ow[239] tt_top1.branch\[1\].mux_I/um_ow[23]
+ tt_top1.branch\[1\].mux_I/um_ow[240] tt_top1.branch\[1\].mux_I/um_ow[241] tt_top1.branch\[1\].mux_I/um_ow[242]
+ tt_top1.branch\[1\].mux_I/um_ow[243] tt_top1.branch\[1\].mux_I/um_ow[244] tt_top1.branch\[1\].mux_I/um_ow[245]
+ tt_top1.branch\[1\].mux_I/um_ow[246] tt_top1.branch\[1\].mux_I/um_ow[247] tt_top1.branch\[1\].mux_I/um_ow[248]
+ tt_top1.branch\[1\].mux_I/um_ow[249] tt_top1.branch\[1\].mux_I/um_ow[24] tt_top1.branch\[1\].mux_I/um_ow[250]
+ tt_top1.branch\[1\].mux_I/um_ow[251] tt_top1.branch\[1\].mux_I/um_ow[252] tt_top1.branch\[1\].mux_I/um_ow[253]
+ tt_top1.branch\[1\].mux_I/um_ow[254] tt_top1.branch\[1\].mux_I/um_ow[255] tt_top1.branch\[1\].mux_I/um_ow[256]
+ tt_top1.branch\[1\].mux_I/um_ow[257] tt_top1.branch\[1\].mux_I/um_ow[258] tt_top1.branch\[1\].mux_I/um_ow[259]
+ tt_top1.branch\[1\].mux_I/um_ow[25] tt_top1.branch\[1\].mux_I/um_ow[260] tt_top1.branch\[1\].mux_I/um_ow[261]
+ tt_top1.branch\[1\].mux_I/um_ow[262] tt_top1.branch\[1\].mux_I/um_ow[263] tt_top1.branch\[1\].mux_I/um_ow[264]
+ tt_top1.branch\[1\].mux_I/um_ow[265] tt_top1.branch\[1\].mux_I/um_ow[266] tt_top1.branch\[1\].mux_I/um_ow[267]
+ tt_top1.branch\[1\].mux_I/um_ow[268] tt_top1.branch\[1\].mux_I/um_ow[269] tt_top1.branch\[1\].mux_I/um_ow[26]
+ tt_top1.branch\[1\].mux_I/um_ow[270] tt_top1.branch\[1\].mux_I/um_ow[271] tt_top1.branch\[1\].mux_I/um_ow[272]
+ tt_top1.branch\[1\].mux_I/um_ow[273] tt_top1.branch\[1\].mux_I/um_ow[274] tt_top1.branch\[1\].mux_I/um_ow[275]
+ tt_top1.branch\[1\].mux_I/um_ow[276] tt_top1.branch\[1\].mux_I/um_ow[277] tt_top1.branch\[1\].mux_I/um_ow[278]
+ tt_top1.branch\[1\].mux_I/um_ow[279] tt_top1.branch\[1\].mux_I/um_ow[27] tt_top1.branch\[1\].mux_I/um_ow[280]
+ tt_top1.branch\[1\].mux_I/um_ow[281] tt_top1.branch\[1\].mux_I/um_ow[282] tt_top1.branch\[1\].mux_I/um_ow[283]
+ tt_top1.branch\[1\].mux_I/um_ow[284] tt_top1.branch\[1\].mux_I/um_ow[285] tt_top1.branch\[1\].mux_I/um_ow[286]
+ tt_top1.branch\[1\].mux_I/um_ow[287] tt_top1.branch\[1\].mux_I/um_ow[288] tt_top1.branch\[1\].mux_I/um_ow[289]
+ tt_top1.branch\[1\].mux_I/um_ow[28] tt_top1.branch\[1\].mux_I/um_ow[290] tt_top1.branch\[1\].mux_I/um_ow[291]
+ tt_top1.branch\[1\].mux_I/um_ow[292] tt_top1.branch\[1\].mux_I/um_ow[293] tt_top1.branch\[1\].mux_I/um_ow[294]
+ tt_top1.branch\[1\].mux_I/um_ow[295] tt_top1.branch\[1\].mux_I/um_ow[296] tt_top1.branch\[1\].mux_I/um_ow[297]
+ tt_top1.branch\[1\].mux_I/um_ow[298] tt_top1.branch\[1\].mux_I/um_ow[299] tt_top1.branch\[1\].mux_I/um_ow[29]
+ tt_top1.branch\[1\].mux_I/um_ow[2] tt_top1.branch\[1\].mux_I/um_ow[300] tt_top1.branch\[1\].mux_I/um_ow[301]
+ tt_top1.branch\[1\].mux_I/um_ow[302] tt_top1.branch\[1\].mux_I/um_ow[303] tt_top1.branch\[1\].mux_I/um_ow[304]
+ tt_top1.branch\[1\].mux_I/um_ow[305] tt_top1.branch\[1\].mux_I/um_ow[306] tt_top1.branch\[1\].mux_I/um_ow[307]
+ tt_top1.branch\[1\].mux_I/um_ow[308] tt_top1.branch\[1\].mux_I/um_ow[309] tt_top1.branch\[1\].mux_I/um_ow[30]
+ tt_top1.branch\[1\].mux_I/um_ow[310] tt_top1.branch\[1\].mux_I/um_ow[311] tt_top1.branch\[1\].mux_I/um_ow[312]
+ tt_top1.branch\[1\].mux_I/um_ow[313] tt_top1.branch\[1\].mux_I/um_ow[314] tt_top1.branch\[1\].mux_I/um_ow[315]
+ tt_top1.branch\[1\].mux_I/um_ow[316] tt_top1.branch\[1\].mux_I/um_ow[317] tt_top1.branch\[1\].mux_I/um_ow[318]
+ tt_top1.branch\[1\].mux_I/um_ow[319] tt_top1.branch\[1\].mux_I/um_ow[31] tt_top1.branch\[1\].mux_I/um_ow[320]
+ tt_top1.branch\[1\].mux_I/um_ow[321] tt_top1.branch\[1\].mux_I/um_ow[322] tt_top1.branch\[1\].mux_I/um_ow[323]
+ tt_top1.branch\[1\].mux_I/um_ow[324] tt_top1.branch\[1\].mux_I/um_ow[325] tt_top1.branch\[1\].mux_I/um_ow[326]
+ tt_top1.branch\[1\].mux_I/um_ow[327] tt_top1.branch\[1\].mux_I/um_ow[328] tt_top1.branch\[1\].mux_I/um_ow[329]
+ tt_top1.branch\[1\].mux_I/um_ow[32] tt_top1.branch\[1\].mux_I/um_ow[330] tt_top1.branch\[1\].mux_I/um_ow[331]
+ tt_top1.branch\[1\].mux_I/um_ow[332] tt_top1.branch\[1\].mux_I/um_ow[333] tt_top1.branch\[1\].mux_I/um_ow[334]
+ tt_top1.branch\[1\].mux_I/um_ow[335] tt_top1.branch\[1\].mux_I/um_ow[336] tt_top1.branch\[1\].mux_I/um_ow[337]
+ tt_top1.branch\[1\].mux_I/um_ow[338] tt_top1.branch\[1\].mux_I/um_ow[339] tt_top1.branch\[1\].mux_I/um_ow[33]
+ tt_top1.branch\[1\].mux_I/um_ow[340] tt_top1.branch\[1\].mux_I/um_ow[341] tt_top1.branch\[1\].mux_I/um_ow[342]
+ tt_top1.branch\[1\].mux_I/um_ow[343] tt_top1.branch\[1\].mux_I/um_ow[344] tt_top1.branch\[1\].mux_I/um_ow[345]
+ tt_top1.branch\[1\].mux_I/um_ow[346] tt_top1.branch\[1\].mux_I/um_ow[347] tt_top1.branch\[1\].mux_I/um_ow[348]
+ tt_top1.branch\[1\].mux_I/um_ow[349] tt_top1.branch\[1\].mux_I/um_ow[34] tt_top1.branch\[1\].mux_I/um_ow[350]
+ tt_top1.branch\[1\].mux_I/um_ow[351] tt_top1.branch\[1\].mux_I/um_ow[352] tt_top1.branch\[1\].mux_I/um_ow[353]
+ tt_top1.branch\[1\].mux_I/um_ow[354] tt_top1.branch\[1\].mux_I/um_ow[355] tt_top1.branch\[1\].mux_I/um_ow[356]
+ tt_top1.branch\[1\].mux_I/um_ow[357] tt_top1.branch\[1\].mux_I/um_ow[358] tt_top1.branch\[1\].mux_I/um_ow[359]
+ tt_top1.branch\[1\].mux_I/um_ow[35] tt_top1.branch\[1\].mux_I/um_ow[360] tt_top1.branch\[1\].mux_I/um_ow[361]
+ tt_top1.branch\[1\].mux_I/um_ow[362] tt_top1.branch\[1\].mux_I/um_ow[363] tt_top1.branch\[1\].mux_I/um_ow[364]
+ tt_top1.branch\[1\].mux_I/um_ow[365] tt_top1.branch\[1\].mux_I/um_ow[366] tt_top1.branch\[1\].mux_I/um_ow[367]
+ tt_top1.branch\[1\].mux_I/um_ow[368] tt_top1.branch\[1\].mux_I/um_ow[369] tt_top1.branch\[1\].mux_I/um_ow[36]
+ tt_top1.branch\[1\].mux_I/um_ow[370] tt_top1.branch\[1\].mux_I/um_ow[371] tt_top1.branch\[1\].mux_I/um_ow[372]
+ tt_top1.branch\[1\].mux_I/um_ow[373] tt_top1.branch\[1\].mux_I/um_ow[374] tt_top1.branch\[1\].mux_I/um_ow[375]
+ tt_top1.branch\[1\].mux_I/um_ow[376] tt_top1.branch\[1\].mux_I/um_ow[377] tt_top1.branch\[1\].mux_I/um_ow[378]
+ tt_top1.branch\[1\].mux_I/um_ow[379] tt_top1.branch\[1\].mux_I/um_ow[37] tt_top1.branch\[1\].mux_I/um_ow[380]
+ tt_top1.branch\[1\].mux_I/um_ow[381] tt_top1.branch\[1\].mux_I/um_ow[382] tt_top1.branch\[1\].mux_I/um_ow[383]
+ tt_top1.branch\[1\].mux_I/um_ow[38] tt_top1.branch\[1\].mux_I/um_ow[39] tt_top1.branch\[1\].mux_I/um_ow[3]
+ tt_top1.branch\[1\].mux_I/um_ow[40] tt_top1.branch\[1\].mux_I/um_ow[41] tt_top1.branch\[1\].mux_I/um_ow[42]
+ tt_top1.branch\[1\].mux_I/um_ow[43] tt_top1.branch\[1\].mux_I/um_ow[44] tt_top1.branch\[1\].mux_I/um_ow[45]
+ tt_top1.branch\[1\].mux_I/um_ow[46] tt_top1.branch\[1\].mux_I/um_ow[47] tt_top1.branch\[1\].mux_I/um_ow[48]
+ tt_top1.branch\[1\].mux_I/um_ow[49] tt_top1.branch\[1\].mux_I/um_ow[4] tt_top1.branch\[1\].mux_I/um_ow[50]
+ tt_top1.branch\[1\].mux_I/um_ow[51] tt_top1.branch\[1\].mux_I/um_ow[52] tt_top1.branch\[1\].mux_I/um_ow[53]
+ tt_top1.branch\[1\].mux_I/um_ow[54] tt_top1.branch\[1\].mux_I/um_ow[55] tt_top1.branch\[1\].mux_I/um_ow[56]
+ tt_top1.branch\[1\].mux_I/um_ow[57] tt_top1.branch\[1\].mux_I/um_ow[58] tt_top1.branch\[1\].mux_I/um_ow[59]
+ tt_top1.branch\[1\].mux_I/um_ow[5] tt_top1.branch\[1\].mux_I/um_ow[60] tt_top1.branch\[1\].mux_I/um_ow[61]
+ tt_top1.branch\[1\].mux_I/um_ow[62] tt_top1.branch\[1\].mux_I/um_ow[63] tt_top1.branch\[1\].mux_I/um_ow[64]
+ tt_top1.branch\[1\].mux_I/um_ow[65] tt_top1.branch\[1\].mux_I/um_ow[66] tt_top1.branch\[1\].mux_I/um_ow[67]
+ tt_top1.branch\[1\].mux_I/um_ow[68] tt_top1.branch\[1\].mux_I/um_ow[69] tt_top1.branch\[1\].mux_I/um_ow[6]
+ tt_top1.branch\[1\].mux_I/um_ow[70] tt_top1.branch\[1\].mux_I/um_ow[71] tt_top1.branch\[1\].mux_I/um_ow[72]
+ tt_top1.branch\[1\].mux_I/um_ow[73] tt_top1.branch\[1\].mux_I/um_ow[74] tt_top1.branch\[1\].mux_I/um_ow[75]
+ tt_top1.branch\[1\].mux_I/um_ow[76] tt_top1.branch\[1\].mux_I/um_ow[77] tt_top1.branch\[1\].mux_I/um_ow[78]
+ tt_top1.branch\[1\].mux_I/um_ow[79] tt_top1.branch\[1\].mux_I/um_ow[7] tt_top1.branch\[1\].mux_I/um_ow[80]
+ tt_top1.branch\[1\].mux_I/um_ow[81] tt_top1.branch\[1\].mux_I/um_ow[82] tt_top1.branch\[1\].mux_I/um_ow[83]
+ tt_top1.branch\[1\].mux_I/um_ow[84] tt_top1.branch\[1\].mux_I/um_ow[85] tt_top1.branch\[1\].mux_I/um_ow[86]
+ tt_top1.branch\[1\].mux_I/um_ow[87] tt_top1.branch\[1\].mux_I/um_ow[88] tt_top1.branch\[1\].mux_I/um_ow[89]
+ tt_top1.branch\[1\].mux_I/um_ow[8] tt_top1.branch\[1\].mux_I/um_ow[90] tt_top1.branch\[1\].mux_I/um_ow[91]
+ tt_top1.branch\[1\].mux_I/um_ow[92] tt_top1.branch\[1\].mux_I/um_ow[93] tt_top1.branch\[1\].mux_I/um_ow[94]
+ tt_top1.branch\[1\].mux_I/um_ow[95] tt_top1.branch\[1\].mux_I/um_ow[96] tt_top1.branch\[1\].mux_I/um_ow[97]
+ tt_top1.branch\[1\].mux_I/um_ow[98] tt_top1.branch\[1\].mux_I/um_ow[99] tt_top1.branch\[1\].mux_I/um_ow[9]
+ vccd1 vssd1 tt_mux
Xtt_top1.branch\[0\].col_um\[1\].um_top_I.block_1_1.tt_um_I tt_top1.branch\[0\].mux_I/um_iw[54]
+ tt_top1.branch\[0\].mux_I/um_ena[3] tt_top1.branch\[0\].mux_I/um_iw[55] tt_top1.branch\[0\].mux_I/um_iw[56]
+ tt_top1.branch\[0\].mux_I/um_iw[57] tt_top1.branch\[0\].mux_I/um_iw[58] tt_top1.branch\[0\].mux_I/um_iw[59]
+ tt_top1.branch\[0\].mux_I/um_iw[60] tt_top1.branch\[0\].mux_I/um_iw[61] tt_top1.branch\[0\].mux_I/um_iw[62]
+ tt_top1.branch\[0\].mux_I/um_iw[63] tt_top1.branch\[0\].mux_I/um_iw[64] tt_top1.branch\[0\].mux_I/um_iw[65]
+ tt_top1.branch\[0\].mux_I/um_iw[66] tt_top1.branch\[0\].mux_I/um_iw[67] tt_top1.branch\[0\].mux_I/um_iw[68]
+ tt_top1.branch\[0\].mux_I/um_iw[69] tt_top1.branch\[0\].mux_I/um_iw[70] tt_top1.branch\[0\].mux_I/um_iw[71]
+ tt_top1.branch\[0\].mux_I/um_ow[88] tt_top1.branch\[0\].mux_I/um_ow[89] tt_top1.branch\[0\].mux_I/um_ow[90]
+ tt_top1.branch\[0\].mux_I/um_ow[91] tt_top1.branch\[0\].mux_I/um_ow[92] tt_top1.branch\[0\].mux_I/um_ow[93]
+ tt_top1.branch\[0\].mux_I/um_ow[94] tt_top1.branch\[0\].mux_I/um_ow[95] tt_top1.branch\[0\].mux_I/um_ow[80]
+ tt_top1.branch\[0\].mux_I/um_ow[81] tt_top1.branch\[0\].mux_I/um_ow[82] tt_top1.branch\[0\].mux_I/um_ow[83]
+ tt_top1.branch\[0\].mux_I/um_ow[84] tt_top1.branch\[0\].mux_I/um_ow[85] tt_top1.branch\[0\].mux_I/um_ow[86]
+ tt_top1.branch\[0\].mux_I/um_ow[87] tt_top1.branch\[0\].mux_I/um_ow[72] tt_top1.branch\[0\].mux_I/um_ow[73]
+ tt_top1.branch\[0\].mux_I/um_ow[74] tt_top1.branch\[0\].mux_I/um_ow[75] tt_top1.branch\[0\].mux_I/um_ow[76]
+ tt_top1.branch\[0\].mux_I/um_ow[77] tt_top1.branch\[0\].mux_I/um_ow[78] tt_top1.branch\[0\].mux_I/um_ow[79]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[1\].col_um\[6\].um_top_I.block_1_22.tt_um_I tt_top1.branch\[1\].mux_I/um_iw[234]
+ tt_top1.branch\[1\].mux_I/um_ena[13] tt_top1.branch\[1\].mux_I/um_iw[235] tt_top1.branch\[1\].mux_I/um_iw[236]
+ tt_top1.branch\[1\].mux_I/um_iw[237] tt_top1.branch\[1\].mux_I/um_iw[238] tt_top1.branch\[1\].mux_I/um_iw[239]
+ tt_top1.branch\[1\].mux_I/um_iw[240] tt_top1.branch\[1\].mux_I/um_iw[241] tt_top1.branch\[1\].mux_I/um_iw[242]
+ tt_top1.branch\[1\].mux_I/um_iw[243] tt_top1.branch\[1\].mux_I/um_iw[244] tt_top1.branch\[1\].mux_I/um_iw[245]
+ tt_top1.branch\[1\].mux_I/um_iw[246] tt_top1.branch\[1\].mux_I/um_iw[247] tt_top1.branch\[1\].mux_I/um_iw[248]
+ tt_top1.branch\[1\].mux_I/um_iw[249] tt_top1.branch\[1\].mux_I/um_iw[250] tt_top1.branch\[1\].mux_I/um_iw[251]
+ tt_top1.branch\[1\].mux_I/um_ow[328] tt_top1.branch\[1\].mux_I/um_ow[329] tt_top1.branch\[1\].mux_I/um_ow[330]
+ tt_top1.branch\[1\].mux_I/um_ow[331] tt_top1.branch\[1\].mux_I/um_ow[332] tt_top1.branch\[1\].mux_I/um_ow[333]
+ tt_top1.branch\[1\].mux_I/um_ow[334] tt_top1.branch\[1\].mux_I/um_ow[335] tt_top1.branch\[1\].mux_I/um_ow[320]
+ tt_top1.branch\[1\].mux_I/um_ow[321] tt_top1.branch\[1\].mux_I/um_ow[322] tt_top1.branch\[1\].mux_I/um_ow[323]
+ tt_top1.branch\[1\].mux_I/um_ow[324] tt_top1.branch\[1\].mux_I/um_ow[325] tt_top1.branch\[1\].mux_I/um_ow[326]
+ tt_top1.branch\[1\].mux_I/um_ow[327] tt_top1.branch\[1\].mux_I/um_ow[312] tt_top1.branch\[1\].mux_I/um_ow[313]
+ tt_top1.branch\[1\].mux_I/um_ow[314] tt_top1.branch\[1\].mux_I/um_ow[315] tt_top1.branch\[1\].mux_I/um_ow[316]
+ tt_top1.branch\[1\].mux_I/um_ow[317] tt_top1.branch\[1\].mux_I/um_ow[318] tt_top1.branch\[1\].mux_I/um_ow[319]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[1\].col_um\[7\].um_bot_I.block_0_23.tt_um_I tt_top1.branch\[1\].mux_I/um_iw[252]
+ tt_top1.branch\[1\].mux_I/um_ena[14] tt_top1.branch\[1\].mux_I/um_iw[253] tt_top1.branch\[1\].mux_I/um_iw[254]
+ tt_top1.branch\[1\].mux_I/um_iw[255] tt_top1.branch\[1\].mux_I/um_iw[256] tt_top1.branch\[1\].mux_I/um_iw[257]
+ tt_top1.branch\[1\].mux_I/um_iw[258] tt_top1.branch\[1\].mux_I/um_iw[259] tt_top1.branch\[1\].mux_I/um_iw[260]
+ tt_top1.branch\[1\].mux_I/um_iw[261] tt_top1.branch\[1\].mux_I/um_iw[262] tt_top1.branch\[1\].mux_I/um_iw[263]
+ tt_top1.branch\[1\].mux_I/um_iw[264] tt_top1.branch\[1\].mux_I/um_iw[265] tt_top1.branch\[1\].mux_I/um_iw[266]
+ tt_top1.branch\[1\].mux_I/um_iw[267] tt_top1.branch\[1\].mux_I/um_iw[268] tt_top1.branch\[1\].mux_I/um_iw[269]
+ tt_top1.branch\[1\].mux_I/um_ow[352] tt_top1.branch\[1\].mux_I/um_ow[353] tt_top1.branch\[1\].mux_I/um_ow[354]
+ tt_top1.branch\[1\].mux_I/um_ow[355] tt_top1.branch\[1\].mux_I/um_ow[356] tt_top1.branch\[1\].mux_I/um_ow[357]
+ tt_top1.branch\[1\].mux_I/um_ow[358] tt_top1.branch\[1\].mux_I/um_ow[359] tt_top1.branch\[1\].mux_I/um_ow[344]
+ tt_top1.branch\[1\].mux_I/um_ow[345] tt_top1.branch\[1\].mux_I/um_ow[346] tt_top1.branch\[1\].mux_I/um_ow[347]
+ tt_top1.branch\[1\].mux_I/um_ow[348] tt_top1.branch\[1\].mux_I/um_ow[349] tt_top1.branch\[1\].mux_I/um_ow[350]
+ tt_top1.branch\[1\].mux_I/um_ow[351] tt_top1.branch\[1\].mux_I/um_ow[336] tt_top1.branch\[1\].mux_I/um_ow[337]
+ tt_top1.branch\[1\].mux_I/um_ow[338] tt_top1.branch\[1\].mux_I/um_ow[339] tt_top1.branch\[1\].mux_I/um_ow[340]
+ tt_top1.branch\[1\].mux_I/um_ow[341] tt_top1.branch\[1\].mux_I/um_ow[342] tt_top1.branch\[1\].mux_I/um_ow[343]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[1\].col_um\[0\].um_top_I.block_1_16.tt_um_I tt_top1.branch\[1\].mux_I/um_iw[18]
+ tt_top1.branch\[1\].mux_I/um_ena[1] tt_top1.branch\[1\].mux_I/um_iw[19] tt_top1.branch\[1\].mux_I/um_iw[20]
+ tt_top1.branch\[1\].mux_I/um_iw[21] tt_top1.branch\[1\].mux_I/um_iw[22] tt_top1.branch\[1\].mux_I/um_iw[23]
+ tt_top1.branch\[1\].mux_I/um_iw[24] tt_top1.branch\[1\].mux_I/um_iw[25] tt_top1.branch\[1\].mux_I/um_iw[26]
+ tt_top1.branch\[1\].mux_I/um_iw[27] tt_top1.branch\[1\].mux_I/um_iw[28] tt_top1.branch\[1\].mux_I/um_iw[29]
+ tt_top1.branch\[1\].mux_I/um_iw[30] tt_top1.branch\[1\].mux_I/um_iw[31] tt_top1.branch\[1\].mux_I/um_iw[32]
+ tt_top1.branch\[1\].mux_I/um_iw[33] tt_top1.branch\[1\].mux_I/um_iw[34] tt_top1.branch\[1\].mux_I/um_iw[35]
+ tt_top1.branch\[1\].mux_I/um_ow[40] tt_top1.branch\[1\].mux_I/um_ow[41] tt_top1.branch\[1\].mux_I/um_ow[42]
+ tt_top1.branch\[1\].mux_I/um_ow[43] tt_top1.branch\[1\].mux_I/um_ow[44] tt_top1.branch\[1\].mux_I/um_ow[45]
+ tt_top1.branch\[1\].mux_I/um_ow[46] tt_top1.branch\[1\].mux_I/um_ow[47] tt_top1.branch\[1\].mux_I/um_ow[32]
+ tt_top1.branch\[1\].mux_I/um_ow[33] tt_top1.branch\[1\].mux_I/um_ow[34] tt_top1.branch\[1\].mux_I/um_ow[35]
+ tt_top1.branch\[1\].mux_I/um_ow[36] tt_top1.branch\[1\].mux_I/um_ow[37] tt_top1.branch\[1\].mux_I/um_ow[38]
+ tt_top1.branch\[1\].mux_I/um_ow[39] tt_top1.branch\[1\].mux_I/um_ow[24] tt_top1.branch\[1\].mux_I/um_ow[25]
+ tt_top1.branch\[1\].mux_I/um_ow[26] tt_top1.branch\[1\].mux_I/um_ow[27] tt_top1.branch\[1\].mux_I/um_ow[28]
+ tt_top1.branch\[1\].mux_I/um_ow[29] tt_top1.branch\[1\].mux_I/um_ow[30] tt_top1.branch\[1\].mux_I/um_ow[31]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[0\].col_um\[0\].um_top_I.block_1_0.tt_um_I tt_top1.branch\[0\].mux_I/um_iw[18]
+ tt_top1.branch\[0\].mux_I/um_ena[1] tt_top1.branch\[0\].mux_I/um_iw[19] tt_top1.branch\[0\].mux_I/um_iw[20]
+ tt_top1.branch\[0\].mux_I/um_iw[21] tt_top1.branch\[0\].mux_I/um_iw[22] tt_top1.branch\[0\].mux_I/um_iw[23]
+ tt_top1.branch\[0\].mux_I/um_iw[24] tt_top1.branch\[0\].mux_I/um_iw[25] tt_top1.branch\[0\].mux_I/um_iw[26]
+ tt_top1.branch\[0\].mux_I/um_iw[27] tt_top1.branch\[0\].mux_I/um_iw[28] tt_top1.branch\[0\].mux_I/um_iw[29]
+ tt_top1.branch\[0\].mux_I/um_iw[30] tt_top1.branch\[0\].mux_I/um_iw[31] tt_top1.branch\[0\].mux_I/um_iw[32]
+ tt_top1.branch\[0\].mux_I/um_iw[33] tt_top1.branch\[0\].mux_I/um_iw[34] tt_top1.branch\[0\].mux_I/um_iw[35]
+ tt_top1.branch\[0\].mux_I/um_ow[40] tt_top1.branch\[0\].mux_I/um_ow[41] tt_top1.branch\[0\].mux_I/um_ow[42]
+ tt_top1.branch\[0\].mux_I/um_ow[43] tt_top1.branch\[0\].mux_I/um_ow[44] tt_top1.branch\[0\].mux_I/um_ow[45]
+ tt_top1.branch\[0\].mux_I/um_ow[46] tt_top1.branch\[0\].mux_I/um_ow[47] tt_top1.branch\[0\].mux_I/um_ow[32]
+ tt_top1.branch\[0\].mux_I/um_ow[33] tt_top1.branch\[0\].mux_I/um_ow[34] tt_top1.branch\[0\].mux_I/um_ow[35]
+ tt_top1.branch\[0\].mux_I/um_ow[36] tt_top1.branch\[0\].mux_I/um_ow[37] tt_top1.branch\[0\].mux_I/um_ow[38]
+ tt_top1.branch\[0\].mux_I/um_ow[39] tt_top1.branch\[0\].mux_I/um_ow[24] tt_top1.branch\[0\].mux_I/um_ow[25]
+ tt_top1.branch\[0\].mux_I/um_ow[26] tt_top1.branch\[0\].mux_I/um_ow[27] tt_top1.branch\[0\].mux_I/um_ow[28]
+ tt_top1.branch\[0\].mux_I/um_ow[29] tt_top1.branch\[0\].mux_I/um_ow[30] tt_top1.branch\[0\].mux_I/um_ow[31]
+ vccd1 vssd1 tt_um_test
Xtt_top1.ctrl_I io_in[32] io_in[34] io_in[36] io_out[9] io_out[4] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[24]
+ io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[30] io_in[31] io_oeb[24]
+ io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[30] io_oeb[31] io_out[24]
+ io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[30] io_out[31] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[20] io_out[21] io_out[22] io_out[23] tt_top1.ctrl_I/spine_iw[0]
+ tt_top1.ctrl_I/spine_iw[10] tt_top1.ctrl_I/spine_iw[11] tt_top1.ctrl_I/spine_iw[12]
+ tt_top1.ctrl_I/spine_iw[13] tt_top1.ctrl_I/spine_iw[14] tt_top1.ctrl_I/spine_iw[15]
+ tt_top1.ctrl_I/spine_iw[16] tt_top1.ctrl_I/spine_iw[17] tt_top1.ctrl_I/spine_iw[18]
+ tt_top1.ctrl_I/spine_iw[19] tt_top1.ctrl_I/spine_iw[1] tt_top1.ctrl_I/spine_iw[20]
+ tt_top1.ctrl_I/spine_iw[21] tt_top1.ctrl_I/spine_iw[22] tt_top1.ctrl_I/spine_iw[23]
+ tt_top1.ctrl_I/spine_iw[24] tt_top1.ctrl_I/spine_iw[25] tt_top1.ctrl_I/spine_iw[26]
+ tt_top1.ctrl_I/spine_iw[27] tt_top1.ctrl_I/spine_iw[28] tt_top1.ctrl_I/spine_iw[29]
+ tt_top1.ctrl_I/spine_iw[2] tt_top1.ctrl_I/spine_iw[30] tt_top1.ctrl_I/spine_iw[3]
+ tt_top1.ctrl_I/spine_iw[4] tt_top1.ctrl_I/spine_iw[5] tt_top1.ctrl_I/spine_iw[6]
+ tt_top1.ctrl_I/spine_iw[7] tt_top1.ctrl_I/spine_iw[8] tt_top1.ctrl_I/spine_iw[9]
+ tt_top1.ctrl_I/spine_ow[0] tt_top1.ctrl_I/spine_ow[10] tt_top1.ctrl_I/spine_ow[11]
+ tt_top1.ctrl_I/spine_ow[12] tt_top1.ctrl_I/spine_ow[13] tt_top1.ctrl_I/spine_ow[14]
+ tt_top1.ctrl_I/spine_ow[15] tt_top1.ctrl_I/spine_ow[16] tt_top1.ctrl_I/spine_ow[17]
+ tt_top1.ctrl_I/spine_ow[18] tt_top1.ctrl_I/spine_ow[19] tt_top1.ctrl_I/spine_ow[1]
+ tt_top1.ctrl_I/spine_ow[20] tt_top1.ctrl_I/spine_ow[21] tt_top1.ctrl_I/spine_ow[22]
+ tt_top1.ctrl_I/spine_ow[23] tt_top1.ctrl_I/spine_ow[24] tt_top1.ctrl_I/spine_ow[25]
+ tt_top1.ctrl_I/spine_ow[2] tt_top1.ctrl_I/spine_ow[3] tt_top1.ctrl_I/spine_ow[4]
+ tt_top1.ctrl_I/spine_ow[5] tt_top1.ctrl_I/spine_ow[6] tt_top1.ctrl_I/spine_ow[7]
+ tt_top1.ctrl_I/spine_ow[8] tt_top1.ctrl_I/spine_ow[9] vccd1 vssd1 tt_ctrl
Xtt_top1.branch\[1\].col_um\[1\].um_bot_I.block_0_17.tt_um_I tt_top1.branch\[1\].mux_I/um_iw[36]
+ tt_top1.branch\[1\].mux_I/um_ena[2] tt_top1.branch\[1\].mux_I/um_iw[37] tt_top1.branch\[1\].mux_I/um_iw[38]
+ tt_top1.branch\[1\].mux_I/um_iw[39] tt_top1.branch\[1\].mux_I/um_iw[40] tt_top1.branch\[1\].mux_I/um_iw[41]
+ tt_top1.branch\[1\].mux_I/um_iw[42] tt_top1.branch\[1\].mux_I/um_iw[43] tt_top1.branch\[1\].mux_I/um_iw[44]
+ tt_top1.branch\[1\].mux_I/um_iw[45] tt_top1.branch\[1\].mux_I/um_iw[46] tt_top1.branch\[1\].mux_I/um_iw[47]
+ tt_top1.branch\[1\].mux_I/um_iw[48] tt_top1.branch\[1\].mux_I/um_iw[49] tt_top1.branch\[1\].mux_I/um_iw[50]
+ tt_top1.branch\[1\].mux_I/um_iw[51] tt_top1.branch\[1\].mux_I/um_iw[52] tt_top1.branch\[1\].mux_I/um_iw[53]
+ tt_top1.branch\[1\].mux_I/um_ow[64] tt_top1.branch\[1\].mux_I/um_ow[65] tt_top1.branch\[1\].mux_I/um_ow[66]
+ tt_top1.branch\[1\].mux_I/um_ow[67] tt_top1.branch\[1\].mux_I/um_ow[68] tt_top1.branch\[1\].mux_I/um_ow[69]
+ tt_top1.branch\[1\].mux_I/um_ow[70] tt_top1.branch\[1\].mux_I/um_ow[71] tt_top1.branch\[1\].mux_I/um_ow[56]
+ tt_top1.branch\[1\].mux_I/um_ow[57] tt_top1.branch\[1\].mux_I/um_ow[58] tt_top1.branch\[1\].mux_I/um_ow[59]
+ tt_top1.branch\[1\].mux_I/um_ow[60] tt_top1.branch\[1\].mux_I/um_ow[61] tt_top1.branch\[1\].mux_I/um_ow[62]
+ tt_top1.branch\[1\].mux_I/um_ow[63] tt_top1.branch\[1\].mux_I/um_ow[48] tt_top1.branch\[1\].mux_I/um_ow[49]
+ tt_top1.branch\[1\].mux_I/um_ow[50] tt_top1.branch\[1\].mux_I/um_ow[51] tt_top1.branch\[1\].mux_I/um_ow[52]
+ tt_top1.branch\[1\].mux_I/um_ow[53] tt_top1.branch\[1\].mux_I/um_ow[54] tt_top1.branch\[1\].mux_I/um_ow[55]
+ vccd1 vssd1 tt_um_moyes0_top_module
Xtt_top1.branch\[1\].col_um\[4\].um_bot_I.block_0_20.tt_um_I tt_top1.branch\[1\].mux_I/um_iw[144]
+ tt_top1.branch\[1\].mux_I/um_ena[8] tt_top1.branch\[1\].mux_I/um_iw[145] tt_top1.branch\[1\].mux_I/um_iw[146]
+ tt_top1.branch\[1\].mux_I/um_iw[147] tt_top1.branch\[1\].mux_I/um_iw[148] tt_top1.branch\[1\].mux_I/um_iw[149]
+ tt_top1.branch\[1\].mux_I/um_iw[150] tt_top1.branch\[1\].mux_I/um_iw[151] tt_top1.branch\[1\].mux_I/um_iw[152]
+ tt_top1.branch\[1\].mux_I/um_iw[153] tt_top1.branch\[1\].mux_I/um_iw[154] tt_top1.branch\[1\].mux_I/um_iw[155]
+ tt_top1.branch\[1\].mux_I/um_iw[156] tt_top1.branch\[1\].mux_I/um_iw[157] tt_top1.branch\[1\].mux_I/um_iw[158]
+ tt_top1.branch\[1\].mux_I/um_iw[159] tt_top1.branch\[1\].mux_I/um_iw[160] tt_top1.branch\[1\].mux_I/um_iw[161]
+ tt_top1.branch\[1\].mux_I/um_ow[208] tt_top1.branch\[1\].mux_I/um_ow[209] tt_top1.branch\[1\].mux_I/um_ow[210]
+ tt_top1.branch\[1\].mux_I/um_ow[211] tt_top1.branch\[1\].mux_I/um_ow[212] tt_top1.branch\[1\].mux_I/um_ow[213]
+ tt_top1.branch\[1\].mux_I/um_ow[214] tt_top1.branch\[1\].mux_I/um_ow[215] tt_top1.branch\[1\].mux_I/um_ow[200]
+ tt_top1.branch\[1\].mux_I/um_ow[201] tt_top1.branch\[1\].mux_I/um_ow[202] tt_top1.branch\[1\].mux_I/um_ow[203]
+ tt_top1.branch\[1\].mux_I/um_ow[204] tt_top1.branch\[1\].mux_I/um_ow[205] tt_top1.branch\[1\].mux_I/um_ow[206]
+ tt_top1.branch\[1\].mux_I/um_ow[207] tt_top1.branch\[1\].mux_I/um_ow[192] tt_top1.branch\[1\].mux_I/um_ow[193]
+ tt_top1.branch\[1\].mux_I/um_ow[194] tt_top1.branch\[1\].mux_I/um_ow[195] tt_top1.branch\[1\].mux_I/um_ow[196]
+ tt_top1.branch\[1\].mux_I/um_ow[197] tt_top1.branch\[1\].mux_I/um_ow[198] tt_top1.branch\[1\].mux_I/um_ow[199]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[0\].mux_I tt_top1.branch\[0\].mux_I/k_zero tt_top1.branch\[0\].mux_I/k_zero
+ tt_top1.branch\[0\].mux_I/k_zero tt_top1.branch\[0\].mux_I/k_zero tt_top1.branch\[0\].mux_I/k_zero
+ tt_top1.branch\[0\].mux_I/k_one tt_top1.branch\[0\].mux_I/k_zero tt_top1.ctrl_I/spine_iw[0]
+ tt_top1.ctrl_I/spine_iw[10] tt_top1.ctrl_I/spine_iw[11] tt_top1.ctrl_I/spine_iw[12]
+ tt_top1.ctrl_I/spine_iw[13] tt_top1.ctrl_I/spine_iw[14] tt_top1.ctrl_I/spine_iw[15]
+ tt_top1.ctrl_I/spine_iw[16] tt_top1.ctrl_I/spine_iw[17] tt_top1.ctrl_I/spine_iw[18]
+ tt_top1.ctrl_I/spine_iw[19] tt_top1.ctrl_I/spine_iw[1] tt_top1.ctrl_I/spine_iw[20]
+ tt_top1.ctrl_I/spine_iw[21] tt_top1.ctrl_I/spine_iw[22] tt_top1.ctrl_I/spine_iw[23]
+ tt_top1.ctrl_I/spine_iw[24] tt_top1.ctrl_I/spine_iw[25] tt_top1.ctrl_I/spine_iw[26]
+ tt_top1.ctrl_I/spine_iw[27] tt_top1.ctrl_I/spine_iw[28] tt_top1.ctrl_I/spine_iw[29]
+ tt_top1.ctrl_I/spine_iw[2] tt_top1.ctrl_I/spine_iw[30] tt_top1.ctrl_I/spine_iw[3]
+ tt_top1.ctrl_I/spine_iw[4] tt_top1.ctrl_I/spine_iw[5] tt_top1.ctrl_I/spine_iw[6]
+ tt_top1.ctrl_I/spine_iw[7] tt_top1.ctrl_I/spine_iw[8] tt_top1.ctrl_I/spine_iw[9]
+ tt_top1.ctrl_I/spine_ow[0] tt_top1.ctrl_I/spine_ow[10] tt_top1.ctrl_I/spine_ow[11]
+ tt_top1.ctrl_I/spine_ow[12] tt_top1.ctrl_I/spine_ow[13] tt_top1.ctrl_I/spine_ow[14]
+ tt_top1.ctrl_I/spine_ow[15] tt_top1.ctrl_I/spine_ow[16] tt_top1.ctrl_I/spine_ow[17]
+ tt_top1.ctrl_I/spine_ow[18] tt_top1.ctrl_I/spine_ow[19] tt_top1.ctrl_I/spine_ow[1]
+ tt_top1.ctrl_I/spine_ow[20] tt_top1.ctrl_I/spine_ow[21] tt_top1.ctrl_I/spine_ow[22]
+ tt_top1.ctrl_I/spine_ow[23] tt_top1.ctrl_I/spine_ow[24] tt_top1.ctrl_I/spine_ow[25]
+ tt_top1.ctrl_I/spine_ow[2] tt_top1.ctrl_I/spine_ow[3] tt_top1.ctrl_I/spine_ow[4]
+ tt_top1.ctrl_I/spine_ow[5] tt_top1.ctrl_I/spine_ow[6] tt_top1.ctrl_I/spine_ow[7]
+ tt_top1.ctrl_I/spine_ow[8] tt_top1.ctrl_I/spine_ow[9] tt_top1.branch\[0\].mux_I/um_ena[0]
+ tt_top1.branch\[0\].mux_I/um_ena[10] tt_top1.branch\[0\].mux_I/um_ena[11] tt_top1.branch\[0\].mux_I/um_ena[12]
+ tt_top1.branch\[0\].mux_I/um_ena[13] tt_top1.branch\[0\].mux_I/um_ena[14] tt_top1.branch\[0\].mux_I/um_ena[15]
+ tt_top1.branch\[0\].mux_I/um_ena[1] tt_top1.branch\[0\].mux_I/um_ena[2] tt_top1.branch\[0\].mux_I/um_ena[3]
+ tt_top1.branch\[0\].mux_I/um_ena[4] tt_top1.branch\[0\].mux_I/um_ena[5] tt_top1.branch\[0\].mux_I/um_ena[6]
+ tt_top1.branch\[0\].mux_I/um_ena[7] tt_top1.branch\[0\].mux_I/um_ena[8] tt_top1.branch\[0\].mux_I/um_ena[9]
+ tt_top1.branch\[0\].mux_I/um_iw[0] tt_top1.branch\[0\].mux_I/um_iw[100] tt_top1.branch\[0\].mux_I/um_iw[101]
+ tt_top1.branch\[0\].mux_I/um_iw[102] tt_top1.branch\[0\].mux_I/um_iw[103] tt_top1.branch\[0\].mux_I/um_iw[104]
+ tt_top1.branch\[0\].mux_I/um_iw[105] tt_top1.branch\[0\].mux_I/um_iw[106] tt_top1.branch\[0\].mux_I/um_iw[107]
+ tt_top1.branch\[0\].mux_I/um_iw[108] tt_top1.branch\[0\].mux_I/um_iw[109] tt_top1.branch\[0\].mux_I/um_iw[10]
+ tt_top1.branch\[0\].mux_I/um_iw[110] tt_top1.branch\[0\].mux_I/um_iw[111] tt_top1.branch\[0\].mux_I/um_iw[112]
+ tt_top1.branch\[0\].mux_I/um_iw[113] tt_top1.branch\[0\].mux_I/um_iw[114] tt_top1.branch\[0\].mux_I/um_iw[115]
+ tt_top1.branch\[0\].mux_I/um_iw[116] tt_top1.branch\[0\].mux_I/um_iw[117] tt_top1.branch\[0\].mux_I/um_iw[118]
+ tt_top1.branch\[0\].mux_I/um_iw[119] tt_top1.branch\[0\].mux_I/um_iw[11] tt_top1.branch\[0\].mux_I/um_iw[120]
+ tt_top1.branch\[0\].mux_I/um_iw[121] tt_top1.branch\[0\].mux_I/um_iw[122] tt_top1.branch\[0\].mux_I/um_iw[123]
+ tt_top1.branch\[0\].mux_I/um_iw[124] tt_top1.branch\[0\].mux_I/um_iw[125] tt_top1.branch\[0\].mux_I/um_iw[126]
+ tt_top1.branch\[0\].mux_I/um_iw[127] tt_top1.branch\[0\].mux_I/um_iw[128] tt_top1.branch\[0\].mux_I/um_iw[129]
+ tt_top1.branch\[0\].mux_I/um_iw[12] tt_top1.branch\[0\].mux_I/um_iw[130] tt_top1.branch\[0\].mux_I/um_iw[131]
+ tt_top1.branch\[0\].mux_I/um_iw[132] tt_top1.branch\[0\].mux_I/um_iw[133] tt_top1.branch\[0\].mux_I/um_iw[134]
+ tt_top1.branch\[0\].mux_I/um_iw[135] tt_top1.branch\[0\].mux_I/um_iw[136] tt_top1.branch\[0\].mux_I/um_iw[137]
+ tt_top1.branch\[0\].mux_I/um_iw[138] tt_top1.branch\[0\].mux_I/um_iw[139] tt_top1.branch\[0\].mux_I/um_iw[13]
+ tt_top1.branch\[0\].mux_I/um_iw[140] tt_top1.branch\[0\].mux_I/um_iw[141] tt_top1.branch\[0\].mux_I/um_iw[142]
+ tt_top1.branch\[0\].mux_I/um_iw[143] tt_top1.branch\[0\].mux_I/um_iw[144] tt_top1.branch\[0\].mux_I/um_iw[145]
+ tt_top1.branch\[0\].mux_I/um_iw[146] tt_top1.branch\[0\].mux_I/um_iw[147] tt_top1.branch\[0\].mux_I/um_iw[148]
+ tt_top1.branch\[0\].mux_I/um_iw[149] tt_top1.branch\[0\].mux_I/um_iw[14] tt_top1.branch\[0\].mux_I/um_iw[150]
+ tt_top1.branch\[0\].mux_I/um_iw[151] tt_top1.branch\[0\].mux_I/um_iw[152] tt_top1.branch\[0\].mux_I/um_iw[153]
+ tt_top1.branch\[0\].mux_I/um_iw[154] tt_top1.branch\[0\].mux_I/um_iw[155] tt_top1.branch\[0\].mux_I/um_iw[156]
+ tt_top1.branch\[0\].mux_I/um_iw[157] tt_top1.branch\[0\].mux_I/um_iw[158] tt_top1.branch\[0\].mux_I/um_iw[159]
+ tt_top1.branch\[0\].mux_I/um_iw[15] tt_top1.branch\[0\].mux_I/um_iw[160] tt_top1.branch\[0\].mux_I/um_iw[161]
+ tt_top1.branch\[0\].mux_I/um_iw[162] tt_top1.branch\[0\].mux_I/um_iw[163] tt_top1.branch\[0\].mux_I/um_iw[164]
+ tt_top1.branch\[0\].mux_I/um_iw[165] tt_top1.branch\[0\].mux_I/um_iw[166] tt_top1.branch\[0\].mux_I/um_iw[167]
+ tt_top1.branch\[0\].mux_I/um_iw[168] tt_top1.branch\[0\].mux_I/um_iw[169] tt_top1.branch\[0\].mux_I/um_iw[16]
+ tt_top1.branch\[0\].mux_I/um_iw[170] tt_top1.branch\[0\].mux_I/um_iw[171] tt_top1.branch\[0\].mux_I/um_iw[172]
+ tt_top1.branch\[0\].mux_I/um_iw[173] tt_top1.branch\[0\].mux_I/um_iw[174] tt_top1.branch\[0\].mux_I/um_iw[175]
+ tt_top1.branch\[0\].mux_I/um_iw[176] tt_top1.branch\[0\].mux_I/um_iw[177] tt_top1.branch\[0\].mux_I/um_iw[178]
+ tt_top1.branch\[0\].mux_I/um_iw[179] tt_top1.branch\[0\].mux_I/um_iw[17] tt_top1.branch\[0\].mux_I/um_iw[180]
+ tt_top1.branch\[0\].mux_I/um_iw[181] tt_top1.branch\[0\].mux_I/um_iw[182] tt_top1.branch\[0\].mux_I/um_iw[183]
+ tt_top1.branch\[0\].mux_I/um_iw[184] tt_top1.branch\[0\].mux_I/um_iw[185] tt_top1.branch\[0\].mux_I/um_iw[186]
+ tt_top1.branch\[0\].mux_I/um_iw[187] tt_top1.branch\[0\].mux_I/um_iw[188] tt_top1.branch\[0\].mux_I/um_iw[189]
+ tt_top1.branch\[0\].mux_I/um_iw[18] tt_top1.branch\[0\].mux_I/um_iw[190] tt_top1.branch\[0\].mux_I/um_iw[191]
+ tt_top1.branch\[0\].mux_I/um_iw[192] tt_top1.branch\[0\].mux_I/um_iw[193] tt_top1.branch\[0\].mux_I/um_iw[194]
+ tt_top1.branch\[0\].mux_I/um_iw[195] tt_top1.branch\[0\].mux_I/um_iw[196] tt_top1.branch\[0\].mux_I/um_iw[197]
+ tt_top1.branch\[0\].mux_I/um_iw[198] tt_top1.branch\[0\].mux_I/um_iw[199] tt_top1.branch\[0\].mux_I/um_iw[19]
+ tt_top1.branch\[0\].mux_I/um_iw[1] tt_top1.branch\[0\].mux_I/um_iw[200] tt_top1.branch\[0\].mux_I/um_iw[201]
+ tt_top1.branch\[0\].mux_I/um_iw[202] tt_top1.branch\[0\].mux_I/um_iw[203] tt_top1.branch\[0\].mux_I/um_iw[204]
+ tt_top1.branch\[0\].mux_I/um_iw[205] tt_top1.branch\[0\].mux_I/um_iw[206] tt_top1.branch\[0\].mux_I/um_iw[207]
+ tt_top1.branch\[0\].mux_I/um_iw[208] tt_top1.branch\[0\].mux_I/um_iw[209] tt_top1.branch\[0\].mux_I/um_iw[20]
+ tt_top1.branch\[0\].mux_I/um_iw[210] tt_top1.branch\[0\].mux_I/um_iw[211] tt_top1.branch\[0\].mux_I/um_iw[212]
+ tt_top1.branch\[0\].mux_I/um_iw[213] tt_top1.branch\[0\].mux_I/um_iw[214] tt_top1.branch\[0\].mux_I/um_iw[215]
+ tt_top1.branch\[0\].mux_I/um_iw[216] tt_top1.branch\[0\].mux_I/um_iw[217] tt_top1.branch\[0\].mux_I/um_iw[218]
+ tt_top1.branch\[0\].mux_I/um_iw[219] tt_top1.branch\[0\].mux_I/um_iw[21] tt_top1.branch\[0\].mux_I/um_iw[220]
+ tt_top1.branch\[0\].mux_I/um_iw[221] tt_top1.branch\[0\].mux_I/um_iw[222] tt_top1.branch\[0\].mux_I/um_iw[223]
+ tt_top1.branch\[0\].mux_I/um_iw[224] tt_top1.branch\[0\].mux_I/um_iw[225] tt_top1.branch\[0\].mux_I/um_iw[226]
+ tt_top1.branch\[0\].mux_I/um_iw[227] tt_top1.branch\[0\].mux_I/um_iw[228] tt_top1.branch\[0\].mux_I/um_iw[229]
+ tt_top1.branch\[0\].mux_I/um_iw[22] tt_top1.branch\[0\].mux_I/um_iw[230] tt_top1.branch\[0\].mux_I/um_iw[231]
+ tt_top1.branch\[0\].mux_I/um_iw[232] tt_top1.branch\[0\].mux_I/um_iw[233] tt_top1.branch\[0\].mux_I/um_iw[234]
+ tt_top1.branch\[0\].mux_I/um_iw[235] tt_top1.branch\[0\].mux_I/um_iw[236] tt_top1.branch\[0\].mux_I/um_iw[237]
+ tt_top1.branch\[0\].mux_I/um_iw[238] tt_top1.branch\[0\].mux_I/um_iw[239] tt_top1.branch\[0\].mux_I/um_iw[23]
+ tt_top1.branch\[0\].mux_I/um_iw[240] tt_top1.branch\[0\].mux_I/um_iw[241] tt_top1.branch\[0\].mux_I/um_iw[242]
+ tt_top1.branch\[0\].mux_I/um_iw[243] tt_top1.branch\[0\].mux_I/um_iw[244] tt_top1.branch\[0\].mux_I/um_iw[245]
+ tt_top1.branch\[0\].mux_I/um_iw[246] tt_top1.branch\[0\].mux_I/um_iw[247] tt_top1.branch\[0\].mux_I/um_iw[248]
+ tt_top1.branch\[0\].mux_I/um_iw[249] tt_top1.branch\[0\].mux_I/um_iw[24] tt_top1.branch\[0\].mux_I/um_iw[250]
+ tt_top1.branch\[0\].mux_I/um_iw[251] tt_top1.branch\[0\].mux_I/um_iw[252] tt_top1.branch\[0\].mux_I/um_iw[253]
+ tt_top1.branch\[0\].mux_I/um_iw[254] tt_top1.branch\[0\].mux_I/um_iw[255] tt_top1.branch\[0\].mux_I/um_iw[256]
+ tt_top1.branch\[0\].mux_I/um_iw[257] tt_top1.branch\[0\].mux_I/um_iw[258] tt_top1.branch\[0\].mux_I/um_iw[259]
+ tt_top1.branch\[0\].mux_I/um_iw[25] tt_top1.branch\[0\].mux_I/um_iw[260] tt_top1.branch\[0\].mux_I/um_iw[261]
+ tt_top1.branch\[0\].mux_I/um_iw[262] tt_top1.branch\[0\].mux_I/um_iw[263] tt_top1.branch\[0\].mux_I/um_iw[264]
+ tt_top1.branch\[0\].mux_I/um_iw[265] tt_top1.branch\[0\].mux_I/um_iw[266] tt_top1.branch\[0\].mux_I/um_iw[267]
+ tt_top1.branch\[0\].mux_I/um_iw[268] tt_top1.branch\[0\].mux_I/um_iw[269] tt_top1.branch\[0\].mux_I/um_iw[26]
+ tt_top1.branch\[0\].mux_I/um_iw[270] tt_top1.branch\[0\].mux_I/um_iw[271] tt_top1.branch\[0\].mux_I/um_iw[272]
+ tt_top1.branch\[0\].mux_I/um_iw[273] tt_top1.branch\[0\].mux_I/um_iw[274] tt_top1.branch\[0\].mux_I/um_iw[275]
+ tt_top1.branch\[0\].mux_I/um_iw[276] tt_top1.branch\[0\].mux_I/um_iw[277] tt_top1.branch\[0\].mux_I/um_iw[278]
+ tt_top1.branch\[0\].mux_I/um_iw[279] tt_top1.branch\[0\].mux_I/um_iw[27] tt_top1.branch\[0\].mux_I/um_iw[280]
+ tt_top1.branch\[0\].mux_I/um_iw[281] tt_top1.branch\[0\].mux_I/um_iw[282] tt_top1.branch\[0\].mux_I/um_iw[283]
+ tt_top1.branch\[0\].mux_I/um_iw[284] tt_top1.branch\[0\].mux_I/um_iw[285] tt_top1.branch\[0\].mux_I/um_iw[286]
+ tt_top1.branch\[0\].mux_I/um_iw[287] tt_top1.branch\[0\].mux_I/um_iw[28] tt_top1.branch\[0\].mux_I/um_iw[29]
+ tt_top1.branch\[0\].mux_I/um_iw[2] tt_top1.branch\[0\].mux_I/um_iw[30] tt_top1.branch\[0\].mux_I/um_iw[31]
+ tt_top1.branch\[0\].mux_I/um_iw[32] tt_top1.branch\[0\].mux_I/um_iw[33] tt_top1.branch\[0\].mux_I/um_iw[34]
+ tt_top1.branch\[0\].mux_I/um_iw[35] tt_top1.branch\[0\].mux_I/um_iw[36] tt_top1.branch\[0\].mux_I/um_iw[37]
+ tt_top1.branch\[0\].mux_I/um_iw[38] tt_top1.branch\[0\].mux_I/um_iw[39] tt_top1.branch\[0\].mux_I/um_iw[3]
+ tt_top1.branch\[0\].mux_I/um_iw[40] tt_top1.branch\[0\].mux_I/um_iw[41] tt_top1.branch\[0\].mux_I/um_iw[42]
+ tt_top1.branch\[0\].mux_I/um_iw[43] tt_top1.branch\[0\].mux_I/um_iw[44] tt_top1.branch\[0\].mux_I/um_iw[45]
+ tt_top1.branch\[0\].mux_I/um_iw[46] tt_top1.branch\[0\].mux_I/um_iw[47] tt_top1.branch\[0\].mux_I/um_iw[48]
+ tt_top1.branch\[0\].mux_I/um_iw[49] tt_top1.branch\[0\].mux_I/um_iw[4] tt_top1.branch\[0\].mux_I/um_iw[50]
+ tt_top1.branch\[0\].mux_I/um_iw[51] tt_top1.branch\[0\].mux_I/um_iw[52] tt_top1.branch\[0\].mux_I/um_iw[53]
+ tt_top1.branch\[0\].mux_I/um_iw[54] tt_top1.branch\[0\].mux_I/um_iw[55] tt_top1.branch\[0\].mux_I/um_iw[56]
+ tt_top1.branch\[0\].mux_I/um_iw[57] tt_top1.branch\[0\].mux_I/um_iw[58] tt_top1.branch\[0\].mux_I/um_iw[59]
+ tt_top1.branch\[0\].mux_I/um_iw[5] tt_top1.branch\[0\].mux_I/um_iw[60] tt_top1.branch\[0\].mux_I/um_iw[61]
+ tt_top1.branch\[0\].mux_I/um_iw[62] tt_top1.branch\[0\].mux_I/um_iw[63] tt_top1.branch\[0\].mux_I/um_iw[64]
+ tt_top1.branch\[0\].mux_I/um_iw[65] tt_top1.branch\[0\].mux_I/um_iw[66] tt_top1.branch\[0\].mux_I/um_iw[67]
+ tt_top1.branch\[0\].mux_I/um_iw[68] tt_top1.branch\[0\].mux_I/um_iw[69] tt_top1.branch\[0\].mux_I/um_iw[6]
+ tt_top1.branch\[0\].mux_I/um_iw[70] tt_top1.branch\[0\].mux_I/um_iw[71] tt_top1.branch\[0\].mux_I/um_iw[72]
+ tt_top1.branch\[0\].mux_I/um_iw[73] tt_top1.branch\[0\].mux_I/um_iw[74] tt_top1.branch\[0\].mux_I/um_iw[75]
+ tt_top1.branch\[0\].mux_I/um_iw[76] tt_top1.branch\[0\].mux_I/um_iw[77] tt_top1.branch\[0\].mux_I/um_iw[78]
+ tt_top1.branch\[0\].mux_I/um_iw[79] tt_top1.branch\[0\].mux_I/um_iw[7] tt_top1.branch\[0\].mux_I/um_iw[80]
+ tt_top1.branch\[0\].mux_I/um_iw[81] tt_top1.branch\[0\].mux_I/um_iw[82] tt_top1.branch\[0\].mux_I/um_iw[83]
+ tt_top1.branch\[0\].mux_I/um_iw[84] tt_top1.branch\[0\].mux_I/um_iw[85] tt_top1.branch\[0\].mux_I/um_iw[86]
+ tt_top1.branch\[0\].mux_I/um_iw[87] tt_top1.branch\[0\].mux_I/um_iw[88] tt_top1.branch\[0\].mux_I/um_iw[89]
+ tt_top1.branch\[0\].mux_I/um_iw[8] tt_top1.branch\[0\].mux_I/um_iw[90] tt_top1.branch\[0\].mux_I/um_iw[91]
+ tt_top1.branch\[0\].mux_I/um_iw[92] tt_top1.branch\[0\].mux_I/um_iw[93] tt_top1.branch\[0\].mux_I/um_iw[94]
+ tt_top1.branch\[0\].mux_I/um_iw[95] tt_top1.branch\[0\].mux_I/um_iw[96] tt_top1.branch\[0\].mux_I/um_iw[97]
+ tt_top1.branch\[0\].mux_I/um_iw[98] tt_top1.branch\[0\].mux_I/um_iw[99] tt_top1.branch\[0\].mux_I/um_iw[9]
+ tt_top1.branch\[0\].mux_I/um_k_zero[0] tt_top1.branch\[0\].mux_I/um_ow[263] tt_top1.branch\[0\].mux_I/um_k_zero[11]
+ tt_top1.branch\[0\].mux_I/um_ow[311] tt_top1.branch\[0\].mux_I/um_k_zero[13] tt_top1.branch\[0\].mux_I/um_ow[359]
+ tt_top1.branch\[0\].mux_I/um_k_zero[15] tt_top1.branch\[0\].mux_I/um_k_zero[1] tt_top1.branch\[0\].mux_I/um_k_zero[2]
+ tt_top1.branch\[0\].mux_I/um_k_zero[3] tt_top1.branch\[0\].mux_I/um_k_zero[4] tt_top1.branch\[0\].mux_I/um_k_zero[5]
+ tt_top1.branch\[0\].mux_I/um_k_zero[6] tt_top1.branch\[0\].mux_I/um_k_zero[7] tt_top1.branch\[0\].mux_I/um_k_zero[8]
+ tt_top1.branch\[0\].mux_I/um_k_zero[9] tt_top1.branch\[0\].mux_I/um_ow[0] tt_top1.branch\[0\].mux_I/um_ow[100]
+ tt_top1.branch\[0\].mux_I/um_ow[101] tt_top1.branch\[0\].mux_I/um_ow[102] tt_top1.branch\[0\].mux_I/um_ow[103]
+ tt_top1.branch\[0\].mux_I/um_ow[104] tt_top1.branch\[0\].mux_I/um_ow[105] tt_top1.branch\[0\].mux_I/um_ow[106]
+ tt_top1.branch\[0\].mux_I/um_ow[107] tt_top1.branch\[0\].mux_I/um_ow[108] tt_top1.branch\[0\].mux_I/um_ow[109]
+ tt_top1.branch\[0\].mux_I/um_ow[10] tt_top1.branch\[0\].mux_I/um_ow[110] tt_top1.branch\[0\].mux_I/um_ow[111]
+ tt_top1.branch\[0\].mux_I/um_ow[112] tt_top1.branch\[0\].mux_I/um_ow[113] tt_top1.branch\[0\].mux_I/um_ow[114]
+ tt_top1.branch\[0\].mux_I/um_ow[115] tt_top1.branch\[0\].mux_I/um_ow[116] tt_top1.branch\[0\].mux_I/um_ow[117]
+ tt_top1.branch\[0\].mux_I/um_ow[118] tt_top1.branch\[0\].mux_I/um_ow[119] tt_top1.branch\[0\].mux_I/um_ow[11]
+ tt_top1.branch\[0\].mux_I/um_ow[120] tt_top1.branch\[0\].mux_I/um_ow[121] tt_top1.branch\[0\].mux_I/um_ow[122]
+ tt_top1.branch\[0\].mux_I/um_ow[123] tt_top1.branch\[0\].mux_I/um_ow[124] tt_top1.branch\[0\].mux_I/um_ow[125]
+ tt_top1.branch\[0\].mux_I/um_ow[126] tt_top1.branch\[0\].mux_I/um_ow[127] tt_top1.branch\[0\].mux_I/um_ow[128]
+ tt_top1.branch\[0\].mux_I/um_ow[129] tt_top1.branch\[0\].mux_I/um_ow[12] tt_top1.branch\[0\].mux_I/um_ow[130]
+ tt_top1.branch\[0\].mux_I/um_ow[131] tt_top1.branch\[0\].mux_I/um_ow[132] tt_top1.branch\[0\].mux_I/um_ow[133]
+ tt_top1.branch\[0\].mux_I/um_ow[134] tt_top1.branch\[0\].mux_I/um_ow[135] tt_top1.branch\[0\].mux_I/um_ow[136]
+ tt_top1.branch\[0\].mux_I/um_ow[137] tt_top1.branch\[0\].mux_I/um_ow[138] tt_top1.branch\[0\].mux_I/um_ow[139]
+ tt_top1.branch\[0\].mux_I/um_ow[13] tt_top1.branch\[0\].mux_I/um_ow[140] tt_top1.branch\[0\].mux_I/um_ow[141]
+ tt_top1.branch\[0\].mux_I/um_ow[142] tt_top1.branch\[0\].mux_I/um_ow[143] tt_top1.branch\[0\].mux_I/um_ow[144]
+ tt_top1.branch\[0\].mux_I/um_ow[145] tt_top1.branch\[0\].mux_I/um_ow[146] tt_top1.branch\[0\].mux_I/um_ow[147]
+ tt_top1.branch\[0\].mux_I/um_ow[148] tt_top1.branch\[0\].mux_I/um_ow[149] tt_top1.branch\[0\].mux_I/um_ow[14]
+ tt_top1.branch\[0\].mux_I/um_ow[150] tt_top1.branch\[0\].mux_I/um_ow[151] tt_top1.branch\[0\].mux_I/um_ow[152]
+ tt_top1.branch\[0\].mux_I/um_ow[153] tt_top1.branch\[0\].mux_I/um_ow[154] tt_top1.branch\[0\].mux_I/um_ow[155]
+ tt_top1.branch\[0\].mux_I/um_ow[156] tt_top1.branch\[0\].mux_I/um_ow[157] tt_top1.branch\[0\].mux_I/um_ow[158]
+ tt_top1.branch\[0\].mux_I/um_ow[159] tt_top1.branch\[0\].mux_I/um_ow[15] tt_top1.branch\[0\].mux_I/um_ow[160]
+ tt_top1.branch\[0\].mux_I/um_ow[161] tt_top1.branch\[0\].mux_I/um_ow[162] tt_top1.branch\[0\].mux_I/um_ow[163]
+ tt_top1.branch\[0\].mux_I/um_ow[164] tt_top1.branch\[0\].mux_I/um_ow[165] tt_top1.branch\[0\].mux_I/um_ow[166]
+ tt_top1.branch\[0\].mux_I/um_ow[167] tt_top1.branch\[0\].mux_I/um_ow[168] tt_top1.branch\[0\].mux_I/um_ow[169]
+ tt_top1.branch\[0\].mux_I/um_ow[16] tt_top1.branch\[0\].mux_I/um_ow[170] tt_top1.branch\[0\].mux_I/um_ow[171]
+ tt_top1.branch\[0\].mux_I/um_ow[172] tt_top1.branch\[0\].mux_I/um_ow[173] tt_top1.branch\[0\].mux_I/um_ow[174]
+ tt_top1.branch\[0\].mux_I/um_ow[175] tt_top1.branch\[0\].mux_I/um_ow[176] tt_top1.branch\[0\].mux_I/um_ow[177]
+ tt_top1.branch\[0\].mux_I/um_ow[178] tt_top1.branch\[0\].mux_I/um_ow[179] tt_top1.branch\[0\].mux_I/um_ow[17]
+ tt_top1.branch\[0\].mux_I/um_ow[180] tt_top1.branch\[0\].mux_I/um_ow[181] tt_top1.branch\[0\].mux_I/um_ow[182]
+ tt_top1.branch\[0\].mux_I/um_ow[183] tt_top1.branch\[0\].mux_I/um_ow[184] tt_top1.branch\[0\].mux_I/um_ow[185]
+ tt_top1.branch\[0\].mux_I/um_ow[186] tt_top1.branch\[0\].mux_I/um_ow[187] tt_top1.branch\[0\].mux_I/um_ow[188]
+ tt_top1.branch\[0\].mux_I/um_ow[189] tt_top1.branch\[0\].mux_I/um_ow[18] tt_top1.branch\[0\].mux_I/um_ow[190]
+ tt_top1.branch\[0\].mux_I/um_ow[191] tt_top1.branch\[0\].mux_I/um_ow[192] tt_top1.branch\[0\].mux_I/um_ow[193]
+ tt_top1.branch\[0\].mux_I/um_ow[194] tt_top1.branch\[0\].mux_I/um_ow[195] tt_top1.branch\[0\].mux_I/um_ow[196]
+ tt_top1.branch\[0\].mux_I/um_ow[197] tt_top1.branch\[0\].mux_I/um_ow[198] tt_top1.branch\[0\].mux_I/um_ow[199]
+ tt_top1.branch\[0\].mux_I/um_ow[19] tt_top1.branch\[0\].mux_I/um_ow[1] tt_top1.branch\[0\].mux_I/um_ow[200]
+ tt_top1.branch\[0\].mux_I/um_ow[201] tt_top1.branch\[0\].mux_I/um_ow[202] tt_top1.branch\[0\].mux_I/um_ow[203]
+ tt_top1.branch\[0\].mux_I/um_ow[204] tt_top1.branch\[0\].mux_I/um_ow[205] tt_top1.branch\[0\].mux_I/um_ow[206]
+ tt_top1.branch\[0\].mux_I/um_ow[207] tt_top1.branch\[0\].mux_I/um_ow[208] tt_top1.branch\[0\].mux_I/um_ow[209]
+ tt_top1.branch\[0\].mux_I/um_ow[20] tt_top1.branch\[0\].mux_I/um_ow[210] tt_top1.branch\[0\].mux_I/um_ow[211]
+ tt_top1.branch\[0\].mux_I/um_ow[212] tt_top1.branch\[0\].mux_I/um_ow[213] tt_top1.branch\[0\].mux_I/um_ow[214]
+ tt_top1.branch\[0\].mux_I/um_ow[215] tt_top1.branch\[0\].mux_I/um_ow[216] tt_top1.branch\[0\].mux_I/um_ow[217]
+ tt_top1.branch\[0\].mux_I/um_ow[218] tt_top1.branch\[0\].mux_I/um_ow[219] tt_top1.branch\[0\].mux_I/um_ow[21]
+ tt_top1.branch\[0\].mux_I/um_ow[220] tt_top1.branch\[0\].mux_I/um_ow[221] tt_top1.branch\[0\].mux_I/um_ow[222]
+ tt_top1.branch\[0\].mux_I/um_ow[223] tt_top1.branch\[0\].mux_I/um_ow[224] tt_top1.branch\[0\].mux_I/um_ow[225]
+ tt_top1.branch\[0\].mux_I/um_ow[226] tt_top1.branch\[0\].mux_I/um_ow[227] tt_top1.branch\[0\].mux_I/um_ow[228]
+ tt_top1.branch\[0\].mux_I/um_ow[229] tt_top1.branch\[0\].mux_I/um_ow[22] tt_top1.branch\[0\].mux_I/um_ow[230]
+ tt_top1.branch\[0\].mux_I/um_ow[231] tt_top1.branch\[0\].mux_I/um_ow[232] tt_top1.branch\[0\].mux_I/um_ow[233]
+ tt_top1.branch\[0\].mux_I/um_ow[234] tt_top1.branch\[0\].mux_I/um_ow[235] tt_top1.branch\[0\].mux_I/um_ow[236]
+ tt_top1.branch\[0\].mux_I/um_ow[237] tt_top1.branch\[0\].mux_I/um_ow[238] tt_top1.branch\[0\].mux_I/um_ow[239]
+ tt_top1.branch\[0\].mux_I/um_ow[23] tt_top1.branch\[0\].mux_I/um_ow[263] tt_top1.branch\[0\].mux_I/um_ow[263]
+ tt_top1.branch\[0\].mux_I/um_ow[263] tt_top1.branch\[0\].mux_I/um_ow[263] tt_top1.branch\[0\].mux_I/um_ow[263]
+ tt_top1.branch\[0\].mux_I/um_ow[263] tt_top1.branch\[0\].mux_I/um_ow[263] tt_top1.branch\[0\].mux_I/um_ow[263]
+ tt_top1.branch\[0\].mux_I/um_ow[263] tt_top1.branch\[0\].mux_I/um_ow[263] tt_top1.branch\[0\].mux_I/um_ow[24]
+ tt_top1.branch\[0\].mux_I/um_ow[263] tt_top1.branch\[0\].mux_I/um_ow[263] tt_top1.branch\[0\].mux_I/um_ow[263]
+ tt_top1.branch\[0\].mux_I/um_ow[263] tt_top1.branch\[0\].mux_I/um_ow[263] tt_top1.branch\[0\].mux_I/um_ow[263]
+ tt_top1.branch\[0\].mux_I/um_ow[263] tt_top1.branch\[0\].mux_I/um_ow[263] tt_top1.branch\[0\].mux_I/um_ow[263]
+ tt_top1.branch\[0\].mux_I/um_ow[263] tt_top1.branch\[0\].mux_I/um_ow[25] tt_top1.branch\[0\].mux_I/um_ow[263]
+ tt_top1.branch\[0\].mux_I/um_ow[263] tt_top1.branch\[0\].mux_I/um_ow[263] tt_top1.branch\[0\].mux_I/um_ow[263]
+ tt_top1.branch\[0\].mux_I/um_ow[264] tt_top1.branch\[0\].mux_I/um_ow[265] tt_top1.branch\[0\].mux_I/um_ow[266]
+ tt_top1.branch\[0\].mux_I/um_ow[267] tt_top1.branch\[0\].mux_I/um_ow[268] tt_top1.branch\[0\].mux_I/um_ow[269]
+ tt_top1.branch\[0\].mux_I/um_ow[26] tt_top1.branch\[0\].mux_I/um_ow[270] tt_top1.branch\[0\].mux_I/um_ow[271]
+ tt_top1.branch\[0\].mux_I/um_ow[272] tt_top1.branch\[0\].mux_I/um_ow[273] tt_top1.branch\[0\].mux_I/um_ow[274]
+ tt_top1.branch\[0\].mux_I/um_ow[275] tt_top1.branch\[0\].mux_I/um_ow[276] tt_top1.branch\[0\].mux_I/um_ow[277]
+ tt_top1.branch\[0\].mux_I/um_ow[278] tt_top1.branch\[0\].mux_I/um_ow[279] tt_top1.branch\[0\].mux_I/um_ow[27]
+ tt_top1.branch\[0\].mux_I/um_ow[280] tt_top1.branch\[0\].mux_I/um_ow[281] tt_top1.branch\[0\].mux_I/um_ow[282]
+ tt_top1.branch\[0\].mux_I/um_ow[283] tt_top1.branch\[0\].mux_I/um_ow[284] tt_top1.branch\[0\].mux_I/um_ow[285]
+ tt_top1.branch\[0\].mux_I/um_ow[286] tt_top1.branch\[0\].mux_I/um_ow[287] tt_top1.branch\[0\].mux_I/um_ow[311]
+ tt_top1.branch\[0\].mux_I/um_ow[311] tt_top1.branch\[0\].mux_I/um_ow[28] tt_top1.branch\[0\].mux_I/um_ow[311]
+ tt_top1.branch\[0\].mux_I/um_ow[311] tt_top1.branch\[0\].mux_I/um_ow[311] tt_top1.branch\[0\].mux_I/um_ow[311]
+ tt_top1.branch\[0\].mux_I/um_ow[311] tt_top1.branch\[0\].mux_I/um_ow[311] tt_top1.branch\[0\].mux_I/um_ow[311]
+ tt_top1.branch\[0\].mux_I/um_ow[311] tt_top1.branch\[0\].mux_I/um_ow[311] tt_top1.branch\[0\].mux_I/um_ow[311]
+ tt_top1.branch\[0\].mux_I/um_ow[29] tt_top1.branch\[0\].mux_I/um_ow[2] tt_top1.branch\[0\].mux_I/um_ow[311]
+ tt_top1.branch\[0\].mux_I/um_ow[311] tt_top1.branch\[0\].mux_I/um_ow[311] tt_top1.branch\[0\].mux_I/um_ow[311]
+ tt_top1.branch\[0\].mux_I/um_ow[311] tt_top1.branch\[0\].mux_I/um_ow[311] tt_top1.branch\[0\].mux_I/um_ow[311]
+ tt_top1.branch\[0\].mux_I/um_ow[311] tt_top1.branch\[0\].mux_I/um_ow[311] tt_top1.branch\[0\].mux_I/um_ow[311]
+ tt_top1.branch\[0\].mux_I/um_ow[30] tt_top1.branch\[0\].mux_I/um_ow[311] tt_top1.branch\[0\].mux_I/um_ow[311]
+ tt_top1.branch\[0\].mux_I/um_ow[312] tt_top1.branch\[0\].mux_I/um_ow[313] tt_top1.branch\[0\].mux_I/um_ow[314]
+ tt_top1.branch\[0\].mux_I/um_ow[315] tt_top1.branch\[0\].mux_I/um_ow[316] tt_top1.branch\[0\].mux_I/um_ow[317]
+ tt_top1.branch\[0\].mux_I/um_ow[318] tt_top1.branch\[0\].mux_I/um_ow[319] tt_top1.branch\[0\].mux_I/um_ow[31]
+ tt_top1.branch\[0\].mux_I/um_ow[320] tt_top1.branch\[0\].mux_I/um_ow[321] tt_top1.branch\[0\].mux_I/um_ow[322]
+ tt_top1.branch\[0\].mux_I/um_ow[323] tt_top1.branch\[0\].mux_I/um_ow[324] tt_top1.branch\[0\].mux_I/um_ow[325]
+ tt_top1.branch\[0\].mux_I/um_ow[326] tt_top1.branch\[0\].mux_I/um_ow[327] tt_top1.branch\[0\].mux_I/um_ow[328]
+ tt_top1.branch\[0\].mux_I/um_ow[329] tt_top1.branch\[0\].mux_I/um_ow[32] tt_top1.branch\[0\].mux_I/um_ow[330]
+ tt_top1.branch\[0\].mux_I/um_ow[331] tt_top1.branch\[0\].mux_I/um_ow[332] tt_top1.branch\[0\].mux_I/um_ow[333]
+ tt_top1.branch\[0\].mux_I/um_ow[334] tt_top1.branch\[0\].mux_I/um_ow[335] tt_top1.branch\[0\].mux_I/um_ow[359]
+ tt_top1.branch\[0\].mux_I/um_ow[359] tt_top1.branch\[0\].mux_I/um_ow[359] tt_top1.branch\[0\].mux_I/um_ow[359]
+ tt_top1.branch\[0\].mux_I/um_ow[33] tt_top1.branch\[0\].mux_I/um_ow[359] tt_top1.branch\[0\].mux_I/um_ow[359]
+ tt_top1.branch\[0\].mux_I/um_ow[359] tt_top1.branch\[0\].mux_I/um_ow[359] tt_top1.branch\[0\].mux_I/um_ow[359]
+ tt_top1.branch\[0\].mux_I/um_ow[359] tt_top1.branch\[0\].mux_I/um_ow[359] tt_top1.branch\[0\].mux_I/um_ow[359]
+ tt_top1.branch\[0\].mux_I/um_ow[359] tt_top1.branch\[0\].mux_I/um_ow[359] tt_top1.branch\[0\].mux_I/um_ow[34]
+ tt_top1.branch\[0\].mux_I/um_ow[359] tt_top1.branch\[0\].mux_I/um_ow[359] tt_top1.branch\[0\].mux_I/um_ow[359]
+ tt_top1.branch\[0\].mux_I/um_ow[359] tt_top1.branch\[0\].mux_I/um_ow[359] tt_top1.branch\[0\].mux_I/um_ow[359]
+ tt_top1.branch\[0\].mux_I/um_ow[359] tt_top1.branch\[0\].mux_I/um_ow[359] tt_top1.branch\[0\].mux_I/um_ow[359]
+ tt_top1.branch\[0\].mux_I/um_ow[359] tt_top1.branch\[0\].mux_I/um_ow[35] tt_top1.branch\[0\].mux_I/um_ow[360]
+ tt_top1.branch\[0\].mux_I/um_ow[361] tt_top1.branch\[0\].mux_I/um_ow[362] tt_top1.branch\[0\].mux_I/um_ow[363]
+ tt_top1.branch\[0\].mux_I/um_ow[364] tt_top1.branch\[0\].mux_I/um_ow[365] tt_top1.branch\[0\].mux_I/um_ow[366]
+ tt_top1.branch\[0\].mux_I/um_ow[367] tt_top1.branch\[0\].mux_I/um_ow[368] tt_top1.branch\[0\].mux_I/um_ow[369]
+ tt_top1.branch\[0\].mux_I/um_ow[36] tt_top1.branch\[0\].mux_I/um_ow[370] tt_top1.branch\[0\].mux_I/um_ow[371]
+ tt_top1.branch\[0\].mux_I/um_ow[372] tt_top1.branch\[0\].mux_I/um_ow[373] tt_top1.branch\[0\].mux_I/um_ow[374]
+ tt_top1.branch\[0\].mux_I/um_ow[375] tt_top1.branch\[0\].mux_I/um_ow[376] tt_top1.branch\[0\].mux_I/um_ow[377]
+ tt_top1.branch\[0\].mux_I/um_ow[378] tt_top1.branch\[0\].mux_I/um_ow[379] tt_top1.branch\[0\].mux_I/um_ow[37]
+ tt_top1.branch\[0\].mux_I/um_ow[380] tt_top1.branch\[0\].mux_I/um_ow[381] tt_top1.branch\[0\].mux_I/um_ow[382]
+ tt_top1.branch\[0\].mux_I/um_ow[383] tt_top1.branch\[0\].mux_I/um_ow[38] tt_top1.branch\[0\].mux_I/um_ow[39]
+ tt_top1.branch\[0\].mux_I/um_ow[3] tt_top1.branch\[0\].mux_I/um_ow[40] tt_top1.branch\[0\].mux_I/um_ow[41]
+ tt_top1.branch\[0\].mux_I/um_ow[42] tt_top1.branch\[0\].mux_I/um_ow[43] tt_top1.branch\[0\].mux_I/um_ow[44]
+ tt_top1.branch\[0\].mux_I/um_ow[45] tt_top1.branch\[0\].mux_I/um_ow[46] tt_top1.branch\[0\].mux_I/um_ow[47]
+ tt_top1.branch\[0\].mux_I/um_ow[48] tt_top1.branch\[0\].mux_I/um_ow[49] tt_top1.branch\[0\].mux_I/um_ow[4]
+ tt_top1.branch\[0\].mux_I/um_ow[50] tt_top1.branch\[0\].mux_I/um_ow[51] tt_top1.branch\[0\].mux_I/um_ow[52]
+ tt_top1.branch\[0\].mux_I/um_ow[53] tt_top1.branch\[0\].mux_I/um_ow[54] tt_top1.branch\[0\].mux_I/um_ow[55]
+ tt_top1.branch\[0\].mux_I/um_ow[56] tt_top1.branch\[0\].mux_I/um_ow[57] tt_top1.branch\[0\].mux_I/um_ow[58]
+ tt_top1.branch\[0\].mux_I/um_ow[59] tt_top1.branch\[0\].mux_I/um_ow[5] tt_top1.branch\[0\].mux_I/um_ow[60]
+ tt_top1.branch\[0\].mux_I/um_ow[61] tt_top1.branch\[0\].mux_I/um_ow[62] tt_top1.branch\[0\].mux_I/um_ow[63]
+ tt_top1.branch\[0\].mux_I/um_ow[64] tt_top1.branch\[0\].mux_I/um_ow[65] tt_top1.branch\[0\].mux_I/um_ow[66]
+ tt_top1.branch\[0\].mux_I/um_ow[67] tt_top1.branch\[0\].mux_I/um_ow[68] tt_top1.branch\[0\].mux_I/um_ow[69]
+ tt_top1.branch\[0\].mux_I/um_ow[6] tt_top1.branch\[0\].mux_I/um_ow[70] tt_top1.branch\[0\].mux_I/um_ow[71]
+ tt_top1.branch\[0\].mux_I/um_ow[72] tt_top1.branch\[0\].mux_I/um_ow[73] tt_top1.branch\[0\].mux_I/um_ow[74]
+ tt_top1.branch\[0\].mux_I/um_ow[75] tt_top1.branch\[0\].mux_I/um_ow[76] tt_top1.branch\[0\].mux_I/um_ow[77]
+ tt_top1.branch\[0\].mux_I/um_ow[78] tt_top1.branch\[0\].mux_I/um_ow[79] tt_top1.branch\[0\].mux_I/um_ow[7]
+ tt_top1.branch\[0\].mux_I/um_ow[80] tt_top1.branch\[0\].mux_I/um_ow[81] tt_top1.branch\[0\].mux_I/um_ow[82]
+ tt_top1.branch\[0\].mux_I/um_ow[83] tt_top1.branch\[0\].mux_I/um_ow[84] tt_top1.branch\[0\].mux_I/um_ow[85]
+ tt_top1.branch\[0\].mux_I/um_ow[86] tt_top1.branch\[0\].mux_I/um_ow[87] tt_top1.branch\[0\].mux_I/um_ow[88]
+ tt_top1.branch\[0\].mux_I/um_ow[89] tt_top1.branch\[0\].mux_I/um_ow[8] tt_top1.branch\[0\].mux_I/um_ow[90]
+ tt_top1.branch\[0\].mux_I/um_ow[91] tt_top1.branch\[0\].mux_I/um_ow[92] tt_top1.branch\[0\].mux_I/um_ow[93]
+ tt_top1.branch\[0\].mux_I/um_ow[94] tt_top1.branch\[0\].mux_I/um_ow[95] tt_top1.branch\[0\].mux_I/um_ow[96]
+ tt_top1.branch\[0\].mux_I/um_ow[97] tt_top1.branch\[0\].mux_I/um_ow[98] tt_top1.branch\[0\].mux_I/um_ow[99]
+ tt_top1.branch\[0\].mux_I/um_ow[9] vccd1 vssd1 tt_mux
Xtt_top1.branch\[0\].col_um\[4\].um_bot_I.block_0_4.tt_um_I tt_top1.branch\[0\].mux_I/um_iw[144]
+ tt_top1.branch\[0\].mux_I/um_ena[8] tt_top1.branch\[0\].mux_I/um_iw[145] tt_top1.branch\[0\].mux_I/um_iw[146]
+ tt_top1.branch\[0\].mux_I/um_iw[147] tt_top1.branch\[0\].mux_I/um_iw[148] tt_top1.branch\[0\].mux_I/um_iw[149]
+ tt_top1.branch\[0\].mux_I/um_iw[150] tt_top1.branch\[0\].mux_I/um_iw[151] tt_top1.branch\[0\].mux_I/um_iw[152]
+ tt_top1.branch\[0\].mux_I/um_iw[153] tt_top1.branch\[0\].mux_I/um_iw[154] tt_top1.branch\[0\].mux_I/um_iw[155]
+ tt_top1.branch\[0\].mux_I/um_iw[156] tt_top1.branch\[0\].mux_I/um_iw[157] tt_top1.branch\[0\].mux_I/um_iw[158]
+ tt_top1.branch\[0\].mux_I/um_iw[159] tt_top1.branch\[0\].mux_I/um_iw[160] tt_top1.branch\[0\].mux_I/um_iw[161]
+ tt_top1.branch\[0\].mux_I/um_ow[208] tt_top1.branch\[0\].mux_I/um_ow[209] tt_top1.branch\[0\].mux_I/um_ow[210]
+ tt_top1.branch\[0\].mux_I/um_ow[211] tt_top1.branch\[0\].mux_I/um_ow[212] tt_top1.branch\[0\].mux_I/um_ow[213]
+ tt_top1.branch\[0\].mux_I/um_ow[214] tt_top1.branch\[0\].mux_I/um_ow[215] tt_top1.branch\[0\].mux_I/um_ow[200]
+ tt_top1.branch\[0\].mux_I/um_ow[201] tt_top1.branch\[0\].mux_I/um_ow[202] tt_top1.branch\[0\].mux_I/um_ow[203]
+ tt_top1.branch\[0\].mux_I/um_ow[204] tt_top1.branch\[0\].mux_I/um_ow[205] tt_top1.branch\[0\].mux_I/um_ow[206]
+ tt_top1.branch\[0\].mux_I/um_ow[207] tt_top1.branch\[0\].mux_I/um_ow[192] tt_top1.branch\[0\].mux_I/um_ow[193]
+ tt_top1.branch\[0\].mux_I/um_ow[194] tt_top1.branch\[0\].mux_I/um_ow[195] tt_top1.branch\[0\].mux_I/um_ow[196]
+ tt_top1.branch\[0\].mux_I/um_ow[197] tt_top1.branch\[0\].mux_I/um_ow[198] tt_top1.branch\[0\].mux_I/um_ow[199]
+ vccd1 vssd1 tt_um_urish_dffram
Xtt_top1.branch\[1\].col_um\[2\].um_top_I.block_1_18.tt_um_I tt_top1.branch\[1\].mux_I/um_iw[90]
+ tt_top1.branch\[1\].mux_I/um_ena[5] tt_top1.branch\[1\].mux_I/um_iw[91] tt_top1.branch\[1\].mux_I/um_iw[92]
+ tt_top1.branch\[1\].mux_I/um_iw[93] tt_top1.branch\[1\].mux_I/um_iw[94] tt_top1.branch\[1\].mux_I/um_iw[95]
+ tt_top1.branch\[1\].mux_I/um_iw[96] tt_top1.branch\[1\].mux_I/um_iw[97] tt_top1.branch\[1\].mux_I/um_iw[98]
+ tt_top1.branch\[1\].mux_I/um_iw[99] tt_top1.branch\[1\].mux_I/um_iw[100] tt_top1.branch\[1\].mux_I/um_iw[101]
+ tt_top1.branch\[1\].mux_I/um_iw[102] tt_top1.branch\[1\].mux_I/um_iw[103] tt_top1.branch\[1\].mux_I/um_iw[104]
+ tt_top1.branch\[1\].mux_I/um_iw[105] tt_top1.branch\[1\].mux_I/um_iw[106] tt_top1.branch\[1\].mux_I/um_iw[107]
+ tt_top1.branch\[1\].mux_I/um_ow[136] tt_top1.branch\[1\].mux_I/um_ow[137] tt_top1.branch\[1\].mux_I/um_ow[138]
+ tt_top1.branch\[1\].mux_I/um_ow[139] tt_top1.branch\[1\].mux_I/um_ow[140] tt_top1.branch\[1\].mux_I/um_ow[141]
+ tt_top1.branch\[1\].mux_I/um_ow[142] tt_top1.branch\[1\].mux_I/um_ow[143] tt_top1.branch\[1\].mux_I/um_ow[128]
+ tt_top1.branch\[1\].mux_I/um_ow[129] tt_top1.branch\[1\].mux_I/um_ow[130] tt_top1.branch\[1\].mux_I/um_ow[131]
+ tt_top1.branch\[1\].mux_I/um_ow[132] tt_top1.branch\[1\].mux_I/um_ow[133] tt_top1.branch\[1\].mux_I/um_ow[134]
+ tt_top1.branch\[1\].mux_I/um_ow[135] tt_top1.branch\[1\].mux_I/um_ow[120] tt_top1.branch\[1\].mux_I/um_ow[121]
+ tt_top1.branch\[1\].mux_I/um_ow[122] tt_top1.branch\[1\].mux_I/um_ow[123] tt_top1.branch\[1\].mux_I/um_ow[124]
+ tt_top1.branch\[1\].mux_I/um_ow[125] tt_top1.branch\[1\].mux_I/um_ow[126] tt_top1.branch\[1\].mux_I/um_ow[127]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[1\].col_um\[3\].um_bot_I.block_0_19.tt_um_I tt_top1.branch\[1\].mux_I/um_iw[108]
+ tt_top1.branch\[1\].mux_I/um_ena[6] tt_top1.branch\[1\].mux_I/um_iw[109] tt_top1.branch\[1\].mux_I/um_iw[110]
+ tt_top1.branch\[1\].mux_I/um_iw[111] tt_top1.branch\[1\].mux_I/um_iw[112] tt_top1.branch\[1\].mux_I/um_iw[113]
+ tt_top1.branch\[1\].mux_I/um_iw[114] tt_top1.branch\[1\].mux_I/um_iw[115] tt_top1.branch\[1\].mux_I/um_iw[116]
+ tt_top1.branch\[1\].mux_I/um_iw[117] tt_top1.branch\[1\].mux_I/um_iw[118] tt_top1.branch\[1\].mux_I/um_iw[119]
+ tt_top1.branch\[1\].mux_I/um_iw[120] tt_top1.branch\[1\].mux_I/um_iw[121] tt_top1.branch\[1\].mux_I/um_iw[122]
+ tt_top1.branch\[1\].mux_I/um_iw[123] tt_top1.branch\[1\].mux_I/um_iw[124] tt_top1.branch\[1\].mux_I/um_iw[125]
+ tt_top1.branch\[1\].mux_I/um_ow[160] tt_top1.branch\[1\].mux_I/um_ow[161] tt_top1.branch\[1\].mux_I/um_ow[162]
+ tt_top1.branch\[1\].mux_I/um_ow[163] tt_top1.branch\[1\].mux_I/um_ow[164] tt_top1.branch\[1\].mux_I/um_ow[165]
+ tt_top1.branch\[1\].mux_I/um_ow[166] tt_top1.branch\[1\].mux_I/um_ow[167] tt_top1.branch\[1\].mux_I/um_ow[152]
+ tt_top1.branch\[1\].mux_I/um_ow[153] tt_top1.branch\[1\].mux_I/um_ow[154] tt_top1.branch\[1\].mux_I/um_ow[155]
+ tt_top1.branch\[1\].mux_I/um_ow[156] tt_top1.branch\[1\].mux_I/um_ow[157] tt_top1.branch\[1\].mux_I/um_ow[158]
+ tt_top1.branch\[1\].mux_I/um_ow[159] tt_top1.branch\[1\].mux_I/um_ow[144] tt_top1.branch\[1\].mux_I/um_ow[145]
+ tt_top1.branch\[1\].mux_I/um_ow[146] tt_top1.branch\[1\].mux_I/um_ow[147] tt_top1.branch\[1\].mux_I/um_ow[148]
+ tt_top1.branch\[1\].mux_I/um_ow[149] tt_top1.branch\[1\].mux_I/um_ow[150] tt_top1.branch\[1\].mux_I/um_ow[151]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[0\].col_um\[3\].um_bot_I.block_0_3.tt_um_I tt_top1.branch\[0\].mux_I/um_iw[108]
+ tt_top1.branch\[0\].mux_I/um_ena[6] tt_top1.branch\[0\].mux_I/um_iw[109] tt_top1.branch\[0\].mux_I/um_iw[110]
+ tt_top1.branch\[0\].mux_I/um_iw[111] tt_top1.branch\[0\].mux_I/um_iw[112] tt_top1.branch\[0\].mux_I/um_iw[113]
+ tt_top1.branch\[0\].mux_I/um_iw[114] tt_top1.branch\[0\].mux_I/um_iw[115] tt_top1.branch\[0\].mux_I/um_iw[116]
+ tt_top1.branch\[0\].mux_I/um_iw[117] tt_top1.branch\[0\].mux_I/um_iw[118] tt_top1.branch\[0\].mux_I/um_iw[119]
+ tt_top1.branch\[0\].mux_I/um_iw[120] tt_top1.branch\[0\].mux_I/um_iw[121] tt_top1.branch\[0\].mux_I/um_iw[122]
+ tt_top1.branch\[0\].mux_I/um_iw[123] tt_top1.branch\[0\].mux_I/um_iw[124] tt_top1.branch\[0\].mux_I/um_iw[125]
+ tt_top1.branch\[0\].mux_I/um_ow[160] tt_top1.branch\[0\].mux_I/um_ow[161] tt_top1.branch\[0\].mux_I/um_ow[162]
+ tt_top1.branch\[0\].mux_I/um_ow[163] tt_top1.branch\[0\].mux_I/um_ow[164] tt_top1.branch\[0\].mux_I/um_ow[165]
+ tt_top1.branch\[0\].mux_I/um_ow[166] tt_top1.branch\[0\].mux_I/um_ow[167] tt_top1.branch\[0\].mux_I/um_ow[152]
+ tt_top1.branch\[0\].mux_I/um_ow[153] tt_top1.branch\[0\].mux_I/um_ow[154] tt_top1.branch\[0\].mux_I/um_ow[155]
+ tt_top1.branch\[0\].mux_I/um_ow[156] tt_top1.branch\[0\].mux_I/um_ow[157] tt_top1.branch\[0\].mux_I/um_ow[158]
+ tt_top1.branch\[0\].mux_I/um_ow[159] tt_top1.branch\[0\].mux_I/um_ow[144] tt_top1.branch\[0\].mux_I/um_ow[145]
+ tt_top1.branch\[0\].mux_I/um_ow[146] tt_top1.branch\[0\].mux_I/um_ow[147] tt_top1.branch\[0\].mux_I/um_ow[148]
+ tt_top1.branch\[0\].mux_I/um_ow[149] tt_top1.branch\[0\].mux_I/um_ow[150] tt_top1.branch\[0\].mux_I/um_ow[151]
+ vccd1 vssd1 tt_um_cam
Xtt_top1.branch\[0\].col_um\[2\].um_bot_I.block_0_2.tt_um_I tt_top1.branch\[0\].mux_I/um_iw[72]
+ tt_top1.branch\[0\].mux_I/um_ena[4] tt_top1.branch\[0\].mux_I/um_iw[73] tt_top1.branch\[0\].mux_I/um_iw[74]
+ tt_top1.branch\[0\].mux_I/um_iw[75] tt_top1.branch\[0\].mux_I/um_iw[76] tt_top1.branch\[0\].mux_I/um_iw[77]
+ tt_top1.branch\[0\].mux_I/um_iw[78] tt_top1.branch\[0\].mux_I/um_iw[79] tt_top1.branch\[0\].mux_I/um_iw[80]
+ tt_top1.branch\[0\].mux_I/um_iw[81] tt_top1.branch\[0\].mux_I/um_iw[82] tt_top1.branch\[0\].mux_I/um_iw[83]
+ tt_top1.branch\[0\].mux_I/um_iw[84] tt_top1.branch\[0\].mux_I/um_iw[85] tt_top1.branch\[0\].mux_I/um_iw[86]
+ tt_top1.branch\[0\].mux_I/um_iw[87] tt_top1.branch\[0\].mux_I/um_iw[88] tt_top1.branch\[0\].mux_I/um_iw[89]
+ tt_top1.branch\[0\].mux_I/um_ow[112] tt_top1.branch\[0\].mux_I/um_ow[113] tt_top1.branch\[0\].mux_I/um_ow[114]
+ tt_top1.branch\[0\].mux_I/um_ow[115] tt_top1.branch\[0\].mux_I/um_ow[116] tt_top1.branch\[0\].mux_I/um_ow[117]
+ tt_top1.branch\[0\].mux_I/um_ow[118] tt_top1.branch\[0\].mux_I/um_ow[119] tt_top1.branch\[0\].mux_I/um_ow[104]
+ tt_top1.branch\[0\].mux_I/um_ow[105] tt_top1.branch\[0\].mux_I/um_ow[106] tt_top1.branch\[0\].mux_I/um_ow[107]
+ tt_top1.branch\[0\].mux_I/um_ow[108] tt_top1.branch\[0\].mux_I/um_ow[109] tt_top1.branch\[0\].mux_I/um_ow[110]
+ tt_top1.branch\[0\].mux_I/um_ow[111] tt_top1.branch\[0\].mux_I/um_ow[96] tt_top1.branch\[0\].mux_I/um_ow[97]
+ tt_top1.branch\[0\].mux_I/um_ow[98] tt_top1.branch\[0\].mux_I/um_ow[99] tt_top1.branch\[0\].mux_I/um_ow[100]
+ tt_top1.branch\[0\].mux_I/um_ow[101] tt_top1.branch\[0\].mux_I/um_ow[102] tt_top1.branch\[0\].mux_I/um_ow[103]
+ vccd1 vssd1 tt_um_MichaelBell_hovalaag
Xtt_top1.branch\[1\].col_um\[5\].um_top_I.block_1_21.tt_um_I tt_top1.branch\[1\].mux_I/um_iw[198]
+ tt_top1.branch\[1\].mux_I/um_ena[11] tt_top1.branch\[1\].mux_I/um_iw[199] tt_top1.branch\[1\].mux_I/um_iw[200]
+ tt_top1.branch\[1\].mux_I/um_iw[201] tt_top1.branch\[1\].mux_I/um_iw[202] tt_top1.branch\[1\].mux_I/um_iw[203]
+ tt_top1.branch\[1\].mux_I/um_iw[204] tt_top1.branch\[1\].mux_I/um_iw[205] tt_top1.branch\[1\].mux_I/um_iw[206]
+ tt_top1.branch\[1\].mux_I/um_iw[207] tt_top1.branch\[1\].mux_I/um_iw[208] tt_top1.branch\[1\].mux_I/um_iw[209]
+ tt_top1.branch\[1\].mux_I/um_iw[210] tt_top1.branch\[1\].mux_I/um_iw[211] tt_top1.branch\[1\].mux_I/um_iw[212]
+ tt_top1.branch\[1\].mux_I/um_iw[213] tt_top1.branch\[1\].mux_I/um_iw[214] tt_top1.branch\[1\].mux_I/um_iw[215]
+ tt_top1.branch\[1\].mux_I/um_ow[280] tt_top1.branch\[1\].mux_I/um_ow[281] tt_top1.branch\[1\].mux_I/um_ow[282]
+ tt_top1.branch\[1\].mux_I/um_ow[283] tt_top1.branch\[1\].mux_I/um_ow[284] tt_top1.branch\[1\].mux_I/um_ow[285]
+ tt_top1.branch\[1\].mux_I/um_ow[286] tt_top1.branch\[1\].mux_I/um_ow[287] tt_top1.branch\[1\].mux_I/um_ow[272]
+ tt_top1.branch\[1\].mux_I/um_ow[273] tt_top1.branch\[1\].mux_I/um_ow[274] tt_top1.branch\[1\].mux_I/um_ow[275]
+ tt_top1.branch\[1\].mux_I/um_ow[276] tt_top1.branch\[1\].mux_I/um_ow[277] tt_top1.branch\[1\].mux_I/um_ow[278]
+ tt_top1.branch\[1\].mux_I/um_ow[279] tt_top1.branch\[1\].mux_I/um_ow[264] tt_top1.branch\[1\].mux_I/um_ow[265]
+ tt_top1.branch\[1\].mux_I/um_ow[266] tt_top1.branch\[1\].mux_I/um_ow[267] tt_top1.branch\[1\].mux_I/um_ow[268]
+ tt_top1.branch\[1\].mux_I/um_ow[269] tt_top1.branch\[1\].mux_I/um_ow[270] tt_top1.branch\[1\].mux_I/um_ow[271]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[1\].col_um\[6\].um_bot_I.block_0_22.tt_um_I tt_top1.branch\[1\].mux_I/um_iw[216]
+ tt_top1.branch\[1\].mux_I/um_ena[12] tt_top1.branch\[1\].mux_I/um_iw[217] tt_top1.branch\[1\].mux_I/um_iw[218]
+ tt_top1.branch\[1\].mux_I/um_iw[219] tt_top1.branch\[1\].mux_I/um_iw[220] tt_top1.branch\[1\].mux_I/um_iw[221]
+ tt_top1.branch\[1\].mux_I/um_iw[222] tt_top1.branch\[1\].mux_I/um_iw[223] tt_top1.branch\[1\].mux_I/um_iw[224]
+ tt_top1.branch\[1\].mux_I/um_iw[225] tt_top1.branch\[1\].mux_I/um_iw[226] tt_top1.branch\[1\].mux_I/um_iw[227]
+ tt_top1.branch\[1\].mux_I/um_iw[228] tt_top1.branch\[1\].mux_I/um_iw[229] tt_top1.branch\[1\].mux_I/um_iw[230]
+ tt_top1.branch\[1\].mux_I/um_iw[231] tt_top1.branch\[1\].mux_I/um_iw[232] tt_top1.branch\[1\].mux_I/um_iw[233]
+ tt_top1.branch\[1\].mux_I/um_ow[304] tt_top1.branch\[1\].mux_I/um_ow[305] tt_top1.branch\[1\].mux_I/um_ow[306]
+ tt_top1.branch\[1\].mux_I/um_ow[307] tt_top1.branch\[1\].mux_I/um_ow[308] tt_top1.branch\[1\].mux_I/um_ow[309]
+ tt_top1.branch\[1\].mux_I/um_ow[310] tt_top1.branch\[1\].mux_I/um_ow[311] tt_top1.branch\[1\].mux_I/um_ow[296]
+ tt_top1.branch\[1\].mux_I/um_ow[297] tt_top1.branch\[1\].mux_I/um_ow[298] tt_top1.branch\[1\].mux_I/um_ow[299]
+ tt_top1.branch\[1\].mux_I/um_ow[300] tt_top1.branch\[1\].mux_I/um_ow[301] tt_top1.branch\[1\].mux_I/um_ow[302]
+ tt_top1.branch\[1\].mux_I/um_ow[303] tt_top1.branch\[1\].mux_I/um_ow[288] tt_top1.branch\[1\].mux_I/um_ow[289]
+ tt_top1.branch\[1\].mux_I/um_ow[290] tt_top1.branch\[1\].mux_I/um_ow[291] tt_top1.branch\[1\].mux_I/um_ow[292]
+ tt_top1.branch\[1\].mux_I/um_ow[293] tt_top1.branch\[1\].mux_I/um_ow[294] tt_top1.branch\[1\].mux_I/um_ow[295]
+ vccd1 vssd1 tt_um_test
Xtt_top1.branch\[0\].col_um\[1\].um_bot_I.block_0_1.tt_um_I tt_top1.branch\[0\].mux_I/um_iw[36]
+ tt_top1.branch\[0\].mux_I/um_ena[2] tt_top1.branch\[0\].mux_I/um_iw[37] tt_top1.branch\[0\].mux_I/um_iw[38]
+ tt_top1.branch\[0\].mux_I/um_iw[39] tt_top1.branch\[0\].mux_I/um_iw[40] tt_top1.branch\[0\].mux_I/um_iw[41]
+ tt_top1.branch\[0\].mux_I/um_iw[42] tt_top1.branch\[0\].mux_I/um_iw[43] tt_top1.branch\[0\].mux_I/um_iw[44]
+ tt_top1.branch\[0\].mux_I/um_iw[45] tt_top1.branch\[0\].mux_I/um_iw[46] tt_top1.branch\[0\].mux_I/um_iw[47]
+ tt_top1.branch\[0\].mux_I/um_iw[48] tt_top1.branch\[0\].mux_I/um_iw[49] tt_top1.branch\[0\].mux_I/um_iw[50]
+ tt_top1.branch\[0\].mux_I/um_iw[51] tt_top1.branch\[0\].mux_I/um_iw[52] tt_top1.branch\[0\].mux_I/um_iw[53]
+ tt_top1.branch\[0\].mux_I/um_ow[64] tt_top1.branch\[0\].mux_I/um_ow[65] tt_top1.branch\[0\].mux_I/um_ow[66]
+ tt_top1.branch\[0\].mux_I/um_ow[67] tt_top1.branch\[0\].mux_I/um_ow[68] tt_top1.branch\[0\].mux_I/um_ow[69]
+ tt_top1.branch\[0\].mux_I/um_ow[70] tt_top1.branch\[0\].mux_I/um_ow[71] tt_top1.branch\[0\].mux_I/um_ow[56]
+ tt_top1.branch\[0\].mux_I/um_ow[57] tt_top1.branch\[0\].mux_I/um_ow[58] tt_top1.branch\[0\].mux_I/um_ow[59]
+ tt_top1.branch\[0\].mux_I/um_ow[60] tt_top1.branch\[0\].mux_I/um_ow[61] tt_top1.branch\[0\].mux_I/um_ow[62]
+ tt_top1.branch\[0\].mux_I/um_ow[63] tt_top1.branch\[0\].mux_I/um_ow[48] tt_top1.branch\[0\].mux_I/um_ow[49]
+ tt_top1.branch\[0\].mux_I/um_ow[50] tt_top1.branch\[0\].mux_I/um_ow[51] tt_top1.branch\[0\].mux_I/um_ow[52]
+ tt_top1.branch\[0\].mux_I/um_ow[53] tt_top1.branch\[0\].mux_I/um_ow[54] tt_top1.branch\[0\].mux_I/um_ow[55]
+ vccd1 vssd1 tt_um_urish_simon
.ends

