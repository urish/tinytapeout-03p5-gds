magic
tech sky130A
magscale 1 2
timestamp 1685642016
<< obsli1 >>
rect 1104 1071 35880 42449
<< obsm1 >>
rect 1104 1040 35880 42832
<< obsm2 >>
rect 1398 439 35586 43761
<< obsm3 >>
rect 790 443 36010 43757
<< metal4 >>
rect 798 42804 858 44064
rect 1166 42668 1226 44064
rect 1534 42804 1594 44064
rect 1902 43076 1962 44064
rect 2270 41308 2330 44064
rect 2638 42260 2698 44064
rect 3006 43076 3066 44064
rect 3374 42668 3434 44064
rect 3742 42124 3802 44064
rect 4110 43076 4170 44064
rect 4478 42804 4538 44064
rect 1902 0 1962 988
rect 2270 0 2330 3300
rect 2638 0 2698 3436
rect 3006 0 3066 444
rect 3374 0 3434 3436
rect 3742 0 3802 3300
rect 4208 1040 4528 42480
rect 4846 42396 4906 44064
rect 5214 41716 5274 44064
rect 5582 42804 5642 44064
rect 5950 41308 6010 44064
rect 6318 43212 6378 44064
rect 6686 42804 6746 44064
rect 7790 43864 7850 44064
rect 8158 42260 8218 44064
rect 8526 43076 8586 44064
rect 8894 42668 8954 44064
rect 9262 42668 9322 44064
rect 9630 41308 9690 44064
rect 9998 42668 10058 44064
rect 10366 42668 10426 44064
rect 10734 42804 10794 44064
rect 11102 42668 11162 44064
rect 11470 43076 11530 44064
rect 11838 42804 11898 44064
rect 12206 42668 12266 44064
rect 12574 43076 12634 44064
rect 12942 42940 13002 44064
rect 13310 42532 13370 44064
rect 13678 42804 13738 44064
rect 14046 43076 14106 44064
rect 14414 43076 14474 44064
rect 14782 43212 14842 44064
rect 15150 43212 15210 44064
rect 15518 43076 15578 44064
rect 15886 42804 15946 44064
rect 16254 43756 16314 44064
rect 16622 43076 16682 44064
rect 16990 43864 17050 44064
rect 18094 42532 18154 44064
rect 18462 39676 18522 44064
rect 18830 39948 18890 44064
rect 19198 42396 19258 44064
rect 19566 42940 19626 44064
rect 19934 42804 19994 44064
rect 4110 0 4170 852
rect 4478 0 4538 852
rect 4846 0 4906 988
rect 19568 1040 19888 42480
rect 20302 41308 20362 44064
rect 20670 42668 20730 44064
rect 21038 42124 21098 44064
rect 21406 41852 21466 44064
rect 21774 41852 21834 44064
rect 22142 42804 22202 44064
rect 22510 42804 22570 44064
rect 22878 42804 22938 44064
rect 23246 39948 23306 44064
rect 23614 41308 23674 44064
rect 23982 43076 24042 44064
rect 24350 38860 24410 44064
rect 24718 38724 24778 44064
rect 25086 42396 25146 44064
rect 25454 41852 25514 44064
rect 25822 43212 25882 44064
rect 26190 41370 26250 44064
rect 26558 42260 26618 44064
rect 26926 42396 26986 44064
rect 27294 42532 27354 44064
rect 27662 42668 27722 44064
rect 28030 41308 28090 44064
rect 28398 40764 28458 44064
rect 28766 38724 28826 44064
rect 29134 42260 29194 44064
rect 30054 39812 30114 44064
rect 30422 41036 30482 44064
rect 30790 43212 30850 44064
rect 31158 43076 31218 44064
rect 31526 40628 31586 44064
rect 31894 42804 31954 44064
rect 32262 42668 32322 44064
rect 32630 41308 32690 44064
rect 32998 43484 33058 44064
rect 33366 43076 33426 44064
rect 33734 43076 33794 44064
rect 34102 43212 34162 44064
rect 34470 41716 34530 44064
rect 34838 42668 34898 44064
rect 35206 42804 35266 44064
rect 34928 1040 35248 42480
rect 35574 41308 35634 44064
rect 35942 42260 36002 44064
rect 5214 0 5274 580
rect 5582 0 5642 444
rect 32814 0 32874 716
rect 33182 0 33242 716
<< obsm4 >>
rect 938 42724 1086 43757
rect 795 42588 1086 42724
rect 1306 42724 1454 43757
rect 1674 42996 1822 43757
rect 2042 42996 2190 43757
rect 1674 42724 2190 42996
rect 1306 42588 2190 42724
rect 795 41228 2190 42588
rect 2410 42180 2558 43757
rect 2778 42996 2926 43757
rect 3146 42996 3294 43757
rect 2778 42588 3294 42996
rect 3514 42588 3662 43757
rect 2778 42180 3662 42588
rect 2410 42044 3662 42180
rect 3882 42996 4030 43757
rect 4250 42996 4398 43757
rect 3882 42724 4398 42996
rect 4618 42724 4766 43757
rect 3882 42560 4766 42724
rect 3882 42044 4128 42560
rect 2410 41228 4128 42044
rect 795 3516 4128 41228
rect 795 3380 2558 3516
rect 795 1068 2190 3380
rect 795 443 1822 1068
rect 2042 443 2190 1068
rect 2410 443 2558 3380
rect 2778 524 3294 3516
rect 2778 443 2926 524
rect 3146 443 3294 524
rect 3514 3380 4128 3516
rect 3514 443 3662 3380
rect 3882 960 4128 3380
rect 4608 42316 4766 42560
rect 4986 42316 5134 43757
rect 4608 41636 5134 42316
rect 5354 42724 5502 43757
rect 5722 42724 5870 43757
rect 5354 41636 5870 42724
rect 4608 41228 5870 41636
rect 6090 43132 6238 43757
rect 6458 43132 6606 43757
rect 6090 42724 6606 43132
rect 6826 42724 8078 43757
rect 6090 42180 8078 42724
rect 8298 42996 8446 43757
rect 8666 42996 8814 43757
rect 8298 42588 8814 42996
rect 9034 42588 9182 43757
rect 9402 42588 9550 43757
rect 8298 42180 9550 42588
rect 6090 41228 9550 42180
rect 9770 42588 9918 43757
rect 10138 42588 10286 43757
rect 10506 42724 10654 43757
rect 10874 42724 11022 43757
rect 10506 42588 11022 42724
rect 11242 42996 11390 43757
rect 11610 42996 11758 43757
rect 11242 42724 11758 42996
rect 11978 42724 12126 43757
rect 11242 42588 12126 42724
rect 12346 42996 12494 43757
rect 12714 42996 12862 43757
rect 12346 42860 12862 42996
rect 13082 42860 13230 43757
rect 12346 42588 13230 42860
rect 9770 42452 13230 42588
rect 13450 42724 13598 43757
rect 13818 42996 13966 43757
rect 14186 42996 14334 43757
rect 14554 43132 14702 43757
rect 14922 43132 15070 43757
rect 15290 43132 15438 43757
rect 14554 42996 15438 43132
rect 15658 42996 15806 43757
rect 13818 42724 15806 42996
rect 16026 43676 16174 43757
rect 16394 43676 16542 43757
rect 16026 42996 16542 43676
rect 16762 42996 18014 43757
rect 16026 42724 18014 42996
rect 13450 42452 18014 42724
rect 18234 42452 18382 43757
rect 9770 41228 18382 42452
rect 4608 39596 18382 41228
rect 18602 39868 18750 43757
rect 18970 42316 19118 43757
rect 19338 42860 19486 43757
rect 19706 42860 19854 43757
rect 19338 42724 19854 42860
rect 20074 42724 20222 43757
rect 19338 42560 20222 42724
rect 19338 42316 19488 42560
rect 18970 39868 19488 42316
rect 18602 39596 19488 39868
rect 4608 1068 19488 39596
rect 4608 960 4766 1068
rect 3882 932 4766 960
rect 3882 443 4030 932
rect 4250 443 4398 932
rect 4618 443 4766 932
rect 4986 960 19488 1068
rect 19968 41228 20222 42560
rect 20442 42588 20590 43757
rect 20810 42588 20958 43757
rect 20442 42044 20958 42588
rect 21178 42044 21326 43757
rect 20442 41772 21326 42044
rect 21546 41772 21694 43757
rect 21914 42724 22062 43757
rect 22282 42724 22430 43757
rect 22650 42724 22798 43757
rect 23018 42724 23166 43757
rect 21914 41772 23166 42724
rect 20442 41228 23166 41772
rect 19968 39868 23166 41228
rect 23386 41228 23534 43757
rect 23754 42996 23902 43757
rect 24122 42996 24270 43757
rect 23754 41228 24270 42996
rect 23386 39868 24270 41228
rect 19968 38780 24270 39868
rect 24490 38780 24638 43757
rect 19968 38644 24638 38780
rect 24858 42316 25006 43757
rect 25226 42316 25374 43757
rect 24858 41772 25374 42316
rect 25594 43132 25742 43757
rect 25962 43132 26110 43757
rect 25594 41772 26110 43132
rect 24858 41290 26110 41772
rect 26330 42180 26478 43757
rect 26698 42316 26846 43757
rect 27066 42452 27214 43757
rect 27434 42588 27582 43757
rect 27802 42588 27950 43757
rect 27434 42452 27950 42588
rect 27066 42316 27950 42452
rect 26698 42180 27950 42316
rect 26330 41290 27950 42180
rect 24858 41228 27950 41290
rect 28170 41228 28318 43757
rect 24858 40684 28318 41228
rect 28538 40684 28686 43757
rect 24858 38644 28686 40684
rect 28906 42180 29054 43757
rect 29274 42180 29974 43757
rect 28906 39732 29974 42180
rect 30194 40956 30342 43757
rect 30562 43132 30710 43757
rect 30930 43132 31078 43757
rect 30562 42996 31078 43132
rect 31298 42996 31446 43757
rect 30562 40956 31446 42996
rect 30194 40548 31446 40956
rect 31666 42724 31814 43757
rect 32034 42724 32182 43757
rect 31666 42588 32182 42724
rect 32402 42588 32550 43757
rect 31666 41228 32550 42588
rect 32770 43404 32918 43757
rect 33138 43404 33286 43757
rect 32770 42996 33286 43404
rect 33506 42996 33654 43757
rect 33874 43132 34022 43757
rect 34242 43132 34390 43757
rect 33874 42996 34390 43132
rect 32770 41636 34390 42996
rect 34610 42588 34758 43757
rect 34978 42724 35126 43757
rect 35346 42724 35494 43757
rect 34978 42588 35494 42724
rect 34610 42560 35494 42588
rect 34610 41636 34848 42560
rect 32770 41228 34848 41636
rect 31666 40548 34848 41228
rect 30194 39732 34848 40548
rect 28906 38644 34848 39732
rect 19968 960 34848 38644
rect 35328 41228 35494 42560
rect 35714 42180 35862 43757
rect 35714 41228 36005 42180
rect 35328 960 36005 41228
rect 4986 796 36005 960
rect 4986 660 32734 796
rect 4986 443 5134 660
rect 5354 524 32734 660
rect 5354 443 5502 524
rect 5722 443 32734 524
rect 32954 443 33102 796
rect 33322 443 36005 796
<< labels >>
rlabel metal4 s 5582 0 5642 444 6 ctrl_ena
port 1 nsew signal input
rlabel metal4 s 5214 0 5274 580 6 ctrl_sel_inc
port 2 nsew signal input
rlabel metal4 s 4846 0 4906 988 6 ctrl_sel_rst_n
port 3 nsew signal input
rlabel metal4 s 4110 0 4170 852 6 k_one
port 4 nsew signal output
rlabel metal4 s 4478 0 4538 852 6 k_zero
port 5 nsew signal output
rlabel metal4 s 32814 0 32874 716 6 pad_ui_in[0]
port 6 nsew signal input
rlabel metal4 s 33182 0 33242 716 6 pad_ui_in[1]
port 7 nsew signal input
rlabel metal4 s 35942 42260 36002 44064 6 pad_ui_in[2]
port 8 nsew signal input
rlabel metal4 s 35574 41308 35634 44064 6 pad_ui_in[3]
port 9 nsew signal input
rlabel metal4 s 35206 42804 35266 44064 6 pad_ui_in[4]
port 10 nsew signal input
rlabel metal4 s 34838 42668 34898 44064 6 pad_ui_in[5]
port 11 nsew signal input
rlabel metal4 s 34470 41716 34530 44064 6 pad_ui_in[6]
port 12 nsew signal input
rlabel metal4 s 34102 43212 34162 44064 6 pad_ui_in[7]
port 13 nsew signal input
rlabel metal4 s 33734 43076 33794 44064 6 pad_ui_in[8]
port 14 nsew signal input
rlabel metal4 s 33366 43076 33426 44064 6 pad_ui_in[9]
port 15 nsew signal input
rlabel metal4 s 6318 43212 6378 44064 6 pad_uio_in[0]
port 16 nsew signal input
rlabel metal4 s 5214 41716 5274 44064 6 pad_uio_in[1]
port 17 nsew signal input
rlabel metal4 s 4110 43076 4170 44064 6 pad_uio_in[2]
port 18 nsew signal input
rlabel metal4 s 3006 43076 3066 44064 6 pad_uio_in[3]
port 19 nsew signal input
rlabel metal4 s 1902 43076 1962 44064 6 pad_uio_in[4]
port 20 nsew signal input
rlabel metal4 s 798 42804 858 44064 6 pad_uio_in[5]
port 21 nsew signal input
rlabel metal4 s 1902 0 1962 988 6 pad_uio_in[6]
port 22 nsew signal input
rlabel metal4 s 3006 0 3066 444 6 pad_uio_in[7]
port 23 nsew signal input
rlabel metal4 s 30054 39812 30114 44064 6 pad_uio_oe_n[0]
port 24 nsew signal output
rlabel metal4 s 5950 41308 6010 44064 6 pad_uio_oe_n[1]
port 25 nsew signal output
rlabel metal4 s 4846 42396 4906 44064 6 pad_uio_oe_n[2]
port 26 nsew signal output
rlabel metal4 s 3742 42124 3802 44064 6 pad_uio_oe_n[3]
port 27 nsew signal output
rlabel metal4 s 2638 42260 2698 44064 6 pad_uio_oe_n[4]
port 28 nsew signal output
rlabel metal4 s 1534 42804 1594 44064 6 pad_uio_oe_n[5]
port 29 nsew signal output
rlabel metal4 s 2638 0 2698 3436 6 pad_uio_oe_n[6]
port 30 nsew signal output
rlabel metal4 s 3742 0 3802 3300 6 pad_uio_oe_n[7]
port 31 nsew signal output
rlabel metal4 s 6686 42804 6746 44064 6 pad_uio_out[0]
port 32 nsew signal output
rlabel metal4 s 5582 42804 5642 44064 6 pad_uio_out[1]
port 33 nsew signal output
rlabel metal4 s 4478 42804 4538 44064 6 pad_uio_out[2]
port 34 nsew signal output
rlabel metal4 s 3374 42668 3434 44064 6 pad_uio_out[3]
port 35 nsew signal output
rlabel metal4 s 2270 41308 2330 44064 6 pad_uio_out[4]
port 36 nsew signal output
rlabel metal4 s 1166 42668 1226 44064 6 pad_uio_out[5]
port 37 nsew signal output
rlabel metal4 s 2270 0 2330 3300 6 pad_uio_out[6]
port 38 nsew signal output
rlabel metal4 s 3374 0 3434 3436 6 pad_uio_out[7]
port 39 nsew signal output
rlabel metal4 s 32998 43484 33058 44064 6 pad_uo_out[0]
port 40 nsew signal output
rlabel metal4 s 32630 41308 32690 44064 6 pad_uo_out[1]
port 41 nsew signal output
rlabel metal4 s 32262 42668 32322 44064 6 pad_uo_out[2]
port 42 nsew signal output
rlabel metal4 s 31894 42804 31954 44064 6 pad_uo_out[3]
port 43 nsew signal output
rlabel metal4 s 31526 40628 31586 44064 6 pad_uo_out[4]
port 44 nsew signal output
rlabel metal4 s 31158 43076 31218 44064 6 pad_uo_out[5]
port 45 nsew signal output
rlabel metal4 s 30790 43212 30850 44064 6 pad_uo_out[6]
port 46 nsew signal output
rlabel metal4 s 30422 41036 30482 44064 6 pad_uo_out[7]
port 47 nsew signal output
rlabel metal4 s 29134 42260 29194 44064 6 spine_iw[0]
port 48 nsew signal output
rlabel metal4 s 25454 41852 25514 44064 6 spine_iw[10]
port 49 nsew signal output
rlabel metal4 s 25086 42396 25146 44064 6 spine_iw[11]
port 50 nsew signal output
rlabel metal4 s 24718 38724 24778 44064 6 spine_iw[12]
port 51 nsew signal output
rlabel metal4 s 24350 38860 24410 44064 6 spine_iw[13]
port 52 nsew signal output
rlabel metal4 s 23982 43076 24042 44064 6 spine_iw[14]
port 53 nsew signal output
rlabel metal4 s 23614 41308 23674 44064 6 spine_iw[15]
port 54 nsew signal output
rlabel metal4 s 23246 39948 23306 44064 6 spine_iw[16]
port 55 nsew signal output
rlabel metal4 s 22878 42804 22938 44064 6 spine_iw[17]
port 56 nsew signal output
rlabel metal4 s 22510 42804 22570 44064 6 spine_iw[18]
port 57 nsew signal output
rlabel metal4 s 22142 42804 22202 44064 6 spine_iw[19]
port 58 nsew signal output
rlabel metal4 s 28766 38724 28826 44064 6 spine_iw[1]
port 59 nsew signal output
rlabel metal4 s 21774 41852 21834 44064 6 spine_iw[20]
port 60 nsew signal output
rlabel metal4 s 21406 41852 21466 44064 6 spine_iw[21]
port 61 nsew signal output
rlabel metal4 s 21038 42124 21098 44064 6 spine_iw[22]
port 62 nsew signal output
rlabel metal4 s 20670 42668 20730 44064 6 spine_iw[23]
port 63 nsew signal output
rlabel metal4 s 20302 41308 20362 44064 6 spine_iw[24]
port 64 nsew signal output
rlabel metal4 s 19934 42804 19994 44064 6 spine_iw[25]
port 65 nsew signal output
rlabel metal4 s 19566 42940 19626 44064 6 spine_iw[26]
port 66 nsew signal output
rlabel metal4 s 19198 42396 19258 44064 6 spine_iw[27]
port 67 nsew signal output
rlabel metal4 s 18830 39948 18890 44064 6 spine_iw[28]
port 68 nsew signal output
rlabel metal4 s 18462 39676 18522 44064 6 spine_iw[29]
port 69 nsew signal output
rlabel metal4 s 28398 40764 28458 44064 6 spine_iw[2]
port 70 nsew signal output
rlabel metal4 s 18094 42532 18154 44064 6 spine_iw[30]
port 71 nsew signal output
rlabel metal4 s 28030 41308 28090 44064 6 spine_iw[3]
port 72 nsew signal output
rlabel metal4 s 27662 42668 27722 44064 6 spine_iw[4]
port 73 nsew signal output
rlabel metal4 s 27294 42532 27354 44064 6 spine_iw[5]
port 74 nsew signal output
rlabel metal4 s 26926 42396 26986 44064 6 spine_iw[6]
port 75 nsew signal output
rlabel metal4 s 26558 42260 26618 44064 6 spine_iw[7]
port 76 nsew signal output
rlabel metal4 s 26190 41370 26250 44064 6 spine_iw[8]
port 77 nsew signal output
rlabel metal4 s 25822 43212 25882 44064 6 spine_iw[9]
port 78 nsew signal output
rlabel metal4 s 16990 43864 17050 44064 6 spine_ow[0]
port 79 nsew signal input
rlabel metal4 s 13310 42532 13370 44064 6 spine_ow[10]
port 80 nsew signal input
rlabel metal4 s 12942 42940 13002 44064 6 spine_ow[11]
port 81 nsew signal input
rlabel metal4 s 12574 43076 12634 44064 6 spine_ow[12]
port 82 nsew signal input
rlabel metal4 s 12206 42668 12266 44064 6 spine_ow[13]
port 83 nsew signal input
rlabel metal4 s 11838 42804 11898 44064 6 spine_ow[14]
port 84 nsew signal input
rlabel metal4 s 11470 43076 11530 44064 6 spine_ow[15]
port 85 nsew signal input
rlabel metal4 s 11102 42668 11162 44064 6 spine_ow[16]
port 86 nsew signal input
rlabel metal4 s 10734 42804 10794 44064 6 spine_ow[17]
port 87 nsew signal input
rlabel metal4 s 10366 42668 10426 44064 6 spine_ow[18]
port 88 nsew signal input
rlabel metal4 s 9998 42668 10058 44064 6 spine_ow[19]
port 89 nsew signal input
rlabel metal4 s 16622 43076 16682 44064 6 spine_ow[1]
port 90 nsew signal input
rlabel metal4 s 9630 41308 9690 44064 6 spine_ow[20]
port 91 nsew signal input
rlabel metal4 s 9262 42668 9322 44064 6 spine_ow[21]
port 92 nsew signal input
rlabel metal4 s 8894 42668 8954 44064 6 spine_ow[22]
port 93 nsew signal input
rlabel metal4 s 8526 43076 8586 44064 6 spine_ow[23]
port 94 nsew signal input
rlabel metal4 s 8158 42260 8218 44064 6 spine_ow[24]
port 95 nsew signal input
rlabel metal4 s 7790 43864 7850 44064 6 spine_ow[25]
port 96 nsew signal input
rlabel metal4 s 16254 43756 16314 44064 6 spine_ow[2]
port 97 nsew signal input
rlabel metal4 s 15886 42804 15946 44064 6 spine_ow[3]
port 98 nsew signal input
rlabel metal4 s 15518 43076 15578 44064 6 spine_ow[4]
port 99 nsew signal input
rlabel metal4 s 15150 43212 15210 44064 6 spine_ow[5]
port 100 nsew signal input
rlabel metal4 s 14782 43212 14842 44064 6 spine_ow[6]
port 101 nsew signal input
rlabel metal4 s 14414 43076 14474 44064 6 spine_ow[7]
port 102 nsew signal input
rlabel metal4 s 14046 43076 14106 44064 6 spine_ow[8]
port 103 nsew signal input
rlabel metal4 s 13678 42804 13738 44064 6 spine_ow[9]
port 104 nsew signal input
rlabel metal4 s 4208 1040 4528 42480 6 vccd1
port 105 nsew power bidirectional
rlabel metal4 s 34928 1040 35248 42480 6 vccd1
port 105 nsew power bidirectional
rlabel metal4 s 19568 1040 19888 42480 6 vssd1
port 106 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 37000 44000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 797218
string GDS_FILE /home/uri/p/tinytapeout-03p5-gds/openlane/tt_ctrl/runs/23_06_01_20_53/results/signoff/tt_ctrl.magic.gds
string GDS_START 76518
<< end >>

