VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_tomkeddie_a
  CLASS BLOCK ;
  FOREIGN tt_um_tomkeddie_a ;
  ORIGIN 0.000 0.000 ;
  SIZE 338.560 BY 220.320 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 206.850 158.850 220.320 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 162.230 219.320 162.530 220.320 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 214.020 155.170 220.320 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 217.420 151.490 220.320 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 216.740 147.810 220.320 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 219.320 144.130 220.320 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 219.320 140.450 220.320 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 219.320 136.770 220.320 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 219.320 133.090 220.320 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 219.320 129.410 220.320 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 219.320 125.730 220.320 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 219.320 122.050 220.320 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 219.320 118.370 220.320 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 219.320 114.690 220.320 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 219.320 111.010 220.320 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 219.320 107.330 220.320 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 219.320 103.650 220.320 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 219.320 99.970 220.320 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 219.320 96.290 220.320 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 218.780 33.730 220.320 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 218.100 30.050 220.320 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 218.780 26.370 220.320 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 218.780 22.690 220.320 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 214.700 19.010 220.320 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 211.300 15.330 220.320 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 214.700 11.650 220.320 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 211.300 7.970 220.320 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 218.100 63.170 220.320 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 218.780 59.490 220.320 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 218.780 55.810 220.320 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 214.700 52.130 220.320 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 218.780 48.450 220.320 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 218.780 44.770 220.320 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 218.780 41.090 220.320 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 218.780 37.410 220.320 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 218.780 92.610 220.320 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 218.780 88.930 220.320 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 214.700 85.250 220.320 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 218.100 81.570 220.320 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 218.780 77.890 220.320 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 218.780 74.210 220.320 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 214.700 70.530 220.320 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 218.780 66.850 220.320 ;
    END
  END uo_out[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 5.200 22.640 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 5.200 176.240 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 5.200 329.840 215.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 5.200 99.440 215.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 5.200 253.040 215.120 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 213.465 333.230 215.070 ;
        RECT 5.330 208.025 333.230 210.855 ;
        RECT 5.330 202.585 333.230 205.415 ;
        RECT 5.330 197.145 333.230 199.975 ;
        RECT 5.330 191.705 333.230 194.535 ;
        RECT 5.330 186.265 333.230 189.095 ;
        RECT 5.330 180.825 333.230 183.655 ;
        RECT 5.330 175.385 333.230 178.215 ;
        RECT 5.330 169.945 333.230 172.775 ;
        RECT 5.330 164.505 333.230 167.335 ;
        RECT 5.330 159.065 333.230 161.895 ;
        RECT 5.330 153.625 333.230 156.455 ;
        RECT 5.330 148.185 333.230 151.015 ;
        RECT 5.330 142.745 333.230 145.575 ;
        RECT 5.330 137.305 333.230 140.135 ;
        RECT 5.330 131.865 333.230 134.695 ;
        RECT 5.330 126.425 333.230 129.255 ;
        RECT 5.330 120.985 333.230 123.815 ;
        RECT 5.330 115.545 333.230 118.375 ;
        RECT 5.330 110.105 333.230 112.935 ;
        RECT 5.330 104.665 333.230 107.495 ;
        RECT 5.330 99.225 333.230 102.055 ;
        RECT 5.330 93.785 333.230 96.615 ;
        RECT 5.330 88.345 333.230 91.175 ;
        RECT 5.330 82.905 333.230 85.735 ;
        RECT 5.330 77.465 333.230 80.295 ;
        RECT 5.330 72.025 333.230 74.855 ;
        RECT 5.330 66.585 333.230 69.415 ;
        RECT 5.330 61.145 333.230 63.975 ;
        RECT 5.330 55.705 333.230 58.535 ;
        RECT 5.330 50.265 333.230 53.095 ;
        RECT 5.330 44.825 333.230 47.655 ;
        RECT 5.330 39.385 333.230 42.215 ;
        RECT 5.330 33.945 333.230 36.775 ;
        RECT 5.330 28.505 333.230 31.335 ;
        RECT 5.330 23.065 333.230 25.895 ;
        RECT 5.330 17.625 333.230 20.455 ;
        RECT 5.330 12.185 333.230 15.015 ;
        RECT 5.330 6.745 333.230 9.575 ;
      LAYER li1 ;
        RECT 5.520 5.355 333.040 214.965 ;
      LAYER met1 ;
        RECT 5.520 5.200 333.040 220.280 ;
      LAYER met2 ;
        RECT 7.920 5.255 329.810 220.310 ;
      LAYER met3 ;
        RECT 7.630 5.275 329.830 218.785 ;
      LAYER met4 ;
        RECT 8.370 214.300 10.950 218.785 ;
        RECT 12.050 214.300 14.630 218.785 ;
        RECT 8.370 210.900 14.630 214.300 ;
        RECT 15.730 214.300 18.310 218.785 ;
        RECT 19.410 218.380 21.990 218.785 ;
        RECT 23.090 218.380 25.670 218.785 ;
        RECT 26.770 218.380 29.350 218.785 ;
        RECT 19.410 217.700 29.350 218.380 ;
        RECT 30.450 218.380 33.030 218.785 ;
        RECT 34.130 218.380 36.710 218.785 ;
        RECT 37.810 218.380 40.390 218.785 ;
        RECT 41.490 218.380 44.070 218.785 ;
        RECT 45.170 218.380 47.750 218.785 ;
        RECT 48.850 218.380 51.430 218.785 ;
        RECT 30.450 217.700 51.430 218.380 ;
        RECT 19.410 215.520 51.430 217.700 ;
        RECT 19.410 214.300 20.640 215.520 ;
        RECT 15.730 210.900 20.640 214.300 ;
        RECT 7.655 91.295 20.640 210.900 ;
        RECT 23.040 214.300 51.430 215.520 ;
        RECT 52.530 218.380 55.110 218.785 ;
        RECT 56.210 218.380 58.790 218.785 ;
        RECT 59.890 218.380 62.470 218.785 ;
        RECT 52.530 217.700 62.470 218.380 ;
        RECT 63.570 218.380 66.150 218.785 ;
        RECT 67.250 218.380 69.830 218.785 ;
        RECT 63.570 217.700 69.830 218.380 ;
        RECT 52.530 214.300 69.830 217.700 ;
        RECT 70.930 218.380 73.510 218.785 ;
        RECT 74.610 218.380 77.190 218.785 ;
        RECT 78.290 218.380 80.870 218.785 ;
        RECT 70.930 217.700 80.870 218.380 ;
        RECT 81.970 217.700 84.550 218.785 ;
        RECT 70.930 214.300 84.550 217.700 ;
        RECT 85.650 218.380 88.230 218.785 ;
        RECT 89.330 218.380 91.910 218.785 ;
        RECT 93.010 218.380 147.110 218.785 ;
        RECT 85.650 216.340 147.110 218.380 ;
        RECT 148.210 217.020 150.790 218.785 ;
        RECT 151.890 217.020 154.470 218.785 ;
        RECT 148.210 216.340 154.470 217.020 ;
        RECT 85.650 215.520 154.470 216.340 ;
        RECT 85.650 214.300 97.440 215.520 ;
        RECT 23.040 91.295 97.440 214.300 ;
        RECT 99.840 213.620 154.470 215.520 ;
        RECT 155.570 213.620 158.150 218.785 ;
        RECT 99.840 206.450 158.150 213.620 ;
        RECT 159.250 215.520 234.305 218.785 ;
        RECT 159.250 206.450 174.240 215.520 ;
        RECT 99.840 91.295 174.240 206.450 ;
        RECT 176.640 91.295 234.305 215.520 ;
  END
END tt_um_tomkeddie_a
END LIBRARY

