* NGSPICE file created from tt_mux.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

.subckt tt_mux addr[0] addr[1] addr[2] addr[3] addr[4] k_one k_zero spine_iw[0] spine_iw[10]
+ spine_iw[11] spine_iw[12] spine_iw[13] spine_iw[14] spine_iw[15] spine_iw[16] spine_iw[17]
+ spine_iw[18] spine_iw[19] spine_iw[1] spine_iw[20] spine_iw[21] spine_iw[22] spine_iw[23]
+ spine_iw[24] spine_iw[25] spine_iw[26] spine_iw[27] spine_iw[28] spine_iw[29] spine_iw[2]
+ spine_iw[30] spine_iw[3] spine_iw[4] spine_iw[5] spine_iw[6] spine_iw[7] spine_iw[8]
+ spine_iw[9] spine_ow[0] spine_ow[10] spine_ow[11] spine_ow[12] spine_ow[13] spine_ow[14]
+ spine_ow[15] spine_ow[16] spine_ow[17] spine_ow[18] spine_ow[19] spine_ow[1] spine_ow[20]
+ spine_ow[21] spine_ow[22] spine_ow[23] spine_ow[24] spine_ow[25] spine_ow[2] spine_ow[3]
+ spine_ow[4] spine_ow[5] spine_ow[6] spine_ow[7] spine_ow[8] spine_ow[9] um_ena[0]
+ um_ena[10] um_ena[11] um_ena[12] um_ena[13] um_ena[14] um_ena[15] um_ena[1] um_ena[2]
+ um_ena[3] um_ena[4] um_ena[5] um_ena[6] um_ena[7] um_ena[8] um_ena[9] um_iw[0] um_iw[100]
+ um_iw[101] um_iw[102] um_iw[103] um_iw[104] um_iw[105] um_iw[106] um_iw[107] um_iw[108]
+ um_iw[109] um_iw[10] um_iw[110] um_iw[111] um_iw[112] um_iw[113] um_iw[114] um_iw[115]
+ um_iw[116] um_iw[117] um_iw[118] um_iw[119] um_iw[11] um_iw[120] um_iw[121] um_iw[122]
+ um_iw[123] um_iw[124] um_iw[125] um_iw[126] um_iw[127] um_iw[128] um_iw[129] um_iw[12]
+ um_iw[130] um_iw[131] um_iw[132] um_iw[133] um_iw[134] um_iw[135] um_iw[136] um_iw[137]
+ um_iw[138] um_iw[139] um_iw[13] um_iw[140] um_iw[141] um_iw[142] um_iw[143] um_iw[144]
+ um_iw[145] um_iw[146] um_iw[147] um_iw[148] um_iw[149] um_iw[14] um_iw[150] um_iw[151]
+ um_iw[152] um_iw[153] um_iw[154] um_iw[155] um_iw[156] um_iw[157] um_iw[158] um_iw[159]
+ um_iw[15] um_iw[160] um_iw[161] um_iw[162] um_iw[163] um_iw[164] um_iw[165] um_iw[166]
+ um_iw[167] um_iw[168] um_iw[169] um_iw[16] um_iw[170] um_iw[171] um_iw[172] um_iw[173]
+ um_iw[174] um_iw[175] um_iw[176] um_iw[177] um_iw[178] um_iw[179] um_iw[17] um_iw[180]
+ um_iw[181] um_iw[182] um_iw[183] um_iw[184] um_iw[185] um_iw[186] um_iw[187] um_iw[188]
+ um_iw[189] um_iw[18] um_iw[190] um_iw[191] um_iw[192] um_iw[193] um_iw[194] um_iw[195]
+ um_iw[196] um_iw[197] um_iw[198] um_iw[199] um_iw[19] um_iw[1] um_iw[200] um_iw[201]
+ um_iw[202] um_iw[203] um_iw[204] um_iw[205] um_iw[206] um_iw[207] um_iw[208] um_iw[209]
+ um_iw[20] um_iw[210] um_iw[211] um_iw[212] um_iw[213] um_iw[214] um_iw[215] um_iw[216]
+ um_iw[217] um_iw[218] um_iw[219] um_iw[21] um_iw[220] um_iw[221] um_iw[222] um_iw[223]
+ um_iw[224] um_iw[225] um_iw[226] um_iw[227] um_iw[228] um_iw[229] um_iw[22] um_iw[230]
+ um_iw[231] um_iw[232] um_iw[233] um_iw[234] um_iw[235] um_iw[236] um_iw[237] um_iw[238]
+ um_iw[239] um_iw[23] um_iw[240] um_iw[241] um_iw[242] um_iw[243] um_iw[244] um_iw[245]
+ um_iw[246] um_iw[247] um_iw[248] um_iw[249] um_iw[24] um_iw[250] um_iw[251] um_iw[252]
+ um_iw[253] um_iw[254] um_iw[255] um_iw[256] um_iw[257] um_iw[258] um_iw[259] um_iw[25]
+ um_iw[260] um_iw[261] um_iw[262] um_iw[263] um_iw[264] um_iw[265] um_iw[266] um_iw[267]
+ um_iw[268] um_iw[269] um_iw[26] um_iw[270] um_iw[271] um_iw[272] um_iw[273] um_iw[274]
+ um_iw[275] um_iw[276] um_iw[277] um_iw[278] um_iw[279] um_iw[27] um_iw[280] um_iw[281]
+ um_iw[282] um_iw[283] um_iw[284] um_iw[285] um_iw[286] um_iw[287] um_iw[28] um_iw[29]
+ um_iw[2] um_iw[30] um_iw[31] um_iw[32] um_iw[33] um_iw[34] um_iw[35] um_iw[36] um_iw[37]
+ um_iw[38] um_iw[39] um_iw[3] um_iw[40] um_iw[41] um_iw[42] um_iw[43] um_iw[44] um_iw[45]
+ um_iw[46] um_iw[47] um_iw[48] um_iw[49] um_iw[4] um_iw[50] um_iw[51] um_iw[52] um_iw[53]
+ um_iw[54] um_iw[55] um_iw[56] um_iw[57] um_iw[58] um_iw[59] um_iw[5] um_iw[60] um_iw[61]
+ um_iw[62] um_iw[63] um_iw[64] um_iw[65] um_iw[66] um_iw[67] um_iw[68] um_iw[69]
+ um_iw[6] um_iw[70] um_iw[71] um_iw[72] um_iw[73] um_iw[74] um_iw[75] um_iw[76] um_iw[77]
+ um_iw[78] um_iw[79] um_iw[7] um_iw[80] um_iw[81] um_iw[82] um_iw[83] um_iw[84] um_iw[85]
+ um_iw[86] um_iw[87] um_iw[88] um_iw[89] um_iw[8] um_iw[90] um_iw[91] um_iw[92] um_iw[93]
+ um_iw[94] um_iw[95] um_iw[96] um_iw[97] um_iw[98] um_iw[99] um_iw[9] um_k_zero[0]
+ um_k_zero[10] um_k_zero[11] um_k_zero[12] um_k_zero[13] um_k_zero[14] um_k_zero[15]
+ um_k_zero[1] um_k_zero[2] um_k_zero[3] um_k_zero[4] um_k_zero[5] um_k_zero[6] um_k_zero[7]
+ um_k_zero[8] um_k_zero[9] um_ow[0] um_ow[100] um_ow[101] um_ow[102] um_ow[103] um_ow[104]
+ um_ow[105] um_ow[106] um_ow[107] um_ow[108] um_ow[109] um_ow[10] um_ow[110] um_ow[111]
+ um_ow[112] um_ow[113] um_ow[114] um_ow[115] um_ow[116] um_ow[117] um_ow[118] um_ow[119]
+ um_ow[11] um_ow[120] um_ow[121] um_ow[122] um_ow[123] um_ow[124] um_ow[125] um_ow[126]
+ um_ow[127] um_ow[128] um_ow[129] um_ow[12] um_ow[130] um_ow[131] um_ow[132] um_ow[133]
+ um_ow[134] um_ow[135] um_ow[136] um_ow[137] um_ow[138] um_ow[139] um_ow[13] um_ow[140]
+ um_ow[141] um_ow[142] um_ow[143] um_ow[144] um_ow[145] um_ow[146] um_ow[147] um_ow[148]
+ um_ow[149] um_ow[14] um_ow[150] um_ow[151] um_ow[152] um_ow[153] um_ow[154] um_ow[155]
+ um_ow[156] um_ow[157] um_ow[158] um_ow[159] um_ow[15] um_ow[160] um_ow[161] um_ow[162]
+ um_ow[163] um_ow[164] um_ow[165] um_ow[166] um_ow[167] um_ow[168] um_ow[169] um_ow[16]
+ um_ow[170] um_ow[171] um_ow[172] um_ow[173] um_ow[174] um_ow[175] um_ow[176] um_ow[177]
+ um_ow[178] um_ow[179] um_ow[17] um_ow[180] um_ow[181] um_ow[182] um_ow[183] um_ow[184]
+ um_ow[185] um_ow[186] um_ow[187] um_ow[188] um_ow[189] um_ow[18] um_ow[190] um_ow[191]
+ um_ow[192] um_ow[193] um_ow[194] um_ow[195] um_ow[196] um_ow[197] um_ow[198] um_ow[199]
+ um_ow[19] um_ow[1] um_ow[200] um_ow[201] um_ow[202] um_ow[203] um_ow[204] um_ow[205]
+ um_ow[206] um_ow[207] um_ow[208] um_ow[209] um_ow[20] um_ow[210] um_ow[211] um_ow[212]
+ um_ow[213] um_ow[214] um_ow[215] um_ow[216] um_ow[217] um_ow[218] um_ow[219] um_ow[21]
+ um_ow[220] um_ow[221] um_ow[222] um_ow[223] um_ow[224] um_ow[225] um_ow[226] um_ow[227]
+ um_ow[228] um_ow[229] um_ow[22] um_ow[230] um_ow[231] um_ow[232] um_ow[233] um_ow[234]
+ um_ow[235] um_ow[236] um_ow[237] um_ow[238] um_ow[239] um_ow[23] um_ow[240] um_ow[241]
+ um_ow[242] um_ow[243] um_ow[244] um_ow[245] um_ow[246] um_ow[247] um_ow[248] um_ow[249]
+ um_ow[24] um_ow[250] um_ow[251] um_ow[252] um_ow[253] um_ow[254] um_ow[255] um_ow[256]
+ um_ow[257] um_ow[258] um_ow[259] um_ow[25] um_ow[260] um_ow[261] um_ow[262] um_ow[263]
+ um_ow[264] um_ow[265] um_ow[266] um_ow[267] um_ow[268] um_ow[269] um_ow[26] um_ow[270]
+ um_ow[271] um_ow[272] um_ow[273] um_ow[274] um_ow[275] um_ow[276] um_ow[277] um_ow[278]
+ um_ow[279] um_ow[27] um_ow[280] um_ow[281] um_ow[282] um_ow[283] um_ow[284] um_ow[285]
+ um_ow[286] um_ow[287] um_ow[288] um_ow[289] um_ow[28] um_ow[290] um_ow[291] um_ow[292]
+ um_ow[293] um_ow[294] um_ow[295] um_ow[296] um_ow[297] um_ow[298] um_ow[299] um_ow[29]
+ um_ow[2] um_ow[300] um_ow[301] um_ow[302] um_ow[303] um_ow[304] um_ow[305] um_ow[306]
+ um_ow[307] um_ow[308] um_ow[309] um_ow[30] um_ow[310] um_ow[311] um_ow[312] um_ow[313]
+ um_ow[314] um_ow[315] um_ow[316] um_ow[317] um_ow[318] um_ow[319] um_ow[31] um_ow[320]
+ um_ow[321] um_ow[322] um_ow[323] um_ow[324] um_ow[325] um_ow[326] um_ow[327] um_ow[328]
+ um_ow[329] um_ow[32] um_ow[330] um_ow[331] um_ow[332] um_ow[333] um_ow[334] um_ow[335]
+ um_ow[336] um_ow[337] um_ow[338] um_ow[339] um_ow[33] um_ow[340] um_ow[341] um_ow[342]
+ um_ow[343] um_ow[344] um_ow[345] um_ow[346] um_ow[347] um_ow[348] um_ow[349] um_ow[34]
+ um_ow[350] um_ow[351] um_ow[352] um_ow[353] um_ow[354] um_ow[355] um_ow[356] um_ow[357]
+ um_ow[358] um_ow[359] um_ow[35] um_ow[360] um_ow[361] um_ow[362] um_ow[363] um_ow[364]
+ um_ow[365] um_ow[366] um_ow[367] um_ow[368] um_ow[369] um_ow[36] um_ow[370] um_ow[371]
+ um_ow[372] um_ow[373] um_ow[374] um_ow[375] um_ow[376] um_ow[377] um_ow[378] um_ow[379]
+ um_ow[37] um_ow[380] um_ow[381] um_ow[382] um_ow[383] um_ow[38] um_ow[39] um_ow[3]
+ um_ow[40] um_ow[41] um_ow[42] um_ow[43] um_ow[44] um_ow[45] um_ow[46] um_ow[47]
+ um_ow[48] um_ow[49] um_ow[4] um_ow[50] um_ow[51] um_ow[52] um_ow[53] um_ow[54] um_ow[55]
+ um_ow[56] um_ow[57] um_ow[58] um_ow[59] um_ow[5] um_ow[60] um_ow[61] um_ow[62] um_ow[63]
+ um_ow[64] um_ow[65] um_ow[66] um_ow[67] um_ow[68] um_ow[69] um_ow[6] um_ow[70] um_ow[71]
+ um_ow[72] um_ow[73] um_ow[74] um_ow[75] um_ow[76] um_ow[77] um_ow[78] um_ow[79]
+ um_ow[7] um_ow[80] um_ow[81] um_ow[82] um_ow[83] um_ow[84] um_ow[85] um_ow[86] um_ow[87]
+ um_ow[88] um_ow[89] um_ow[8] um_ow[90] um_ow[91] um_ow[92] um_ow[93] um_ow[94] um_ow[95]
+ um_ow[96] um_ow[97] um_ow[98] um_ow[99] um_ow[9] vccd1 vssd1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0367_ _0040_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_2673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[4\].zbuf_bot_iw_I\[10\].genblk1.cell0_I net509 net443 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_bot_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0985_ col\[0\].genblk1.mux4_I\[14\].x _0205_ vssd1 vssd1 vccd1 vccd1 bus_ow\[14\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_14_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.mux4_I\[17\].cell0_I net263 net289 net316 net342 net475 net462 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[17\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_1_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0419_ _0071_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_2334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0770_ col\[4\].zbuf_top_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[167] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[0\].zbuf_bot_iw_I\[5\].genblk1.cell0_I net485 net448 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_bot_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[4\].genblk1.mux4_I\[8\].cell0_I net147 net173 net199 net226 net470 net458 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[8\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_7_2908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0968_ bus_ow\[21\] _0188_ vssd1 vssd1 vccd1 vccd1 spine_ow[22] sky130_fd_sc_hd__ebufn_8
XFILLER_0_6_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].zbuf_bot_iw_I\[0\].genblk1.cell0_I net511 net446 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_bot_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XFILLER_0_15_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0899_ col\[4\].zbuf_bot_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[8] sky130_fd_sc_hd__buf_2
XFILLER_0_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout480 col\[0\].zbuf_bot_iw_I\[8\].a vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_4
Xfanout491 col\[0\].zbuf_bot_iw_I\[2\].a vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__buf_6
Xcol\[0\].genblk1.mux4_I\[6\].cell0_I net385 net268 net368 net394 net466 net452 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[6\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_9_2042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0822_ col\[6\].zbuf_bot_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[219] sky130_fd_sc_hd__buf_2
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0753_ col\[4\].zbuf_bot_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[150] sky130_fd_sc_hd__buf_2
XFILLER_0_3_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0684_ col\[2\].zbuf_bot_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[81] sky130_fd_sc_hd__buf_2
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[3\].zbuf_top_iw_I\[17\].genblk1.cell0_I net495 net425 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_2136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1021_ col\[4\].genblk1.mux4_I\[2\].x _0241_ vssd1 vssd1 vccd1 vccd1 bus_ow\[2\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_2_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_2681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[3\].zbuf_bot_iw_I\[8\].genblk1.cell0_I net479 net427 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_bot_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0805_ col\[5\].zbuf_top_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[202] sky130_fd_sc_hd__buf_2
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0736_ col\[3\].zbuf_top_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[133] sky130_fd_sc_hd__buf_2
XFILLER_0_0_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0667_ col\[1\].zbuf_top_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[64] sky130_fd_sc_hd__buf_2
X_0598_ net474 net460 _0264_ zbuf_bus_ena_I.z vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__or4b_1
XFILLER_0_7_2513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_2557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[5\].zbuf_bot_iw_I\[3\].genblk1.cell0_I net490 net422 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_bot_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_2178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput301 um_ow[33] vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_2
Xinput312 um_ow[34] vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__clkbuf_2
Xinput334 um_ow[36] vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_2
Xinput323 um_ow[35] vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__clkbuf_2
Xinput345 um_ow[37] vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__clkbuf_2
Xinput356 um_ow[43] vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__clkbuf_2
Xinput378 um_ow[63] vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_1
Xinput367 um_ow[53] vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__clkbuf_1
Xinput389 um_ow[73] vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_2001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_5 col\[0\].zbuf_bot_iw_I\[13\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0521_ _0129_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0452_ _0083_ _0089_ _0084_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__or3b_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0383_ _0051_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_2732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1004_ col\[2\].genblk1.mux4_I\[9\].x _0224_ vssd1 vssd1 vccd1 vccd1 bus_ow\[9\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_14_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[5\].zbuf_top_iw_I\[16\].genblk1.cell0_I net498 net419 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[16\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_iw_I\[7\].genblk1.cell0_I net481 net432 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0719_ col\[3\].zbuf_bot_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[116] sky130_fd_sc_hd__buf_2
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[2\].genblk1.mux4_I\[9\].cell0_I net41 net67 net94 net120 net468 net454 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[9\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_9_1929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[3\].zbuf_top_iw_I\[2\].genblk1.cell0_I net491 net426 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput120 um_ow[177] vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__clkbuf_1
Xinput131 um_ow[187] vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__clkbuf_1
Xinput142 um_ow[197] vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_1
Xinput153 um_ow[206] vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__clkbuf_1
Xinput175 um_ow[226] vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_1
Xinput186 um_ow[236] vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_1
Xinput164 um_ow[216] vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_1
Xinput197 um_ow[246] vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_8_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_2039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].genblk1.mux4_I\[12\].cell0_I net44 net71 net97 net124 net468 net454 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[12\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_15_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_2673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_sel_I\[4\].genblk1.cell0_I net30 net516 vssd1 vssd1 vccd1 vccd1 zbuf_bus_sel_I\[4\].genblk1.l
+ sky130_fd_sc_hd__and2_2
XFILLER_0_14_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0504_ _0119_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0435_ _0075_ _0076_ _0077_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__or3b_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0366_ _0001_ _0005_ _0008_ _0012_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_2641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_top_iw_I\[15\].genblk1.cell0_I net500 net437 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0984_ col\[0\].genblk1.mux4_I\[13\].x _0204_ vssd1 vssd1 vccd1 vccd1 bus_ow\[13\]
+ sky130_fd_sc_hd__ebufn_8
Xcol\[4\].genblk1.mux4_I\[22\].cell0_I net162 net188 net215 net241 net471 net458 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[22\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_2_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0418_ _0042_ _0044_ _0066_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__or3_1
X_0349_ _0031_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_2346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_2493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[6\].zbuf_top_iw_I\[5\].genblk1.cell0_I net486 net442 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_2390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0967_ bus_ow\[20\] _0187_ vssd1 vssd1 vccd1 vccd1 spine_ow[21] sky130_fd_sc_hd__ebufn_8
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0898_ col\[3\].zbuf_top_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[7] sky130_fd_sc_hd__buf_2
XFILLER_0_3_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_2029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout492 col\[0\].zbuf_bot_iw_I\[2\].a vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__clkbuf_4
Xfanout481 col\[0\].zbuf_bot_iw_I\[7\].a vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__buf_6
Xfanout470 net471 vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__buf_4
XFILLER_0_13_2841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0821_ col\[6\].zbuf_bot_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[218] sky130_fd_sc_hd__buf_2
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0752_ col\[4\].zbuf_bot_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[149] sky130_fd_sc_hd__buf_2
XFILLER_0_4_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0683_ col\[2\].zbuf_bot_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[80] sky130_fd_sc_hd__buf_2
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_2205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_2115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1020_ col\[4\].genblk1.mux4_I\[1\].x _0240_ vssd1 vssd1 vccd1 vccd1 bus_ow\[1\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_2903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xzbuf_bus_ena_I.genblk1.cell0_I net16 net516 vssd1 vssd1 vccd1 vccd1 zbuf_bus_ena_I.genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0804_ col\[5\].zbuf_top_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[201] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0735_ col\[3\].zbuf_top_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[132] sky130_fd_sc_hd__buf_2
X_0666_ col\[1\].zbuf_top_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[63] sky130_fd_sc_hd__buf_2
XFILLER_0_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0597_ _0161_ vssd1 vssd1 vccd1 vccd1 col\[5\].zbuf_top_ena_I.e sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_2402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput302 um_ow[340] vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput324 um_ow[360] vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput335 um_ow[370] vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__clkbuf_2
Xinput313 um_ow[350] vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput346 um_ow[380] vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__clkbuf_2
Xinput357 um_ow[44] vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__clkbuf_2
Xinput379 um_ow[64] vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__clkbuf_1
Xinput368 um_ow[54] vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_2013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_6 col\[0\].zbuf_bot_iw_I\[16\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0520_ _0124_ _0121_ _0122_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__or3b_1
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0451_ _0090_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__clkbuf_1
X_0382_ _0043_ _0045_ _0047_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__or3_1
Xcol\[0\].zbuf_top_iw_I\[16\].genblk1.cell0_I net497 net435 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1003_ col\[2\].genblk1.mux4_I\[8\].x _0223_ vssd1 vssd1 vccd1 vccd1 bus_ow\[8\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_11_1929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0718_ col\[3\].zbuf_bot_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[115] sky130_fd_sc_hd__buf_2
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0649_ col\[1\].zbuf_bot_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[46] sky130_fd_sc_hd__buf_2
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[3\].zbuf_bot_ena_I.genblk1.cell0_I net542 net428 vssd1 vssd1 vccd1 vccd1 col\[3\].zbuf_bot_ena_I.z
+ sky130_fd_sc_hd__and2_1
XFILLER_0_7_2377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput110 um_ow[168] vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_1
Xinput121 um_ow[178] vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_1
Xinput132 um_ow[188] vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_1
Xinput143 um_ow[198] vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_1
Xinput154 um_ow[207] vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__clkbuf_1
Xinput165 um_ow[217] vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_1
Xinput176 um_ow[227] vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_1
Xinput187 um_ow[237] vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_1
Xinput198 um_ow[247] vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_15_2029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.mux4_I\[16\].cell0_I net49 net75 net102 net128 net467 net456 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[16\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_10_2641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_2685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[1\].zbuf_bot_iw_I\[0\].genblk1.cell0_I net511 net434 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_bot_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0503_ _0111_ _0108_ _0109_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__or3b_1
XFILLER_0_10_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0434_ _0080_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__clkbuf_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0365_ _0039_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_2653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_2517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[14\].genblk1.cell1_I zbuf_bus_iw_I\[14\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[14\].a sky130_fd_sc_hd__buf_6
XFILLER_0_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[2\].zbuf_top_iw_I\[15\].genblk1.cell0_I net499 net429 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0983_ col\[0\].genblk1.mux4_I\[12\].x _0203_ vssd1 vssd1 vccd1 vccd1 bus_ow\[12\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_2460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0417_ _0070_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__clkbuf_1
X_0348_ _0023_ _0024_ _0025_ _0026_ vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_2314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[6\].zbuf_bot_iw_I\[17\].genblk1.cell0_I net496 net450 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_bot_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xzbuf_bus_iw_I\[1\].genblk1.cell1_I zbuf_bus_iw_I\[1\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[1\].a sky130_fd_sc_hd__buf_6
XFILLER_0_12_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].zbuf_bot_iw_I\[8\].genblk1.cell0_I net479 net446 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_bot_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_2601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_2380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_bot_iw_I\[3\].genblk1.cell0_I net489 net444 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_bot_iw_I\[3\].z sky130_fd_sc_hd__and2_1
X_0966_ bus_ow\[19\] _0186_ vssd1 vssd1 vccd1 vccd1 spine_ow[20] sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[4\].zbuf_top_iw_I\[14\].genblk1.cell0_I net501 net423 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0897_ col\[3\].zbuf_bot_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[6] sky130_fd_sc_hd__buf_2
XFILLER_0_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout482 col\[0\].zbuf_bot_iw_I\[7\].a vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__clkbuf_4
Xfanout493 col\[0\].zbuf_bot_iw_I\[1\].a vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__buf_6
Xfanout471 net472 vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__buf_4
Xfanout460 net461 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_2
XFILLER_0_9_2055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_top_iw_I\[7\].genblk1.cell0_I net481 net436 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_2564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0820_ col\[6\].zbuf_bot_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[217] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0751_ col\[4\].zbuf_bot_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[148] sky130_fd_sc_hd__buf_2
XFILLER_0_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0682_ col\[2\].zbuf_bot_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[79] sky130_fd_sc_hd__buf_2
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[2\].zbuf_top_iw_I\[2\].genblk1.cell0_I net491 net430 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[7\].zbuf_top_ena_I.genblk1.cell0_I net551 net438 vssd1 vssd1 vccd1 vccd1 col\[7\].zbuf_top_ena_I.z
+ sky130_fd_sc_hd__and2_1
XFILLER_0_12_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0949_ bus_ow\[2\] _0169_ vssd1 vssd1 vccd1 vccd1 spine_ow[3] sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[6\].zbuf_top_iw_I\[13\].genblk1.cell0_I net504 net441 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0803_ col\[5\].zbuf_top_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[200] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0734_ col\[3\].zbuf_top_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[131] sky130_fd_sc_hd__buf_2
XFILLER_0_13_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xzbuf_bus_iw_I\[10\].genblk1.cell0_I net19 net515 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[10\].genblk1.l
+ sky130_fd_sc_hd__and2_1
X_0665_ col\[1\].zbuf_top_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[62] sky130_fd_sc_hd__buf_2
X_0596_ _0147_ _0148_ net463 _0158_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_2414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[7\].zbuf_bot_iw_I\[6\].genblk1.cell0_I net484 net440 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_bot_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_2136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_2169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput303 um_ow[341] vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput336 um_ow[371] vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput325 um_ow[361] vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput314 um_ow[351] vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput347 um_ow[381] vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_2
Xinput358 um_ow[45] vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__clkbuf_2
Xinput369 um_ow[55] vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_2025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_2069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_7 col\[0\].zbuf_bot_iw_I\[16\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0450_ _0083_ _0089_ _0084_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__or3b_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0381_ _0050_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__clkbuf_1
X_1002_ col\[2\].genblk1.mux4_I\[7\].x _0222_ vssd1 vssd1 vccd1 vccd1 bus_ow\[7\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_8_2879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0717_ col\[3\].zbuf_bot_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[114] sky130_fd_sc_hd__buf_2
XFILLER_0_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0648_ col\[1\].zbuf_bot_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[45] sky130_fd_sc_hd__buf_2
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0579_ _0151_ vssd1 vssd1 vccd1 vccd1 col\[1\].zbuf_top_ena_I.e sky130_fd_sc_hd__clkbuf_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_2200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[5\].zbuf_top_iw_I\[5\].genblk1.cell0_I net486 net420 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput111 um_ow[169] vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_1
Xinput100 um_ow[159] vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_1
Xinput122 um_ow[179] vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__clkbuf_1
Xinput133 um_ow[189] vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_1
Xinput144 um_ow[199] vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_1
Xinput166 um_ow[218] vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_1
Xinput177 um_ow[228] vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_1
Xinput155 um_ow[208] vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__clkbuf_1
Xcol\[7\].zbuf_top_iw_I\[0\].genblk1.cell0_I net512 net438 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[0\].z sky130_fd_sc_hd__and2_1
Xinput188 um_ow[238] vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_1
Xinput199 um_ow[248] vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__dlymetal6s2s_1
Xcol\[0\].genblk1.mux4_I\[21\].cell0_I net168 net358 net384 net411 net464 net451 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[21\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_6_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0502_ _0118_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0433_ _0075_ _0076_ _0077_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__or3b_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0364_ _0001_ _0005_ _0008_ _0012_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_2529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_2687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_2417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_2597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_2253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_2017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0982_ col\[0\].genblk1.mux4_I\[11\].x _0202_ vssd1 vssd1 vccd1 vccd1 bus_ow\[11\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_3_2573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0416_ _0058_ _0059_ _0066_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__or3_1
X_0347_ _0030_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_2372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[1\].zbuf_bot_iw_I\[17\].genblk1.cell0_I net495 net433 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_bot_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_2061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_2781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_2578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0965_ bus_ow\[18\] _0185_ vssd1 vssd1 vccd1 vccd1 spine_ow[19] sky130_fd_sc_hd__ebufn_8
XFILLER_0_12_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0896_ col\[2\].zbuf_top_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[5] sky130_fd_sc_hd__buf_2
XFILLER_0_3_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtt_mux_530 vssd1 vssd1 vccd1 vccd1 tt_mux_530/HI um_k_zero[10] sky130_fd_sc_hd__conb_1
XFILLER_0_13_2309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtt_mux_552 vssd1 vssd1 vccd1 vccd1 k_one tt_mux_552/LO sky130_fd_sc_hd__conb_1
XFILLER_0_6_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout450 col\[6\].zbuf_bot_ena_I.e vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__clkbuf_2
Xfanout483 col\[0\].zbuf_bot_iw_I\[6\].a vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__buf_6
Xfanout461 net462 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__buf_2
Xfanout472 net476 vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__clkbuf_4
Xfanout494 col\[0\].zbuf_bot_iw_I\[1\].a vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_2067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0750_ col\[4\].zbuf_bot_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[147] sky130_fd_sc_hd__buf_2
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0681_ col\[2\].zbuf_bot_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[78] sky130_fd_sc_hd__buf_2
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[3\].zbuf_bot_iw_I\[16\].genblk1.cell0_I net497 net427 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_bot_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_2432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0948_ bus_ow\[1\] _0168_ vssd1 vssd1 vccd1 vccd1 spine_ow[2] sky130_fd_sc_hd__ebufn_8
X_0879_ col\[7\].zbuf_top_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[276] sky130_fd_sc_hd__buf_2
XFILLER_0_2_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].zbuf_bot_iw_I\[0\].genblk1.cell0_I net511 net448 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_bot_iw_I\[0\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_iw_I\[13\].genblk1.cell0_I net503 net431 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_2763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_sel_I\[3\].genblk1.cell1_I zbuf_bus_sel_I\[3\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 zbuf_bus_sel_I\[3\].z sky130_fd_sc_hd__buf_8
XFILLER_0_13_1961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0802_ col\[5\].zbuf_top_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[199] sky130_fd_sc_hd__buf_2
XFILLER_0_13_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0733_ col\[3\].zbuf_top_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[130] sky130_fd_sc_hd__buf_2
X_0664_ col\[1\].zbuf_top_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[61] sky130_fd_sc_hd__buf_2
XFILLER_0_0_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0595_ _0160_ vssd1 vssd1 vccd1 vccd1 col\[5\].zbuf_bot_ena_I.e sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput326 um_ow[362] vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput315 um_ow[352] vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput304 um_ow[342] vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput359 um_ow[46] vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__clkbuf_2
Xinput337 um_ow[372] vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__clkbuf_2
Xinput348 um_ow[382] vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__dlymetal6s2s_1
Xcol\[5\].zbuf_bot_iw_I\[15\].genblk1.cell0_I net500 net421 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_bot_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_2903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_8 col\[0\].zbuf_bot_iw_I\[17\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0380_ _0043_ _0045_ _0047_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__or3_1
X_1001_ col\[2\].genblk1.mux4_I\[6\].x _0221_ vssd1 vssd1 vccd1 vccd1 bus_ow\[6\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_2757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_2468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0716_ col\[3\].zbuf_bot_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[113] sky130_fd_sc_hd__buf_2
XFILLER_0_0_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0647_ col\[1\].zbuf_bot_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[44] sky130_fd_sc_hd__buf_2
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0578_ _0147_ _0148_ _0145_ _0146_ vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__and4_2
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[3\].zbuf_top_iw_I\[12\].genblk1.cell0_I net505 net425 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_2267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[1\].zbuf_bot_iw_I\[8\].genblk1.cell0_I net479 net433 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_bot_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput101 um_ow[15] vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput112 um_ow[16] vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput145 um_ow[19] vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput134 um_ow[18] vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput123 um_ow[17] vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput167 um_ow[219] vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_1
Xinput178 um_ow[229] vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_1
Xinput156 um_ow[209] vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_1
Xinput189 um_ow[239] vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_2880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[3\].zbuf_bot_iw_I\[3\].genblk1.cell0_I net489 net428 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_bot_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_2490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0501_ _0111_ _0108_ _0109_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__or3b_1
XTAP_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0432_ _0079_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__clkbuf_1
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0363_ _0038_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_2543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_2390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[7\].zbuf_bot_iw_I\[14\].genblk1.cell0_I net502 net439 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_bot_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_11_1717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_2165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[5\].zbuf_top_iw_I\[11\].genblk1.cell0_I net508 net419 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[11\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_iw_I\[2\].genblk1.cell0_I net491 net432 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_15_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0981_ col\[0\].genblk1.mux4_I\[10\].x _0201_ vssd1 vssd1 vccd1 vccd1 bus_ow\[10\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_3_1840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0415_ _0069_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__clkbuf_1
X_0346_ _0023_ _0024_ _0025_ _0026_ vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__or4_1
Xzbuf_bus_iw_I\[9\].genblk1.cell1_I zbuf_bus_iw_I\[9\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[9\].a sky130_fd_sc_hd__buf_6
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[6\].zbuf_bot_iw_I\[6\].genblk1.cell0_I net484 net449 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_bot_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_2625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_2647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0964_ bus_ow\[17\] _0184_ vssd1 vssd1 vccd1 vccd1 spine_ow[18] sky130_fd_sc_hd__ebufn_8
XFILLER_0_3_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_2281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0895_ col\[2\].zbuf_bot_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[4] sky130_fd_sc_hd__buf_2
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0329_ _0019_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__clkbuf_1
Xtt_mux_531 vssd1 vssd1 vccd1 vccd1 tt_mux_531/HI um_k_zero[11] sky130_fd_sc_hd__conb_1
Xtt_mux_520 vssd1 vssd1 vccd1 vccd1 tt_mux_520/HI um_k_zero[0] sky130_fd_sc_hd__conb_1
XFILLER_0_4_2113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_2181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[7\].zbuf_top_iw_I\[10\].genblk1.cell0_I net510 net437 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout440 col\[7\].zbuf_bot_ena_I.e vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout484 col\[0\].zbuf_bot_iw_I\[6\].a vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__clkbuf_4
Xcol\[4\].genblk1.mux4_I\[12\].cell0_I net151 net177 net204 net230 net471 net458 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[12\].x sky130_fd_sc_hd__mux4_1
Xfanout451 net453 vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__clkbuf_4
Xfanout473 net474 vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__clkbuf_4
Xfanout462 net463 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__buf_2
Xfanout495 col\[0\].zbuf_bot_iw_I\[17\].a vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_6
XFILLER_0_9_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0680_ col\[2\].zbuf_bot_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[77] sky130_fd_sc_hd__buf_2
XFILLER_0_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[4\].zbuf_top_iw_I\[5\].genblk1.cell0_I net485 net424 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_2477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0947_ bus_ow\[0\] _0167_ vssd1 vssd1 vccd1 vccd1 spine_ow[1] sky130_fd_sc_hd__ebufn_8
XFILLER_0_3_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0878_ col\[7\].zbuf_top_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[275] sky130_fd_sc_hd__buf_2
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].zbuf_top_iw_I\[0\].genblk1.cell0_I net512 net442 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_2107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_2129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.mux4_I\[22\].cell0_I net269 net295 net321 net348 net475 net462 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[22\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_13_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0801_ col\[5\].zbuf_top_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[198] sky130_fd_sc_hd__buf_2
XFILLER_0_13_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0732_ col\[3\].zbuf_top_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[129] sky130_fd_sc_hd__buf_2
X_0663_ col\[1\].zbuf_top_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[60] sky130_fd_sc_hd__buf_2
X_0594_ _0147_ _0148_ _0145_ _0158_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__and4b_1
XFILLER_0_0_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].zbuf_bot_iw_I\[15\].genblk1.cell0_I net499 net447 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_bot_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput327 um_ow[363] vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput316 um_ow[353] vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput305 um_ow[343] vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput338 um_ow[373] vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_2
Xinput349 um_ow[383] vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_6_1326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_2836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_9 col\[0\].zbuf_bot_iw_I\[17\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_2804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1000_ col\[2\].genblk1.mux4_I\[5\].x _0220_ vssd1 vssd1 vccd1 vccd1 bus_ow\[5\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_8_2826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_2561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[5\].genblk1.cell0_I net13 net514 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[5\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_2_1724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0715_ col\[3\].zbuf_bot_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[112] sky130_fd_sc_hd__buf_2
XFILLER_0_0_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0646_ col\[1\].zbuf_bot_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[43] sky130_fd_sc_hd__buf_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0577_ _0150_ vssd1 vssd1 vccd1 vccd1 col\[1\].zbuf_bot_ena_I.e sky130_fd_sc_hd__clkbuf_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[7\].zbuf_top_iw_I\[8\].genblk1.cell0_I net480 net438 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput102 um_ow[160] vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_1
Xinput113 um_ow[170] vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__clkbuf_1
Xinput135 um_ow[190] vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__clkbuf_1
Xinput124 um_ow[180] vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__clkbuf_1
Xinput146 um_ow[1] vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__clkbuf_2
Xinput157 um_ow[20] vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput168 um_ow[21] vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput179 um_ow[22] vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_2712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0500_ _0117_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__clkbuf_1
XTAP_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0431_ _0075_ _0076_ _0077_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__or3b_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0362_ _0001_ _0005_ _0008_ _0012_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__or4_1
Xcol\[2\].zbuf_bot_iw_I\[14\].genblk1.cell0_I net501 net445 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_bot_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_15_2500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_2511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_2907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[0\].zbuf_top_iw_I\[11\].genblk1.cell0_I net507 net435 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_12_2717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0980_ col\[0\].genblk1.mux4_I\[9\].x _0200_ vssd1 vssd1 vccd1 vccd1 bus_ow\[9\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_3_1885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0414_ _0058_ _0059_ _0066_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__or3_1
X_0345_ _0029_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_2330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[4\].zbuf_bot_iw_I\[13\].genblk1.cell0_I net503 net443 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_bot_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_2547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0963_ bus_ow\[16\] _0183_ vssd1 vssd1 vccd1 vccd1 spine_ow[17] sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0894_ col\[1\].zbuf_top_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[3] sky130_fd_sc_hd__buf_2
XFILLER_0_10_2293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0328_ _0002_ _0006_ _0009_ _0013_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__or4_1
Xtt_mux_521 vssd1 vssd1 vccd1 vccd1 tt_mux_521/HI um_k_zero[1] sky130_fd_sc_hd__conb_1
Xtt_mux_532 vssd1 vssd1 vccd1 vccd1 tt_mux_532/HI um_k_zero[12] sky130_fd_sc_hd__conb_1
Xcol\[2\].zbuf_top_iw_I\[10\].genblk1.cell0_I net509 net429 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_2125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout441 col\[6\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__clkbuf_2
Xfanout430 col\[2\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout452 net453 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__buf_2
Xfanout474 net475 vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__clkbuf_4
Xfanout463 zbuf_bus_sel_I\[1\].z vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_6
Xfanout485 col\[0\].zbuf_bot_iw_I\[5\].a vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_6
Xfanout496 col\[0\].zbuf_bot_iw_I\[17\].a vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[16\].cell0_I net155 net182 net208 net235 net470 net457 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[16\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_6_2924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_2670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_2556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_2401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_2489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_bot_iw_I\[8\].genblk1.cell0_I net479 net447 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_bot_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0946_ col\[1\].zbuf_bot_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[39] sky130_fd_sc_hd__buf_2
Xcol\[6\].zbuf_bot_iw_I\[12\].genblk1.cell0_I net506 net450 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_bot_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0877_ col\[7\].zbuf_top_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[274] sky130_fd_sc_hd__buf_2
XFILLER_0_3_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].zbuf_bot_iw_I\[3\].genblk1.cell0_I net489 net446 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_bot_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0800_ col\[5\].zbuf_bot_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[197] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0731_ col\[3\].zbuf_top_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[128] sky130_fd_sc_hd__buf_2
XFILLER_0_13_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0662_ col\[1\].zbuf_top_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[59] sky130_fd_sc_hd__buf_2
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0593_ _0159_ vssd1 vssd1 vccd1 vccd1 col\[4\].zbuf_top_ena_I.e sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_2264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0929_ col\[0\].zbuf_top_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[22] sky130_fd_sc_hd__buf_2
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput306 um_ow[344] vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput317 um_ow[354] vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput328 um_ow[364] vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput339 um_ow[374] vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__dlymetal6s2s_1
Xcol\[0\].zbuf_top_iw_I\[2\].genblk1.cell0_I net491 net436 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_1338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_2816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_2849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_2472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0714_ col\[3\].zbuf_bot_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[111] sky130_fd_sc_hd__buf_2
X_0645_ col\[1\].zbuf_bot_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[42] sky130_fd_sc_hd__buf_2
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0576_ _0147_ _0148_ _0145_ _0146_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__and4b_2
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_2225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1059_ col\[6\].genblk1.mux4_I\[16\].x _0279_ vssd1 vssd1 vccd1 vccd1 bus_ow\[16\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_5_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[3\].zbuf_top_ena_I.genblk1.cell0_I net543 net425 vssd1 vssd1 vccd1 vccd1 col\[3\].zbuf_top_ena_I.z
+ sky130_fd_sc_hd__and2_1
XFILLER_0_4_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput114 um_ow[171] vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkbuf_1
Xinput125 um_ow[181] vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_1
Xinput136 um_ow[191] vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_1
Xinput103 um_ow[161] vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_1
Xinput169 um_ow[220] vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_1
Xinput147 um_ow[200] vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_1
Xinput158 um_ow[210] vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__clkbuf_1
Xcol\[5\].zbuf_bot_iw_I\[6\].genblk1.cell0_I net484 net422 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_bot_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_2757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_2601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_2481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0430_ _0078_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__clkbuf_1
X_0361_ _0037_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__clkbuf_1
Xcol\[7\].zbuf_bot_iw_I\[1\].genblk1.cell0_I net494 net440 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_bot_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_1901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0559_ _0001_ _0005_ _0008_ _0012_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__or4_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_2009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_top_ena_I.genblk1.cell0_I_537 vssd1 vssd1 vccd1 vccd1 net537 col\[0\].zbuf_top_ena_I.genblk1.cell0_I_537/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_9_2911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[3\].zbuf_top_iw_I\[5\].genblk1.cell0_I net485 net426 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_2808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0413_ _0068_ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__clkbuf_1
Xcol\[5\].zbuf_top_iw_I\[0\].genblk1.cell0_I net512 net420 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[0\].z sky130_fd_sc_hd__and2_1
X_0344_ _0023_ _0024_ _0025_ _0026_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_2443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].genblk1.mux4_I\[11\].cell0_I net57 net323 net373 net400 net465 net452 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[11\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_1_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_2896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_2740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_2351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_2537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0962_ bus_ow\[15\] _0182_ vssd1 vssd1 vccd1 vccd1 spine_ow[16] sky130_fd_sc_hd__ebufn_8
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0893_ col\[1\].zbuf_bot_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[2] sky130_fd_sc_hd__buf_2
XFILLER_0_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0327_ _0018_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__clkbuf_1
Xtt_mux_522 vssd1 vssd1 vccd1 vccd1 tt_mux_522/HI um_k_zero[2] sky130_fd_sc_hd__conb_1
Xtt_mux_533 vssd1 vssd1 vccd1 vccd1 tt_mux_533/HI um_k_zero[13] sky130_fd_sc_hd__conb_1
XFILLER_0_8_2262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_2137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout431 col\[1\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__clkbuf_2
Xfanout420 col\[5\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__dlymetal6s2s_1
Xcol\[2\].genblk1.mux4_I\[21\].cell0_I net54 net81 net107 net133 net467 net456 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[21\].x sky130_fd_sc_hd__mux4_1
Xfanout442 col\[6\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout464 net466 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__buf_4
Xfanout453 net463 vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__buf_2
Xfanout475 net476 vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__clkbuf_4
Xfanout486 col\[0\].zbuf_bot_iw_I\[5\].a vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__clkbuf_4
Xfanout497 col\[0\].zbuf_bot_iw_I\[16\].a vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__buf_6
XFILLER_0_9_2015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_2037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].zbuf_top_iw_I\[8\].genblk1.cell0_I net480 net442 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[8\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_ena_I.genblk1.cell0_I_539 vssd1 vssd1 vccd1 vccd1 net539 col\[1\].zbuf_top_ena_I.genblk1.cell0_I_539/LO
+ sky130_fd_sc_hd__conb_1
Xcol\[1\].zbuf_bot_iw_I\[12\].genblk1.cell0_I net505 net433 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_bot_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_2457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_2323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0945_ col\[1\].zbuf_bot_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[38] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0876_ col\[7\].zbuf_top_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[273] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0730_ col\[3\].zbuf_top_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[127] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0661_ col\[1\].zbuf_top_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[58] sky130_fd_sc_hd__buf_2
X_0592_ _0145_ _0158_ net472 zbuf_bus_ena_I.z vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__and4b_1
XFILLER_0_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_2221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0928_ col\[0\].zbuf_top_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[21] sky130_fd_sc_hd__buf_2
X_0859_ col\[7\].zbuf_bot_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[256] sky130_fd_sc_hd__buf_2
XFILLER_0_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput318 um_ow[355] vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput307 um_ow[345] vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput329 um_ow[365] vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_6_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[3\].zbuf_bot_iw_I\[11\].genblk1.cell0_I net507 net427 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_bot_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_2541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_2427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0713_ col\[3\].zbuf_bot_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[110] sky130_fd_sc_hd__buf_2
X_0644_ col\[1\].zbuf_bot_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[41] sky130_fd_sc_hd__buf_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0575_ _0149_ vssd1 vssd1 vccd1 vccd1 col\[0\].zbuf_top_ena_I.e sky130_fd_sc_hd__clkbuf_2
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_2237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1058_ col\[6\].genblk1.mux4_I\[15\].x _0278_ vssd1 vssd1 vccd1 vccd1 bus_ow\[15\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_5_2073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput115 um_ow[172] vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__clkbuf_1
Xinput126 um_ow[182] vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_1
Xinput104 um_ow[162] vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_1
Xinput148 um_ow[201] vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__clkbuf_1
Xinput159 um_ow[211] vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__clkbuf_1
Xinput137 um_ow[192] vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_2850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_2861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_2872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0360_ _0001_ _0005_ _0008_ _0012_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_2603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[5\].zbuf_bot_iw_I\[10\].genblk1.cell0_I net510 net421 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_bot_iw_I\[10\].z sky130_fd_sc_hd__and2_1
X_0558_ _0075_ _0077_ _0047_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__nand3b_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0489_ _0111_ _0108_ _0109_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__or3b_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_2001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0412_ _0058_ _0059_ _0066_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__or3_1
X_0343_ _0028_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_2455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[1\].zbuf_bot_iw_I\[3\].genblk1.cell0_I net489 net434 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_bot_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_1765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[0\].genblk1.mux4_I\[15\].cell0_I net101 net351 net378 net404 net464 net451 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[15\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_1_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_2717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[17\].genblk1.cell1_I zbuf_bus_iw_I\[17\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[17\].a sky130_fd_sc_hd__buf_6
XFILLER_0_11_2730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_2786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0961_ bus_ow\[14\] _0181_ vssd1 vssd1 vccd1 vccd1 spine_ow[15] sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0892_ col\[0\].zbuf_top_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[1] sky130_fd_sc_hd__buf_2
X_0326_ _0002_ _0006_ _0009_ _0013_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__or4_1
Xtt_mux_523 vssd1 vssd1 vccd1 vccd1 tt_mux_523/HI um_k_zero[3] sky130_fd_sc_hd__conb_1
Xtt_mux_534 vssd1 vssd1 vccd1 vccd1 tt_mux_534/HI um_k_zero[14] sky130_fd_sc_hd__conb_1
XFILLER_0_4_2149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout432 col\[1\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout421 col\[5\].zbuf_bot_ena_I.e vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__clkbuf_2
Xfanout443 col\[4\].zbuf_bot_ena_I.e vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__clkbuf_2
Xfanout465 net466 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__clkbuf_4
Xfanout454 net455 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__clkbuf_4
Xfanout487 col\[0\].zbuf_bot_iw_I\[4\].a vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__buf_6
Xfanout498 col\[0\].zbuf_bot_iw_I\[16\].a vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__clkbuf_4
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout476 zbuf_bus_sel_I\[0\].z vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__buf_8
XFILLER_0_6_2915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_2825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_2683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.mux4_I\[2\].cell0_I net246 net273 net299 net326 net473 net460 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[2\].x sky130_fd_sc_hd__mux4_1
Xzbuf_bus_iw_I\[4\].genblk1.cell1_I zbuf_bus_iw_I\[4\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[4\].a sky130_fd_sc_hd__buf_6
XFILLER_0_5_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_2379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0944_ col\[1\].zbuf_bot_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[37] sky130_fd_sc_hd__buf_2
XFILLER_0_10_2070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0875_ col\[7\].zbuf_top_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[272] sky130_fd_sc_hd__buf_2
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[4\].zbuf_bot_iw_I\[6\].genblk1.cell0_I net483 net444 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_bot_iw_I\[6\].z sky130_fd_sc_hd__and2_1
X_0309_ _0005_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_8_2071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_top_iw_I\[17\].genblk1.cell0_I net495 net423 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.mux4_I\[0\].cell0_I net414 net58 net84 net110 net468 net454 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[0\].x sky130_fd_sc_hd__mux4_1
Xcol\[6\].zbuf_bot_iw_I\[1\].genblk1.cell0_I net494 net449 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_bot_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_2633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_2390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0660_ col\[1\].zbuf_top_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[57] sky130_fd_sc_hd__buf_2
X_0591_ _0240_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0927_ col\[0\].zbuf_top_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[20] sky130_fd_sc_hd__buf_2
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0858_ col\[7\].zbuf_bot_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[255] sky130_fd_sc_hd__buf_2
XFILLER_0_3_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0789_ col\[5\].zbuf_bot_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[186] sky130_fd_sc_hd__buf_2
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput308 um_ow[346] vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput319 um_ow[356] vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__dlymetal6s2s_1
Xcol\[2\].zbuf_top_iw_I\[5\].genblk1.cell0_I net485 net430 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_2620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[4\].zbuf_top_iw_I\[0\].genblk1.cell0_I net511 net424 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_2163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0712_ col\[3\].zbuf_bot_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[109] sky130_fd_sc_hd__buf_2
X_0643_ col\[1\].zbuf_bot_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[40] sky130_fd_sc_hd__buf_2
XFILLER_0_0_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].zbuf_top_iw_I\[16\].genblk1.cell0_I net498 net441 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0574_ _0145_ _0146_ _0147_ _0148_ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__and4b_2
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1057_ col\[6\].genblk1.mux4_I\[14\].x _0277_ vssd1 vssd1 vccd1 vccd1 bus_ow\[14\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_5_2085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[13\].genblk1.cell0_I net22 net515 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[13\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_1_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[6\].genblk1.mux4_I\[12\].cell0_I net258 net284 net310 net337 net474 net461 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[12\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_11_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput127 um_ow[183] vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_1
Xinput116 um_ow[173] vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_1
Xinput105 um_ow[163] vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_1
Xcol\[7\].zbuf_bot_iw_I\[9\].genblk1.cell0_I net478 net439 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_bot_iw_I\[9\].z sky130_fd_sc_hd__and2_1
Xinput149 um_ow[202] vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_1
Xinput138 um_ow[193] vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_2737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_2472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_2659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[0\].zbuf_bot_iw_I\[10\].genblk1.cell0_I net509 net447 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_bot_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_1581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0557_ _0075_ _0077_ _0047_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__nand3b_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[4\].genblk1.mux4_I\[3\].cell0_I net140 net167 net194 net220 net472 net459 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[3\].x sky130_fd_sc_hd__mux4_1
X_0488_ _0042_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__clkbuf_2
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[5\].zbuf_top_iw_I\[8\].genblk1.cell0_I net480 net419 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xzbuf_bus_iw_I\[0\].genblk1.cell0_I net8 net513 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[0\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_9_2924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_top_iw_I\[3\].genblk1.cell0_I net490 net438 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[3\].z sky130_fd_sc_hd__and2_1
X_0411_ _0067_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__clkbuf_1
X_0342_ _0023_ _0024_ _0025_ _0026_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_2412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[0\].genblk1.mux4_I\[1\].cell0_I net146 net212 net362 net389 net466 net453 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[1\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_8_2434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[0\].genblk1.mux4_I\[19\].cell0_I net145 net356 net382 net409 net464 net451 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[19\].x sky130_fd_sc_hd__mux4_2
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_2798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0960_ bus_ow\[13\] _0180_ vssd1 vssd1 vccd1 vccd1 spine_ow[14] sky130_fd_sc_hd__ebufn_8
XFILLER_0_7_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0891_ col\[0\].zbuf_bot_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[0] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0325_ _0017_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__clkbuf_1
Xtt_mux_535 vssd1 vssd1 vccd1 vccd1 tt_mux_535/HI um_k_zero[15] sky130_fd_sc_hd__conb_1
Xtt_mux_524 vssd1 vssd1 vccd1 vccd1 tt_mux_524/HI um_k_zero[4] sky130_fd_sc_hd__conb_1
XFILLER_0_8_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout422 col\[5\].zbuf_bot_ena_I.e vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_10_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout433 col\[1\].zbuf_bot_ena_I.e vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__clkbuf_2
Xfanout444 col\[4\].zbuf_bot_ena_I.e vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout455 net463 vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__clkbuf_2
Xfanout466 net476 vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__buf_4
Xfanout488 col\[0\].zbuf_bot_iw_I\[4\].a vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__clkbuf_4
Xfanout477 col\[0\].zbuf_bot_iw_I\[9\].a vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__buf_6
Xfanout499 col\[0\].zbuf_bot_iw_I\[15\].a vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__buf_6
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].genblk1.mux4_I\[6\].cell0_I net250 net277 net304 net330 net473 net460 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[6\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_9_1861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0943_ col\[1\].zbuf_bot_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[36] sky130_fd_sc_hd__buf_2
XFILLER_0_3_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0874_ col\[7\].zbuf_top_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[271] sky130_fd_sc_hd__buf_2
XFILLER_0_10_2082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0308_ _0003_ net34 net1 _0004_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__a22o_2
XFILLER_0_4_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_2083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[2\].genblk1.mux4_I\[4\].cell0_I net36 net62 net88 net115 net468 net454 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[4\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_13_2601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0590_ _0157_ vssd1 vssd1 vccd1 vccd1 col\[4\].zbuf_bot_ena_I.e sky130_fd_sc_hd__inv_2
XFILLER_0_5_2289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0926_ col\[0\].zbuf_top_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[19] sky130_fd_sc_hd__buf_2
XFILLER_0_7_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0857_ col\[7\].zbuf_bot_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[254] sky130_fd_sc_hd__buf_2
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0788_ col\[5\].zbuf_bot_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[185] sky130_fd_sc_hd__buf_2
Xinput309 um_ow[347] vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_10_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[1\].zbuf_top_iw_I\[16\].genblk1.cell0_I net497 net431 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[16\].z sky130_fd_sc_hd__and2_1
Xcol\[0\].zbuf_bot_iw_I\[3\].genblk1.cell0_I net489 net448 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_bot_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0711_ col\[3\].zbuf_bot_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[108] sky130_fd_sc_hd__buf_2
XFILLER_0_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0573_ zbuf_bus_ena_I.z vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__buf_4
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1056_ col\[6\].genblk1.mux4_I\[13\].x _0276_ vssd1 vssd1 vccd1 vccd1 bus_ow\[13\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_5_2053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_2097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0909_ col\[0\].zbuf_bot_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[2] sky130_fd_sc_hd__buf_2
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput117 um_ow[174] vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_1
Xinput106 um_ow[164] vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_1
Xinput128 um_ow[184] vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__clkbuf_1
Xinput139 um_ow[194] vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__clkbuf_1
Xcol\[6\].genblk1.mux4_I\[16\].cell0_I net262 net288 net315 net341 net474 net461 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[16\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_14_2740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_90 spine_iw[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_2605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0556_ _0137_ _0138_ _0139_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__nand3b_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0487_ _0110_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__clkbuf_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[7\].cell0_I net144 net172 net198 net225 net470 net457 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[7\].x sky130_fd_sc_hd__mux4_1
X_1039_ col\[4\].genblk1.mux4_I\[20\].x _0259_ vssd1 vssd1 vccd1 vccd1 bus_ow\[20\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_7_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[3\].zbuf_top_iw_I\[15\].genblk1.cell0_I net499 net425 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0410_ _0058_ _0059_ _0066_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__or3_1
X_0341_ _0027_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__clkbuf_1
Xcol\[3\].zbuf_bot_iw_I\[6\].genblk1.cell0_I net483 net428 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_bot_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_1745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[0\].genblk1.mux4_I\[5\].cell0_I net374 net256 net367 net393 net466 net453 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[5\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_6_2181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0539_ _0134_ _0135_ _0136_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__nand3b_2
Xcol\[5\].zbuf_bot_iw_I\[1\].genblk1.cell0_I net494 net422 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_bot_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[7\].zbuf_bot_iw_I\[17\].genblk1.cell0_I net496 net439 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_bot_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_2822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_2710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0890_ col\[7\].zbuf_top_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[287] sky130_fd_sc_hd__buf_2
XFILLER_0_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[5\].zbuf_top_iw_I\[14\].genblk1.cell0_I net502 net419 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[14\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_iw_I\[5\].genblk1.cell0_I net485 net432 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[5\].z sky130_fd_sc_hd__and2_1
X_0324_ _0002_ _0006_ _0009_ _0013_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__or4_1
Xtt_mux_525 vssd1 vssd1 vccd1 vccd1 tt_mux_525/HI um_k_zero[5] sky130_fd_sc_hd__conb_1
XFILLER_0_8_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_2017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[3\].zbuf_top_iw_I\[0\].genblk1.cell0_I net511 net426 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[0\].z sky130_fd_sc_hd__and2_1
Xfanout423 col\[4\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__clkbuf_2
Xfanout445 col\[2\].zbuf_bot_ena_I.e vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__clkbuf_2
Xfanout434 col\[1\].zbuf_bot_ena_I.e vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout456 net463 vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout478 col\[0\].zbuf_bot_iw_I\[9\].a vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__clkbuf_4
Xfanout489 col\[0\].zbuf_bot_iw_I\[3\].a vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_6
Xfanout467 net476 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_4
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_2641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xzbuf_bus_sel_I\[2\].genblk1.cell0_I net28 net516 vssd1 vssd1 vccd1 vccd1 zbuf_bus_sel_I\[2\].genblk1.l
+ sky130_fd_sc_hd__and2_2
XFILLER_0_5_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0942_ col\[0\].zbuf_top_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[35] sky130_fd_sc_hd__clkbuf_4
X_0873_ col\[7\].zbuf_top_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[270] sky130_fd_sc_hd__buf_2
XFILLER_0_10_2094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].zbuf_bot_iw_I\[9\].genblk1.cell0_I net478 net449 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_bot_iw_I\[9\].z sky130_fd_sc_hd__and2_1
X_0307_ net31 vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_2095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_2613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_top_iw_I\[13\].genblk1.cell0_I net504 net437 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_2657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].genblk1.mux4_I\[8\].cell0_I net40 net66 net93 net119 net468 net454 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[8\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_4_2493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.mux4_I\[11\].cell0_I net43 net70 net96 net122 net468 net454 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[11\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0925_ col\[0\].zbuf_top_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[18] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0856_ col\[7\].zbuf_bot_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[253] sky130_fd_sc_hd__buf_2
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0787_ col\[5\].zbuf_bot_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[184] sky130_fd_sc_hd__buf_2
Xcol\[4\].zbuf_top_iw_I\[8\].genblk1.cell0_I net479 net423 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_2933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].zbuf_top_iw_I\[3\].genblk1.cell0_I net490 net442 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_15_2708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_2432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0710_ col\[2\].zbuf_top_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[107] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0572_ net471 vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__buf_4
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1055_ col\[6\].genblk1.mux4_I\[12\].x _0275_ vssd1 vssd1 vccd1 vccd1 bus_ow\[12\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_8_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0908_ col\[0\].zbuf_bot_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[1] sky130_fd_sc_hd__buf_2
X_0839_ col\[6\].zbuf_top_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[236] sky130_fd_sc_hd__buf_2
Xcol\[4\].genblk1.mux4_I\[21\].cell0_I net161 net187 net214 net240 net471 net458 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[21\].x sky130_fd_sc_hd__mux4_1
Xinput118 um_ow[175] vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_1
Xinput107 um_ow[165] vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_1
Xinput129 um_ow[185] vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_2820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_2842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_91 net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_80 _0145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_2617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_bot_ena_I.genblk1.cell0_I net544 net444 vssd1 vssd1 vccd1 vccd1 col\[4\].zbuf_bot_ena_I.z
+ sky130_fd_sc_hd__and2_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0555_ _0137_ _0138_ _0139_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__nand3b_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0486_ _0096_ _0108_ _0109_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__or3b_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xzbuf_bus_iw_I\[8\].genblk1.cell0_I net17 net513 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[8\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1038_ col\[4\].genblk1.mux4_I\[19\].x _0258_ vssd1 vssd1 vccd1 vccd1 bus_ow\[19\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_14_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0340_ _0023_ _0024_ _0025_ _0026_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_2302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_2193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].genblk1.mux4_I\[9\].cell0_I net418 net301 net371 net398 net465 net452 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[9\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].zbuf_bot_iw_I\[17\].genblk1.cell0_I net495 net445 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_bot_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0538_ _0134_ _0135_ _0136_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__nand3b_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0469_ _0100_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__clkbuf_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_top_iw_I\[14\].genblk1.cell0_I net501 net435 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_10_1597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0323_ _0016_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__clkbuf_1
Xinput290 um_ow[32] vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_8_2211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtt_mux_526 vssd1 vssd1 vccd1 vccd1 tt_mux_526/HI um_k_zero[6] sky130_fd_sc_hd__conb_1
XFILLER_0_15_2121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_2299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout424 col\[4\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout435 net436 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout446 col\[2\].zbuf_bot_ena_I.e vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout457 net458 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_2
Xfanout479 col\[0\].zbuf_bot_iw_I\[8\].a vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__buf_6
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout468 net469 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_1827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[4\].zbuf_bot_iw_I\[16\].genblk1.cell0_I net497 net443 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_bot_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0941_ col\[0\].zbuf_top_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[34] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0872_ col\[7\].zbuf_bot_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[269] sky130_fd_sc_hd__buf_2
XFILLER_0_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0306_ net3 vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__inv_2
Xzbuf_bus_iw_I\[12\].genblk1.cell1_I zbuf_bus_iw_I\[12\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[12\].a sky130_fd_sc_hd__buf_6
XFILLER_0_8_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_2883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].zbuf_top_iw_I\[13\].genblk1.cell0_I net503 net429 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_2669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0924_ col\[0\].zbuf_bot_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[17] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0855_ col\[7\].zbuf_bot_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[252] sky130_fd_sc_hd__buf_2
Xcol\[2\].genblk1.mux4_I\[15\].cell0_I net48 net74 net100 net127 net476 net456 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[15\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_10_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0786_ col\[5\].zbuf_bot_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[183] sky130_fd_sc_hd__buf_2
XFILLER_0_3_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_2781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[6\].zbuf_bot_iw_I\[15\].genblk1.cell0_I net500 net450 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_bot_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[2\].zbuf_bot_iw_I\[6\].genblk1.cell0_I net483 net446 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_bot_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_2422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0571_ _0192_ vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__inv_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[4\].zbuf_bot_iw_I\[1\].genblk1.cell0_I net493 net444 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_bot_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_2208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1054_ col\[6\].genblk1.mux4_I\[11\].x _0274_ vssd1 vssd1 vccd1 vccd1 bus_ow\[11\]
+ sky130_fd_sc_hd__ebufn_8
Xcol\[4\].zbuf_top_iw_I\[12\].genblk1.cell0_I net505 net423 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0907_ col\[0\].zbuf_bot_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[0] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0838_ col\[6\].zbuf_top_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[235] sky130_fd_sc_hd__buf_2
X_0769_ col\[4\].zbuf_top_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[166] sky130_fd_sc_hd__buf_2
Xinput108 um_ow[166] vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_1
Xinput119 um_ow[176] vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_2854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_2617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_70 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_92 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_81 _0145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcol\[0\].zbuf_top_iw_I\[5\].genblk1.cell0_I net485 net436 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_2386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_2241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[2\].zbuf_top_iw_I\[0\].genblk1.cell0_I net511 net430 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[0\].z sky130_fd_sc_hd__and2_1
X_0554_ _0137_ _0138_ _0139_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__nand3b_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0485_ _0046_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1037_ col\[4\].genblk1.mux4_I\[18\].x _0257_ vssd1 vssd1 vccd1 vccd1 bus_ow\[18\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_7_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_2740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput90 um_ow[14] vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_bot_ena_I.genblk1.cell0_I_550 vssd1 vssd1 vccd1 vccd1 net550 col\[7\].zbuf_bot_ena_I.genblk1.cell0_I_550/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_7_1961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].zbuf_top_iw_I\[11\].genblk1.cell0_I net508 net441 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_10_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[5\].zbuf_bot_iw_I\[9\].genblk1.cell0_I net478 net421 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_bot_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[7\].zbuf_bot_iw_I\[4\].genblk1.cell0_I net488 net440 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_bot_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0606_ _0166_ vssd1 vssd1 vccd1 vccd1 col\[7\].zbuf_top_ena_I.e sky130_fd_sc_hd__clkbuf_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0537_ _0134_ _0135_ _0136_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__nand3b_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0468_ _0096_ _0089_ _0097_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__or3b_1
X_0399_ _0058_ _0059_ _0053_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_2345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_2211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[3\].zbuf_top_iw_I\[8\].genblk1.cell0_I net479 net426 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0322_ _0002_ _0006_ _0009_ _0013_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__or4_1
Xinput280 um_ow[320] vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_1
Xinput291 um_ow[330] vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_1
Xtt_mux_527 vssd1 vssd1 vccd1 vccd1 tt_mux_527/HI um_k_zero[7] sky130_fd_sc_hd__conb_1
XFILLER_0_15_2133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[5\].zbuf_top_iw_I\[3\].genblk1.cell0_I net490 net420 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout425 col\[3\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__clkbuf_2
Xfanout436 col\[0\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__clkbuf_2
Xfanout447 net448 vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout469 net476 vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__clkbuf_2
Xfanout458 net459 vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__clkbuf_4
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_2807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_2575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_2317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0940_ col\[0\].zbuf_top_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[33] sky130_fd_sc_hd__buf_2
XFILLER_0_15_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0871_ col\[7\].zbuf_bot_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[268] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0305_ _0001_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_8_2042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_2350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_2361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_2395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[0\].genblk1.mux4_I\[20\].cell0_I net157 net357 net383 net410 net464 net451 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[20\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_9_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0923_ col\[0\].zbuf_bot_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[16] sky130_fd_sc_hd__clkbuf_4
X_0854_ col\[6\].zbuf_top_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[251] sky130_fd_sc_hd__buf_2
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0785_ col\[5\].zbuf_bot_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[182] sky130_fd_sc_hd__buf_2
Xcol\[2\].genblk1.mux4_I\[19\].cell0_I net52 net78 net105 net131 net467 net456 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[19\].x sky130_fd_sc_hd__mux4_1
Xcol\[1\].zbuf_bot_iw_I\[15\].genblk1.cell0_I net499 net433 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_bot_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0570_ net458 vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__buf_4
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1053_ col\[6\].genblk1.mux4_I\[10\].x _0273_ vssd1 vssd1 vccd1 vccd1 bus_ow\[10\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_14_1508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0906_ col\[7\].zbuf_top_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[15] sky130_fd_sc_hd__buf_2
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0837_ col\[6\].zbuf_top_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[234] sky130_fd_sc_hd__buf_2
XFILLER_0_3_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0768_ col\[4\].zbuf_top_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[165] sky130_fd_sc_hd__buf_2
X_0699_ col\[2\].zbuf_top_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[96] sky130_fd_sc_hd__buf_2
Xinput109 um_ow[167] vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_2833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_2629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_71 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_93 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_82 _0145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_60 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcol\[3\].zbuf_bot_iw_I\[14\].genblk1.cell0_I net501 net427 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_bot_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_2253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0553_ _0137_ _0138_ _0139_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__nand3b_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0484_ _0044_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__clkbuf_2
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1036_ col\[4\].genblk1.mux4_I\[17\].x _0256_ vssd1 vssd1 vccd1 vccd1 bus_ow\[17\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_8_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput80 um_ow[140] vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput91 um_ow[150] vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[1\].zbuf_top_iw_I\[11\].genblk1.cell0_I net507 net431 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xzbuf_bus_sel_I\[1\].genblk1.cell1_I zbuf_bus_sel_I\[1\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 zbuf_bus_sel_I\[1\].z sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0605_ _0147_ _0148_ net461 _0163_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0536_ _0134_ _0135_ _0136_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__nand3b_2
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0467_ _0099_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__clkbuf_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0398_ _0060_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1019_ col\[4\].genblk1.mux4_I\[0\].x _0239_ vssd1 vssd1 vccd1 vccd1 bus_ow\[0\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[5\].zbuf_bot_iw_I\[13\].genblk1.cell0_I net504 net421 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_bot_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_2769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0321_ _0015_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__clkbuf_1
Xinput281 um_ow[321] vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__clkbuf_1
Xinput270 um_ow[311] vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_2213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput292 um_ow[331] vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_1
Xtt_mux_517 vssd1 vssd1 vccd1 vccd1 tt_mux_517/HI k_zero sky130_fd_sc_hd__conb_1
Xtt_mux_528 vssd1 vssd1 vccd1 vccd1 tt_mux_528/HI um_k_zero[8] sky130_fd_sc_hd__conb_1
XFILLER_0_8_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[3\].zbuf_top_iw_I\[10\].genblk1.cell0_I net509 net425 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout437 col\[7\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__clkbuf_2
Xfanout426 col\[3\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout448 col\[0\].zbuf_bot_ena_I.e vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__clkbuf_2
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0519_ _0128_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__clkbuf_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout459 net463 vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_2
Xcol\[1\].zbuf_bot_iw_I\[6\].genblk1.cell0_I net483 net434 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_bot_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_2519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[3\].zbuf_bot_iw_I\[1\].genblk1.cell0_I net493 net428 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_bot_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0870_ col\[7\].zbuf_bot_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[267] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0304_ net2 _0000_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__nor2_2
Xcol\[7\].zbuf_bot_iw_I\[12\].genblk1.cell0_I net506 net439 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_bot_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0999_ col\[2\].genblk1.mux4_I\[4\].x _0219_ vssd1 vssd1 vccd1 vccd1 bus_ow\[4\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[1\].zbuf_top_iw_I\[0\].genblk1.cell0_I net511 net432 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_2238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0922_ col\[0\].zbuf_bot_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0853_ col\[6\].zbuf_top_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[250] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0784_ col\[5\].zbuf_bot_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[181] sky130_fd_sc_hd__buf_2
XFILLER_0_12_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[7\].genblk1.cell1_I zbuf_bus_iw_I\[7\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[7\].a sky130_fd_sc_hd__buf_6
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput1 addr[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_14_2903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_90 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[4\].zbuf_bot_iw_I\[9\].genblk1.cell0_I net477 net443 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_bot_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_2547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[6\].zbuf_bot_iw_I\[4\].genblk1.cell0_I net488 net449 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_bot_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1052_ col\[6\].genblk1.mux4_I\[9\].x _0272_ vssd1 vssd1 vccd1 vccd1 bus_ow\[9\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_5_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0905_ col\[7\].zbuf_bot_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[14] sky130_fd_sc_hd__buf_2
XFILLER_0_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0836_ col\[6\].zbuf_bot_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[233] sky130_fd_sc_hd__buf_2
XFILLER_0_3_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0767_ col\[4\].zbuf_top_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[164] sky130_fd_sc_hd__buf_2
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0698_ col\[2\].zbuf_top_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[95] sky130_fd_sc_hd__buf_2
XFILLER_0_7_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_2889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_50 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_72 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_61 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_83 _0145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_94 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcol\[2\].zbuf_top_iw_I\[8\].genblk1.cell0_I net479 net429 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_15_2519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_2322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_2265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[4\].zbuf_top_iw_I\[3\].genblk1.cell0_I net489 net424 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0552_ _0137_ _0138_ _0139_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__nand3b_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0483_ _0107_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__clkbuf_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_2029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1035_ col\[4\].genblk1.mux4_I\[16\].x _0255_ vssd1 vssd1 vccd1 vccd1 bus_ow\[16\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_14_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput81 um_ow[141] vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_1
Xinput70 um_ow[131] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dlymetal6s2s_1
X_0819_ col\[6\].zbuf_bot_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[216] sky130_fd_sc_hd__buf_2
Xinput92 um_ow[151] vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_2907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xzbuf_bus_iw_I\[16\].genblk1.cell0_I net25 net513 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[16\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_7_2631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_2686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_2316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[4\].genblk1.mux4_I\[11\].cell0_I net150 net176 net203 net229 net471 net457 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[11\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_15_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0604_ _0165_ vssd1 vssd1 vccd1 vccd1 col\[7\].zbuf_bot_ena_I.e sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0535_ _0134_ _0135_ _0136_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__nand3b_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0466_ _0096_ _0089_ _0097_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__or3b_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0397_ _0058_ _0059_ _0053_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__or3_1
Xcol\[0\].zbuf_bot_iw_I\[13\].genblk1.cell0_I net503 net447 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_bot_iw_I\[13\].z sky130_fd_sc_hd__and2_1
X_1018_ col\[2\].genblk1.mux4_I\[23\].x _0238_ vssd1 vssd1 vccd1 vccd1 bus_ow\[23\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_2894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_2759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[3\].genblk1.cell0_I net11 net513 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[3\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0320_ _0002_ _0006_ _0009_ _0013_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__or4_1
Xinput271 um_ow[312] vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_1
Xinput260 um_ow[302] vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_1
Xinput282 um_ow[322] vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__clkbuf_1
Xinput293 um_ow[332] vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_1
Xtt_mux_529 vssd1 vssd1 vccd1 vccd1 tt_mux_529/HI um_k_zero[9] sky130_fd_sc_hd__conb_1
Xtt_mux_518 vssd1 vssd1 vccd1 vccd1 tt_mux_518/HI spine_ow[0] sky130_fd_sc_hd__conb_1
XFILLER_0_8_2225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_top_iw_I\[6\].genblk1.cell0_I net484 net438 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.mux4_I\[21\].cell0_I net267 net294 net320 net347 net475 net462 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[21\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[0\].zbuf_bot_ena_I.genblk1.cell0_I net536 net448 vssd1 vssd1 vccd1 vccd1 col\[0\].zbuf_bot_ena_I.z
+ sky130_fd_sc_hd__and2_1
Xfanout438 col\[7\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout427 col\[3\].zbuf_bot_ena_I.e vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__clkbuf_2
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0518_ _0124_ _0121_ _0122_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__or3b_1
Xfanout449 net450 vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__clkbuf_2
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0449_ zbuf_bus_sel_I\[3\].z vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_2770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[2\].zbuf_bot_iw_I\[12\].genblk1.cell0_I net505 net445 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_bot_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_10_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0303_ net33 vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_2055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_2099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0998_ col\[2\].genblk1.mux4_I\[3\].x _0218_ vssd1 vssd1 vccd1 vccd1 bus_ow\[3\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0921_ col\[0\].zbuf_bot_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[14] sky130_fd_sc_hd__buf_2
XFILLER_0_12_2149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0852_ col\[6\].zbuf_top_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[249] sky130_fd_sc_hd__buf_2
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0783_ col\[5\].zbuf_bot_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[180] sky130_fd_sc_hd__buf_2
XFILLER_0_3_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput2 addr[1] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XTAP_91 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_2661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[4\].zbuf_bot_iw_I\[11\].genblk1.cell0_I net507 net443 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_bot_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_2436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1051_ col\[6\].genblk1.mux4_I\[8\].x _0271_ vssd1 vssd1 vccd1 vccd1 bus_ow\[8\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_9_2183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0904_ col\[6\].zbuf_top_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[13] sky130_fd_sc_hd__buf_2
XFILLER_0_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0835_ col\[6\].zbuf_bot_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[232] sky130_fd_sc_hd__buf_2
XFILLER_0_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0766_ col\[4\].zbuf_top_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[163] sky130_fd_sc_hd__buf_2
XFILLER_0_3_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0697_ col\[2\].zbuf_top_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[94] sky130_fd_sc_hd__buf_2
XFILLER_0_7_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_2756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_40 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_2491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_73 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_62 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_51 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_84 _0147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_95 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_2356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_2378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0551_ _0137_ _0138_ _0139_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_1_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0482_ _0096_ _0097_ _0066_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__or3b_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[0\].zbuf_bot_iw_I\[6\].genblk1.cell0_I net483 net448 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_bot_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_2109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1034_ col\[4\].genblk1.mux4_I\[15\].x _0254_ vssd1 vssd1 vccd1 vccd1 bus_ow\[15\]
+ sky130_fd_sc_hd__ebufn_8
Xcol\[6\].zbuf_bot_iw_I\[10\].genblk1.cell0_I net510 net450 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_bot_iw_I\[10\].z sky130_fd_sc_hd__and2_1
Xcol\[4\].zbuf_top_ena_I.genblk1.cell0_I net545 net424 vssd1 vssd1 vccd1 vccd1 col\[4\].zbuf_top_ena_I.z
+ sky130_fd_sc_hd__and2_1
XFILLER_0_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput60 um_ow[122] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_2
Xinput71 um_ow[132] vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput82 um_ow[142] vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dlymetal6s2s_1
X_0818_ col\[5\].zbuf_top_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[215] sky130_fd_sc_hd__buf_2
Xinput93 um_ow[152] vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_1
X_0749_ col\[4\].zbuf_bot_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[146] sky130_fd_sc_hd__buf_2
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[2\].zbuf_bot_iw_I\[1\].genblk1.cell0_I net493 net446 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_bot_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_2676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_2564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_2030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[4\].genblk1.mux4_I\[15\].cell0_I net154 net181 net207 net233 net470 net457 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[15\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_13_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0603_ _0147_ _0148_ _0145_ _0163_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__and4b_1
XFILLER_0_0_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0534_ _0134_ _0135_ _0136_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__nand3b_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0465_ _0098_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__clkbuf_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0396_ _0044_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_8_2930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1017_ col\[2\].genblk1.mux4_I\[22\].x _0237_ vssd1 vssd1 vccd1 vccd1 bus_ow\[22\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_8_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[0\].zbuf_top_iw_I\[0\].genblk1.cell0_I net511 net436 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_1761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_2269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput272 um_ow[313] vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_1
Xinput261 um_ow[303] vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_1
Xinput250 um_ow[294] vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_1
Xinput283 um_ow[323] vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_1
Xinput294 um_ow[333] vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_1
Xtt_mux_519 vssd1 vssd1 vccd1 vccd1 tt_mux_519/HI spine_ow[25] sky130_fd_sc_hd__conb_1
XFILLER_0_8_2237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[3\].zbuf_bot_iw_I\[9\].genblk1.cell0_I net477 net427 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_bot_iw_I\[9\].z sky130_fd_sc_hd__and2_1
Xfanout428 col\[3\].zbuf_bot_ena_I.e vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout439 col\[7\].zbuf_bot_ena_I.e vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__clkbuf_2
X_0517_ _0127_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__clkbuf_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0448_ _0088_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__clkbuf_1
X_0379_ _0049_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_1901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[5\].zbuf_bot_iw_I\[4\].genblk1.cell0_I net488 net422 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_bot_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0997_ col\[2\].genblk1.mux4_I\[2\].x _0217_ vssd1 vssd1 vccd1 vccd1 bus_ow\[2\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[5\].zbuf_top_iw_I\[17\].genblk1.cell0_I net496 net419 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[17\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_iw_I\[8\].genblk1.cell0_I net479 net431 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[3\].zbuf_top_iw_I\[3\].genblk1.cell0_I net489 net426 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_2365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_2387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_130 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0920_ col\[0\].zbuf_bot_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[13] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0851_ col\[6\].zbuf_top_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[248] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0782_ col\[4\].zbuf_top_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[179] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput3 addr[2] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XTAP_92 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_70 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_2183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[7\].zbuf_top_iw_I\[16\].genblk1.cell0_I net498 net437 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[16\].z sky130_fd_sc_hd__and2_1
X_1050_ col\[6\].genblk1.mux4_I\[7\].x _0270_ vssd1 vssd1 vccd1 vccd1 bus_ow\[7\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_5_2015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_2059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0903_ col\[6\].zbuf_bot_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[12] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0834_ col\[6\].zbuf_bot_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[231] sky130_fd_sc_hd__buf_2
XFILLER_0_4_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0765_ col\[4\].zbuf_top_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[162] sky130_fd_sc_hd__buf_2
XFILLER_0_3_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0696_ col\[2\].zbuf_top_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[93] sky130_fd_sc_hd__buf_2
XFILLER_0_12_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_41 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_30 zbuf_bus_ena_I.z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_63 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_74 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_52 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_85 _0147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_96 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].genblk1.mux4_I\[10\].cell0_I net46 net312 net372 net399 net465 net452 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[10\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_13_2201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_2081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].zbuf_top_iw_I\[6\].genblk1.cell0_I net484 net442 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[1\].zbuf_bot_iw_I\[10\].genblk1.cell0_I net509 net433 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_bot_iw_I\[10\].z sky130_fd_sc_hd__and2_1
X_0550_ _0137_ _0138_ _0139_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__nand3b_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0481_ _0106_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__clkbuf_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1033_ col\[4\].genblk1.mux4_I\[14\].x _0253_ vssd1 vssd1 vccd1 vccd1 bus_ow\[14\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_5_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput61 um_ow[123] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_2
X_0817_ col\[5\].zbuf_top_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[214] sky130_fd_sc_hd__buf_2
XFILLER_0_13_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput72 um_ow[133] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput50 um_ow[113] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput83 um_ow[143] vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__clkbuf_1
Xinput94 um_ow[153] vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__clkbuf_1
X_0748_ col\[4\].zbuf_bot_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[145] sky130_fd_sc_hd__buf_2
X_0679_ col\[2\].zbuf_bot_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[76] sky130_fd_sc_hd__buf_2
XFILLER_0_7_2633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput410 um_ow[92] vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_1
Xcol\[2\].genblk1.mux4_I\[20\].cell0_I net53 net80 net106 net132 net467 net456 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[20\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_13_2042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[4\].genblk1.mux4_I\[19\].cell0_I net159 net185 net211 net238 net471 net458 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[19\].x sky130_fd_sc_hd__mux4_1
X_0602_ _0164_ vssd1 vssd1 vccd1 vccd1 col\[6\].zbuf_top_ena_I.e sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0533_ _0047_ vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__clkbuf_4
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0464_ _0096_ _0089_ _0097_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__or3b_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0395_ zbuf_bus_sel_I\[4\].z vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_2806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1016_ col\[2\].genblk1.mux4_I\[21\].x _0236_ vssd1 vssd1 vccd1 vccd1 bus_ow\[21\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_2706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_2463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_2237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput240 um_ow[285] vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_2
Xinput251 um_ow[295] vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_1
Xinput262 um_ow[304] vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_1
Xinput284 um_ow[324] vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_1
Xinput295 um_ow[334] vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_1
Xinput273 um_ow[314] vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_2205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_2115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_2126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout429 col\[2\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__clkbuf_2
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0516_ _0124_ _0121_ _0122_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__or3b_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0447_ _0083_ _0076_ _0084_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__or3b_1
X_0378_ _0043_ _0045_ _0047_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_2603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_2513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_2013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_top_iw_I\[17\].genblk1.cell0_I net495 net435 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_2934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0996_ col\[2\].genblk1.mux4_I\[1\].x _0216_ vssd1 vssd1 vccd1 vccd1 bus_ow\[1\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_120 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0850_ col\[6\].zbuf_top_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[247] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0781_ col\[4\].zbuf_top_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[178] sky130_fd_sc_hd__buf_2
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[1\].zbuf_bot_iw_I\[1\].genblk1.cell0_I net493 net434 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_bot_iw_I\[1\].z sky130_fd_sc_hd__and2_1
Xinput4 addr[3] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_2917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_60 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_93 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_2742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_2641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0979_ col\[0\].genblk1.mux4_I\[8\].x _0199_ vssd1 vssd1 vccd1 vccd1 bus_ow\[8\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_14_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xzbuf_bus_iw_I\[15\].genblk1.cell1_I zbuf_bus_iw_I\[15\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[15\].a sky130_fd_sc_hd__buf_6
XFILLER_0_11_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].zbuf_top_iw_I\[16\].genblk1.cell0_I net497 net429 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0902_ col\[5\].zbuf_top_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[11] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0833_ col\[6\].zbuf_bot_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[230] sky130_fd_sc_hd__buf_2
XFILLER_0_4_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0764_ col\[4\].zbuf_bot_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[161] sky130_fd_sc_hd__buf_2
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0695_ col\[2\].zbuf_top_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[92] sky130_fd_sc_hd__buf_2
XFILLER_0_12_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_20 col\[0\].zbuf_bot_iw_I\[8\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_31 net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_2493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_64 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_75 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_42 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_97 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_86 _0147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[0\].genblk1.mux4_I\[14\].cell0_I net90 net350 net377 net403 net464 net451 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[14\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_6_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xzbuf_bus_iw_I\[2\].genblk1.cell1_I zbuf_bus_iw_I\[2\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[2\].a sky130_fd_sc_hd__buf_6
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[2\].zbuf_bot_iw_I\[9\].genblk1.cell0_I net477 net445 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_bot_iw_I\[9\].z sky130_fd_sc_hd__and2_1
X_0480_ _0096_ _0097_ _0066_ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__or3b_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1032_ col\[4\].genblk1.mux4_I\[13\].x _0252_ vssd1 vssd1 vccd1 vccd1 bus_ow\[13\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput40 um_ow[104] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__dlymetal6s2s_1
X_0816_ col\[5\].zbuf_top_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[213] sky130_fd_sc_hd__buf_2
Xinput62 um_ow[124] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput73 um_ow[134] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dlymetal6s2s_1
Xcol\[4\].zbuf_bot_iw_I\[4\].genblk1.cell0_I net487 net444 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_bot_iw_I\[4\].z sky130_fd_sc_hd__and2_1
Xinput51 um_ow[114] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
X_0747_ col\[4\].zbuf_bot_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[144] sky130_fd_sc_hd__buf_2
Xinput84 um_ow[144] vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__clkbuf_1
Xinput95 um_ow[154] vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0678_ col\[2\].zbuf_bot_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[75] sky130_fd_sc_hd__buf_2
Xcol\[4\].zbuf_top_iw_I\[15\].genblk1.cell0_I net499 net423 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput400 um_ow[83] vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__clkbuf_1
Xinput411 um_ow[93] vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_top_iw_I\[8\].genblk1.cell0_I net479 net435 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0601_ _0145_ _0163_ net474 zbuf_bus_ena_I.z vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__and4b_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0532_ _0077_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0463_ _0044_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__clkbuf_4
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0394_ _0057_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__clkbuf_1
Xcol\[6\].genblk1.mux4_I\[1\].cell0_I net244 net272 net298 net325 net473 net460 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[1\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_4_2829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1015_ col\[2\].genblk1.mux4_I\[20\].x _0235_ vssd1 vssd1 vccd1 vccd1 bus_ow\[20\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_14_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].zbuf_top_iw_I\[3\].genblk1.cell0_I net489 net430 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_2249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput241 um_ow[286] vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput230 um_ow[276] vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_2
Xinput263 um_ow[305] vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__clkbuf_1
Xinput252 um_ow[296] vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_1
Xinput274 um_ow[315] vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_1
Xinput285 um_ow[325] vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_1
Xinput296 um_ow[335] vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].zbuf_top_iw_I\[14\].genblk1.cell0_I net502 net441 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_15_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout419 col\[5\].zbuf_top_ena_I.e vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__clkbuf_2
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0515_ _0126_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__clkbuf_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0446_ _0087_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__clkbuf_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xzbuf_bus_iw_I\[11\].genblk1.cell0_I net20 net515 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[11\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0377_ _0048_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[7\].zbuf_bot_iw_I\[7\].genblk1.cell0_I net482 net440 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_bot_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_11_1835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0995_ col\[2\].genblk1.mux4_I\[0\].x _0215_ vssd1 vssd1 vccd1 vccd1 bus_ow\[0\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_2_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0429_ _0075_ _0076_ _0077_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__or3b_1
XFILLER_0_4_2412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[5\].zbuf_top_iw_I\[6\].genblk1.cell0_I net484 net420 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_1733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_2301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].genblk1.mux4_I\[11\].cell0_I net255 net283 net309 net336 net473 net460 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[11\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_9_2345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_121 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_110 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[7\].zbuf_top_iw_I\[1\].genblk1.cell0_I net494 net438 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_12_1407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0780_ col\[4\].zbuf_top_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[177] sky130_fd_sc_hd__buf_2
XFILLER_0_11_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput5 addr[4] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XTAP_50 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_94 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_2798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0978_ col\[0\].genblk1.mux4_I\[7\].x _0198_ vssd1 vssd1 vccd1 vccd1 bus_ow\[7\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_2529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[4\].genblk1.mux4_I\[2\].cell0_I net139 net166 net193 net219 net472 net459 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[2\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_6_1839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_2141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0901_ col\[5\].zbuf_bot_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[10] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0832_ col\[6\].zbuf_bot_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[229] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0763_ col\[4\].zbuf_bot_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[160] sky130_fd_sc_hd__buf_2
XFILLER_0_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0694_ col\[2\].zbuf_top_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[91] sky130_fd_sc_hd__buf_2
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].genblk1.mux4_I\[0\].cell0_I net35 net201 net361 net388 net466 net453 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[0\].x sky130_fd_sc_hd__mux4_2
XANTENNA_21 col\[0\].zbuf_bot_iw_I\[8\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 col\[0\].zbuf_bot_iw_I\[1\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_32 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_65 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_54 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_98 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_76 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_87 _0147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcol\[0\].genblk1.mux4_I\[18\].cell0_I net134 net355 net381 net408 net464 net451 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[18\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_6_2348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_2225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1031_ col\[4\].genblk1.mux4_I\[12\].x _0251_ vssd1 vssd1 vccd1 vccd1 bus_ow\[12\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_2_2713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput30 spine_iw[5] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
X_0815_ col\[5\].zbuf_top_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[212] sky130_fd_sc_hd__buf_2
Xinput63 um_ow[125] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput41 um_ow[105] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput52 um_ow[115] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0746_ col\[3\].zbuf_top_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[143] sky130_fd_sc_hd__buf_2
Xinput74 um_ow[135] vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_13_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput85 um_ow[145] vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_1
Xinput96 um_ow[155] vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0677_ col\[2\].zbuf_bot_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[74] sky130_fd_sc_hd__buf_2
XFILLER_0_7_2613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput401 um_ow[84] vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__clkbuf_1
Xinput412 um_ow[94] vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_2101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_2099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_2790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0600_ _0264_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0531_ _0075_ vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0462_ _0042_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__clkbuf_4
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0393_ _0043_ _0045_ _0053_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__or3_1
Xcol\[3\].zbuf_bot_iw_I\[17\].genblk1.cell0_I net495 net427 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_bot_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1014_ col\[2\].genblk1.mux4_I\[19\].x _0234_ vssd1 vssd1 vccd1 vccd1 bus_ow\[19\]
+ sky130_fd_sc_hd__ebufn_8
Xcol\[6\].genblk1.mux4_I\[5\].cell0_I net249 net276 net303 net329 net473 net460 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[5\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_15_2865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0729_ col\[3\].zbuf_top_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[126] sky130_fd_sc_hd__buf_2
XFILLER_0_0_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_2465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_bot_iw_I\[1\].genblk1.cell0_I net493 net448 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_bot_iw_I\[1\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_iw_I\[14\].genblk1.cell0_I net501 net431 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[14\].z sky130_fd_sc_hd__and2_1
Xinput220 um_ow[267] vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput231 um_ow[277] vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_2
Xinput242 um_ow[287] vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput253 um_ow[297] vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_1
Xinput275 um_ow[316] vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_1
Xinput286 um_ow[326] vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_1
Xinput264 um_ow[306] vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_1
Xinput297 um_ow[336] vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_15_2139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_2830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[2\].genblk1.mux4_I\[3\].cell0_I net417 net61 net87 net114 net469 net455 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[3\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_3_2896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xzbuf_bus_sel_I\[4\].genblk1.cell1_I zbuf_bus_sel_I\[4\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 zbuf_bus_sel_I\[4\].z sky130_fd_sc_hd__buf_8
XFILLER_0_10_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0514_ _0124_ _0121_ _0122_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__or3b_1
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0445_ _0083_ _0076_ _0084_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__or3b_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0376_ _0043_ _0045_ _0047_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_2741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_top_ena_I.genblk1.cell0_I net537 net436 vssd1 vssd1 vccd1 vccd1 col\[0\].zbuf_top_ena_I.z
+ sky130_fd_sc_hd__and2_1
XFILLER_0_8_2785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[5\].zbuf_bot_iw_I\[16\].genblk1.cell0_I net498 net421 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_bot_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_2058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_2903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_2671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0994_ col\[0\].genblk1.mux4_I\[23\].x _0214_ vssd1 vssd1 vccd1 vccd1 bus_ow\[23\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_2_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0428_ _0044_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__buf_4
X_0359_ _0036_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__clkbuf_1
Xcol\[3\].zbuf_top_iw_I\[13\].genblk1.cell0_I net503 net425 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[1\].zbuf_bot_iw_I\[9\].genblk1.cell0_I net477 net433 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_bot_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_2335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_100 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_122 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_111 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcol\[6\].genblk1.mux4_I\[15\].cell0_I net261 net287 net314 net340 net474 net461 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[15\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_9_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_2844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_2899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[3\].zbuf_bot_iw_I\[4\].genblk1.cell0_I net487 net428 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_bot_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput6 spine_iw[10] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_40 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_51 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_84 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_95 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0977_ col\[0\].genblk1.mux4_I\[6\].x _0197_ vssd1 vssd1 vccd1 vccd1 bus_ow\[6\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_6_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[7\].zbuf_bot_iw_I\[15\].genblk1.cell0_I net500 net439 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_bot_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_2107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[4\].genblk1.mux4_I\[6\].cell0_I net143 net171 net197 net224 net470 net457 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[6\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_2197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_2165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0900_ col\[4\].zbuf_top_ena_I.z vssd1 vssd1 vccd1 vccd1 um_ena[9] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[5\].zbuf_top_iw_I\[12\].genblk1.cell0_I net506 net419 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[12\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_iw_I\[3\].genblk1.cell0_I net489 net432 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[3\].z sky130_fd_sc_hd__and2_1
X_0831_ col\[6\].zbuf_bot_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[228] sky130_fd_sc_hd__buf_2
XFILLER_0_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0762_ col\[4\].zbuf_bot_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[159] sky130_fd_sc_hd__buf_2
XFILLER_0_4_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0693_ col\[2\].zbuf_top_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[90] sky130_fd_sc_hd__buf_2
XFILLER_0_11_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_11 col\[0\].zbuf_bot_iw_I\[1\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 col\[0\].zbuf_bot_iw_I\[9\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_66 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_44 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_33 net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_55 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcol\[0\].genblk1.mux4_I\[4\].cell0_I net363 net245 net366 net392 net466 net453 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[4\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_99 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_77 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_88 bus_ow\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xzbuf_bus_sel_I\[0\].genblk1.cell0_I net32 net516 vssd1 vssd1 vccd1 vccd1 zbuf_bus_sel_I\[0\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_0_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1030_ col\[4\].genblk1.mux4_I\[11\].x _0250_ vssd1 vssd1 vccd1 vccd1 bus_ow\[11\]
+ sky130_fd_sc_hd__ebufn_8
Xzbuf_bus_ena_I.genblk1.cell1_I zbuf_bus_ena_I.genblk1.l vssd1 vssd1 vccd1 vccd1 zbuf_bus_ena_I.z
+ sky130_fd_sc_hd__buf_8
XFILLER_0_6_2861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].zbuf_bot_iw_I\[7\].genblk1.cell0_I net482 net449 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_bot_iw_I\[7\].z sky130_fd_sc_hd__and2_1
X_0814_ col\[5\].zbuf_top_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[211] sky130_fd_sc_hd__buf_2
Xinput31 spine_iw[6] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_2471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput20 spine_iw[23] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput64 um_ow[126] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_2
Xinput42 um_ow[106] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput53 um_ow[116] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0745_ col\[3\].zbuf_top_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[142] sky130_fd_sc_hd__buf_2
Xinput75 um_ow[136] vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput86 um_ow[146] vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput97 um_ow[156] vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_1
X_0676_ col\[2\].zbuf_bot_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[73] sky130_fd_sc_hd__buf_2
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[7\].zbuf_top_iw_I\[11\].genblk1.cell0_I net508 net437 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[11\].z sky130_fd_sc_hd__and2_1
Xinput402 um_ow[85] vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__clkbuf_1
Xinput413 um_ow[95] vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_2113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[5\].zbuf_bot_ena_I.genblk1.cell0_I net546 net422 vssd1 vssd1 vccd1 vccd1 col\[5\].zbuf_bot_ena_I.z
+ sky130_fd_sc_hd__and2_1
XFILLER_0_1_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0530_ zbuf_bus_sel_I\[4\].z zbuf_bus_sel_I\[2\].z zbuf_bus_sel_I\[3\].z vssd1 vssd1
+ vccd1 vccd1 _0264_ sky130_fd_sc_hd__nand3b_4
XFILLER_0_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0461_ _0095_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__clkbuf_1
X_0392_ _0056_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__clkbuf_1
X_1013_ col\[2\].genblk1.mux4_I\[18\].x _0233_ vssd1 vssd1 vccd1 vccd1 bus_ow\[18\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_2_2511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[4\].zbuf_top_iw_I\[6\].genblk1.cell0_I net483 net424 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.mux4_I\[9\].cell0_I net253 net281 net307 net333 net474 net461 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[9\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_5_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0728_ col\[3\].zbuf_bot_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[125] sky130_fd_sc_hd__buf_2
XFILLER_0_12_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0659_ col\[1\].zbuf_top_iw_I\[2\].z vssd1 vssd1 vccd1 vccd1 um_iw[56] sky130_fd_sc_hd__buf_2
XFILLER_0_0_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[6\].zbuf_top_iw_I\[1\].genblk1.cell0_I net494 net442 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_2477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput210 um_ow[258] vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput232 um_ow[278] vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput221 um_ow[268] vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput254 um_ow[298] vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_1
Xinput243 um_ow[288] vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_1
Xinput276 um_ow[317] vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_1
Xinput287 um_ow[327] vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_1
Xinput265 um_ow[307] vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_1
Xinput298 um_ow[337] vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_15_2129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.mux4_I\[7\].cell0_I net39 net65 net92 net118 net468 net454 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[7\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_2_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0513_ _0125_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0444_ _0086_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__clkbuf_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0375_ _0046_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_7_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.mux4_I\[10\].cell0_I net42 net69 net95 net121 net468 net454 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[10\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_13_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[0\].zbuf_bot_iw_I\[16\].genblk1.cell0_I net497 net447 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_bot_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_2274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0993_ col\[0\].genblk1.mux4_I\[22\].x _0213_ vssd1 vssd1 vccd1 vccd1 bus_ow\[22\]
+ sky130_fd_sc_hd__ebufn_8
Xzbuf_bus_iw_I\[6\].genblk1.cell0_I net14 net514 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[6\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_14_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0427_ _0046_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__buf_2
X_0358_ _0023_ _0024_ _0025_ _0026_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__or4_1
Xcol\[7\].zbuf_top_iw_I\[9\].genblk1.cell0_I net478 net437 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[20\].cell0_I net160 net186 net213 net239 net471 net458 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[20\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_9_2314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_101 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_112 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_123 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_2071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.mux4_I\[19\].cell0_I net265 net292 net318 net344 net475 net462 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[19\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_3_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput7 spine_iw[11] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XTAP_41 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_2712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_2881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_85 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[2\].zbuf_bot_iw_I\[15\].genblk1.cell0_I net499 net445 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_bot_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XTAP_63 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_52 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_2734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_96 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0976_ col\[0\].genblk1.mux4_I\[5\].x _0196_ vssd1 vssd1 vccd1 vccd1 bus_ow\[5\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].zbuf_top_iw_I\[12\].genblk1.cell0_I net505 net435 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0830_ col\[6\].zbuf_bot_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[227] sky130_fd_sc_hd__buf_2
XFILLER_0_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0761_ col\[4\].zbuf_bot_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[158] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0692_ col\[2\].zbuf_bot_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[89] sky130_fd_sc_hd__buf_2
XFILLER_0_11_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_12 col\[0\].zbuf_bot_iw_I\[3\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 col\[0\].zbuf_bot_iw_I\[9\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_34 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_56 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_45 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_78 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_67 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_89 bus_ow\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0959_ bus_ow\[12\] _0179_ vssd1 vssd1 vccd1 vccd1 spine_ow[13] sky130_fd_sc_hd__ebufn_8
Xcol\[0\].genblk1.mux4_I\[8\].cell0_I net407 net290 net370 net397 net465 net452 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[8\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_13_1537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_bot_iw_I\[14\].genblk1.cell0_I net501 net443 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_bot_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_11_1294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0813_ col\[5\].zbuf_top_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[210] sky130_fd_sc_hd__buf_2
Xinput10 spine_iw[14] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput21 spine_iw[24] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
Xinput32 spine_iw[7] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
Xinput43 um_ow[107] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_0_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput54 um_ow[117] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput65 um_ow[127] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dlymetal6s2s_1
X_0744_ col\[3\].zbuf_top_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[141] sky130_fd_sc_hd__buf_2
Xinput76 um_ow[137] vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput87 um_ow[147] vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[10\].genblk1.cell1_I zbuf_bus_iw_I\[10\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[10\].a sky130_fd_sc_hd__buf_6
Xinput98 um_ow[157] vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_1
X_0675_ col\[2\].zbuf_bot_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[72] sky130_fd_sc_hd__buf_2
XFILLER_0_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[2\].zbuf_top_iw_I\[11\].genblk1.cell0_I net507 net429 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_2293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput403 um_ow[86] vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__clkbuf_1
Xinput414 um_ow[96] vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_6_2125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0460_ _0083_ _0089_ _0084_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__or3b_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0391_ _0043_ _0045_ _0053_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1012_ col\[2\].genblk1.mux4_I\[17\].x _0232_ vssd1 vssd1 vccd1 vccd1 bus_ow\[17\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_2845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0727_ col\[3\].zbuf_bot_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[124] sky130_fd_sc_hd__buf_2
Xcol\[0\].zbuf_bot_iw_I\[9\].genblk1.cell0_I net477 net447 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_bot_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0658_ col\[1\].zbuf_top_iw_I\[1\].z vssd1 vssd1 vccd1 vccd1 um_iw[55] sky130_fd_sc_hd__buf_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[6\].zbuf_bot_iw_I\[13\].genblk1.cell0_I net504 net450 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_bot_iw_I\[13\].z sky130_fd_sc_hd__and2_1
X_0589_ net472 net459 _0240_ zbuf_bus_ena_I.z vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__or4b_1
XFILLER_0_14_2322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[2\].zbuf_bot_iw_I\[4\].genblk1.cell0_I net487 net446 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_bot_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput200 um_ow[249] vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput211 um_ow[259] vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput222 um_ow[269] vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput233 um_ow[279] vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput244 um_ow[289] vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_1
Xinput277 um_ow[318] vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_1
Xinput288 um_ow[328] vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_1
Xinput266 um_ow[308] vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_1
Xinput255 um_ow[299] vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_1
Xinput299 um_ow[338] vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_15_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[4\].zbuf_top_iw_I\[10\].genblk1.cell0_I net509 net423 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0512_ _0124_ _0121_ _0122_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__or3b_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0443_ _0083_ _0076_ _0084_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__or3b_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0374_ zbuf_bus_sel_I\[3\].z vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_2631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_2629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[2\].genblk1.mux4_I\[14\].cell0_I net47 net73 net99 net126 net467 net456 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[14\].x sky130_fd_sc_hd__mux4_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_2286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[0\].zbuf_top_iw_I\[3\].genblk1.cell0_I net489 net436 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_2927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_2826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0992_ col\[0\].genblk1.mux4_I\[21\].x _0212_ vssd1 vssd1 vccd1 vccd1 bus_ow\[21\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_3_1961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0426_ _0042_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__buf_4
X_0357_ _0035_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_2573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_2172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_113 col\[0\].zbuf_bot_iw_I\[13\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_102 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_124 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_2813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[5\].zbuf_bot_iw_I\[7\].genblk1.cell0_I net482 net422 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_bot_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput8 spine_iw[12] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XTAP_42 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_53 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[7\].zbuf_bot_iw_I\[2\].genblk1.cell0_I net492 net440 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_bot_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XTAP_97 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0975_ col\[0\].genblk1.mux4_I\[4\].x _0195_ vssd1 vssd1 vccd1 vccd1 bus_ow\[4\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0409_ _0046_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[3\].zbuf_top_iw_I\[6\].genblk1.cell0_I net483 net426 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_12_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0760_ col\[4\].zbuf_bot_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[157] sky130_fd_sc_hd__buf_2
X_0691_ col\[2\].zbuf_bot_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[88] sky130_fd_sc_hd__buf_2
Xcol\[5\].zbuf_top_iw_I\[1\].genblk1.cell0_I net494 net420 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_2521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_13 col\[0\].zbuf_bot_iw_I\[4\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_46 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_24 spine_iw[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_57 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_79 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_68 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0958_ bus_ow\[11\] _0178_ vssd1 vssd1 vccd1 vccd1 spine_ow[12] sky130_fd_sc_hd__ebufn_8
XFILLER_0_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0889_ col\[7\].zbuf_top_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[286] sky130_fd_sc_hd__buf_2
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0812_ col\[5\].zbuf_top_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[209] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput22 spine_iw[25] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
Xinput11 spine_iw[15] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput55 um_ow[118] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput44 um_ow[108] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput33 spine_iw[8] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
X_0743_ col\[3\].zbuf_top_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[140] sky130_fd_sc_hd__buf_2
Xinput66 um_ow[128] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput77 um_ow[138] vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput88 um_ow[148] vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0674_ col\[1\].zbuf_top_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[71] sky130_fd_sc_hd__buf_2
XFILLER_0_0_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput99 um_ow[158] vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_1959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput404 um_ow[87] vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__clkbuf_1
Xinput415 um_ow[97] vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_6_2137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[2\].zbuf_bot_ena_I.genblk1.cell0_I_540 vssd1 vssd1 vccd1 vccd1 net540 col\[2\].zbuf_bot_ena_I.genblk1.cell0_I_540/LO
+ sky130_fd_sc_hd__conb_1
X_0390_ _0055_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_2903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1011_ col\[2\].genblk1.mux4_I\[16\].x _0231_ vssd1 vssd1 vccd1 vccd1 bus_ow\[16\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_2813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].zbuf_top_iw_I\[9\].genblk1.cell0_I net478 net441 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_15_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[1\].zbuf_bot_iw_I\[13\].genblk1.cell0_I net503 net433 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_bot_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_1845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0726_ col\[3\].zbuf_bot_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[123] sky130_fd_sc_hd__buf_2
XFILLER_0_4_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0657_ col\[1\].zbuf_top_iw_I\[0\].z vssd1 vssd1 vccd1 vccd1 um_iw[54] sky130_fd_sc_hd__buf_2
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0588_ _0156_ vssd1 vssd1 vccd1 vccd1 col\[3\].zbuf_top_ena_I.e sky130_fd_sc_hd__clkbuf_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_2457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_2378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_2089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput201 um_ow[24] vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_2
Xinput212 um_ow[25] vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__clkbuf_2
Xinput245 um_ow[28] vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_2
Xinput234 um_ow[27] vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_2
Xinput223 um_ow[26] vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_2
Xinput278 um_ow[319] vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_1
Xinput256 um_ow[29] vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_2
Xinput267 um_ow[309] vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_1
Xinput289 um_ow[329] vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_2822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0511_ _0042_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__clkbuf_2
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0442_ _0085_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__clkbuf_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0373_ _0044_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__buf_2
XFILLER_0_15_2676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_2665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0709_ col\[2\].zbuf_top_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[106] sky130_fd_sc_hd__buf_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[2\].genblk1.mux4_I\[18\].cell0_I net51 net77 net104 net130 net467 net456 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[18\].x sky130_fd_sc_hd__mux4_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_2221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[3\].zbuf_bot_iw_I\[12\].genblk1.cell0_I net505 net427 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_bot_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_2805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0991_ col\[0\].genblk1.mux4_I\[20\].x _0211_ vssd1 vssd1 vccd1 vccd1 bus_ow\[20\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_3_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[3\].zbuf_bot_ena_I.genblk1.cell0_I_542 vssd1 vssd1 vccd1 vccd1 net542 col\[3\].zbuf_bot_ena_I.genblk1.cell0_I_542/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_10_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0425_ _0074_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__clkbuf_2
X_0356_ _0023_ _0024_ _0025_ _0026_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_2541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_2585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_125 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_103 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_114 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_2073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput9 spine_iw[13] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XTAP_32 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_76 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_43 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_54 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_98 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0974_ col\[0\].genblk1.mux4_I\[3\].x _0194_ vssd1 vssd1 vccd1 vccd1 bus_ow\[3\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_10_2381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0408_ _0065_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__clkbuf_1
X_0339_ _0012_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__dlymetal6s2s_1
Xcol\[5\].zbuf_bot_iw_I\[11\].genblk1.cell0_I net508 net421 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_bot_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_2213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0690_ col\[2\].zbuf_bot_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[87] sky130_fd_sc_hd__buf_2
XFILLER_0_2_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_14 col\[0\].zbuf_bot_iw_I\[4\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_25 spine_iw[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_36 net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_47 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_69 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcol\[1\].zbuf_bot_iw_I\[4\].genblk1.cell0_I net487 net434 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_bot_iw_I\[4\].z sky130_fd_sc_hd__and2_1
X_0957_ bus_ow\[10\] _0177_ vssd1 vssd1 vccd1 vccd1 spine_ow[11] sky130_fd_sc_hd__ebufn_8
XANTENNA_58 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0888_ col\[7\].zbuf_top_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[285] sky130_fd_sc_hd__buf_2
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_bot_ena_I.genblk1.cell0_I_544 vssd1 vssd1 vccd1 vccd1 net544 col\[4\].zbuf_bot_ena_I.genblk1.cell0_I_544/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_2043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0811_ col\[5\].zbuf_top_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[208] sky130_fd_sc_hd__buf_2
Xcol\[7\].zbuf_bot_iw_I\[10\].genblk1.cell0_I net510 net439 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_bot_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_2463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 spine_iw[16] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
X_0742_ col\[3\].zbuf_top_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[139] sky130_fd_sc_hd__buf_2
Xinput45 um_ow[109] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput23 spine_iw[26] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 spine_iw[9] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
Xinput67 um_ow[129] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput78 um_ow[139] vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput89 um_ow[149] vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_1
Xinput56 um_ow[119] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0673_ col\[1\].zbuf_top_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[70] sky130_fd_sc_hd__buf_2
XFILLER_0_0_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput405 um_ow[88] vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__clkbuf_1
Xinput416 um_ow[98] vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_6_2149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_2015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1010_ col\[2\].genblk1.mux4_I\[15\].x _0230_ vssd1 vssd1 vccd1 vccd1 bus_ow\[15\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_2836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xzbuf_bus_iw_I\[5\].genblk1.cell1_I zbuf_bus_iw_I\[5\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[5\].a sky130_fd_sc_hd__buf_6
XFILLER_0_0_2260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0725_ col\[3\].zbuf_bot_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[122] sky130_fd_sc_hd__buf_2
X_0656_ col\[1\].zbuf_bot_iw_I\[17\].z vssd1 vssd1 vccd1 vccd1 um_iw[53] sky130_fd_sc_hd__buf_2
XFILLER_0_0_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0587_ _0147_ _0148_ _0145_ _0153_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__and4_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_2302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[4\].zbuf_bot_iw_I\[7\].genblk1.cell0_I net481 net444 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_bot_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_2057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput202 um_ow[250] vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput224 um_ow[270] vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput235 um_ow[280] vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_2
Xinput213 um_ow[260] vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__dlymetal6s2s_1
Xcol\[5\].zbuf_bot_ena_I.genblk1.cell0_I_546 vssd1 vssd1 vccd1 vccd1 net546 col\[5\].zbuf_bot_ena_I.genblk1.cell0_I_546/LO
+ sky130_fd_sc_hd__conb_1
Xinput268 um_ow[30] vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_2
Xinput279 um_ow[31] vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_2
Xinput257 um_ow[2] vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput246 um_ow[290] vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_2801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[6\].zbuf_bot_iw_I\[2\].genblk1.cell0_I net492 net449 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_bot_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0510_ _0123_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__clkbuf_1
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0441_ _0083_ _0076_ _0084_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__or3b_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0372_ zbuf_bus_sel_I\[2\].z vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_2756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[0\].genblk1.mux4_I\[23\].cell0_I net190 net360 net387 net413 net464 net451 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[23\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_1_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0708_ col\[2\].zbuf_top_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[105] sky130_fd_sc_hd__buf_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].zbuf_top_iw_I\[6\].genblk1.cell0_I net483 net430 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_2154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_top_iw_I\[1\].genblk1.cell0_I net493 net424 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0990_ col\[0\].genblk1.mux4_I\[19\].x _0210_ vssd1 vssd1 vccd1 vccd1 bus_ow\[19\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_3_1941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[1\].zbuf_bot_ena_I.genblk1.cell0_I net538 net434 vssd1 vssd1 vccd1 vccd1 col\[1\].zbuf_bot_ena_I.z
+ sky130_fd_sc_hd__and2_1
XFILLER_0_2_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0424_ zbuf_bus_sel_I\[4\].z zbuf_bus_sel_I\[3\].z zbuf_bus_sel_I\[2\].z vssd1 vssd1
+ vccd1 vccd1 _0074_ sky130_fd_sc_hd__or3b_1
Xcol\[6\].zbuf_top_iw_I\[17\].genblk1.cell0_I net496 net441 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[17\].z sky130_fd_sc_hd__and2_1
X_0355_ _0034_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_1830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_2597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xzbuf_bus_iw_I\[14\].genblk1.cell0_I net23 net513 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[14\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_14_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_104 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_2041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_115 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_126 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_2085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[6\].zbuf_bot_ena_I.genblk1.cell0_I_548 vssd1 vssd1 vccd1 vccd1 net548 col\[6\].zbuf_bot_ena_I.genblk1.cell0_I_548/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_9_2840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_33 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_66 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_44 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_2726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_99 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0973_ col\[0\].genblk1.mux4_I\[2\].x _0193_ vssd1 vssd1 vccd1 vccd1 bus_ow\[2\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_3_1793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_bot_iw_I\[11\].genblk1.cell0_I net507 net447 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_bot_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_10_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0407_ _0058_ _0059_ _0053_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__or3_1
X_0338_ _0008_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_15_2260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_2225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[5\].zbuf_top_iw_I\[9\].genblk1.cell0_I net478 net419 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xzbuf_bus_iw_I\[1\].genblk1.cell0_I net9 net513 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[1\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_0_2645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[7\].zbuf_top_iw_I\[4\].genblk1.cell0_I net488 net438 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_15 col\[0\].zbuf_bot_iw_I\[5\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcol\[4\].genblk1.mux4_I\[10\].cell0_I net149 net175 net202 net228 net470 net457 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[10\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_3_2280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_48 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 spine_iw[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0956_ bus_ow\[9\] _0176_ vssd1 vssd1 vccd1 vccd1 spine_ow[10] sky130_fd_sc_hd__ebufn_8
XANTENNA_59 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0887_ col\[7\].zbuf_top_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[284] sky130_fd_sc_hd__buf_2
XFILLER_0_3_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].zbuf_bot_iw_I\[10\].genblk1.cell0_I net509 net445 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_bot_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0810_ col\[5\].zbuf_top_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[207] sky130_fd_sc_hd__buf_2
Xinput13 spine_iw[17] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
X_0741_ col\[3\].zbuf_top_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[138] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput35 um_ow[0] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_2
Xinput46 um_ow[10] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput24 spine_iw[27] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput68 um_ow[12] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput57 um_ow[11] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput79 um_ow[13] vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0672_ col\[1\].zbuf_top_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[69] sky130_fd_sc_hd__buf_2
XFILLER_0_7_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0939_ col\[0\].zbuf_top_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[32] sky130_fd_sc_hd__buf_2
XFILLER_0_15_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.mux4_I\[20\].cell0_I net266 net293 net319 net346 net475 net462 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[20\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_11_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput406 um_ow[89] vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__clkbuf_1
Xinput417 um_ow[99] vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_6_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[5\].zbuf_top_ena_I.genblk1.cell0_I net547 net420 vssd1 vssd1 vccd1 vccd1 col\[5\].zbuf_top_ena_I.z
+ sky130_fd_sc_hd__and2_1
XFILLER_0_15_2826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0724_ col\[3\].zbuf_bot_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[121] sky130_fd_sc_hd__buf_2
X_0655_ col\[1\].zbuf_bot_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[52] sky130_fd_sc_hd__buf_2
XFILLER_0_12_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0586_ _0155_ vssd1 vssd1 vccd1 vccd1 col\[3\].zbuf_bot_ena_I.e sky130_fd_sc_hd__clkbuf_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_2325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_2358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput225 um_ow[271] vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput236 um_ow[281] vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__clkbuf_2
Xinput203 um_ow[251] vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput214 um_ow[261] vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput258 um_ow[300] vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_1
Xinput269 um_ow[310] vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_1
Xinput247 um_ow[291] vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_2813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0440_ _0044_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__dlymetal6s2s_1
X_0371_ _0042_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_15_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_2323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0707_ col\[2\].zbuf_top_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[104] sky130_fd_sc_hd__buf_2
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0569_ _0144_ vssd1 vssd1 vccd1 vccd1 col\[0\].zbuf_bot_ena_I.e sky130_fd_sc_hd__inv_2
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_2109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].zbuf_bot_iw_I\[4\].genblk1.cell0_I net487 net448 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_bot_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_1953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[1\].zbuf_top_iw_I\[17\].genblk1.cell0_I net495 net431 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0423_ _0073_ vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__clkbuf_1
X_0354_ _0023_ _0024_ _0025_ _0026_ vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_2420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_116 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_127 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_2053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_67 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_34 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_45 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_89 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_2749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_2451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0972_ col\[0\].genblk1.mux4_I\[1\].x _0192_ vssd1 vssd1 vccd1 vccd1 bus_ow\[1\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_12_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0406_ _0064_ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__clkbuf_1
X_0337_ _0005_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_2237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[7\].zbuf_top_ena_I.genblk1.cell0_I_551 vssd1 vssd1 vccd1 vccd1 net551 col\[7\].zbuf_top_ena_I.genblk1.cell0_I_551/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_8_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[3\].zbuf_top_iw_I\[16\].genblk1.cell0_I net497 net425 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_2657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_2681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[3\].zbuf_bot_iw_I\[7\].genblk1.cell0_I net481 net428 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_bot_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_2557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_2467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_16 col\[0\].zbuf_bot_iw_I\[5\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 spine_iw[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_49 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0955_ bus_ow\[8\] _0175_ vssd1 vssd1 vccd1 vccd1 spine_ow[9] sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0886_ col\[7\].zbuf_top_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[283] sky130_fd_sc_hd__buf_2
XFILLER_0_3_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[14\].cell0_I net153 net180 net206 net232 net470 net457 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[14\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[5\].zbuf_bot_iw_I\[2\].genblk1.cell0_I net492 net422 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_bot_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_2001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_2476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0740_ col\[3\].zbuf_top_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[137] sky130_fd_sc_hd__buf_2
Xinput36 um_ow[100] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput25 spine_iw[28] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
Xinput14 spine_iw[18] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
Xinput58 um_ow[120] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput69 um_ow[130] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_2
Xinput47 um_ow[110] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dlymetal6s2s_1
X_0671_ col\[1\].zbuf_top_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[68] sky130_fd_sc_hd__buf_2
XFILLER_0_0_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[1\].zbuf_top_iw_I\[6\].genblk1.cell0_I net483 net432 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_1929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[5\].zbuf_top_iw_I\[15\].genblk1.cell0_I net500 net419 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_2376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0938_ col\[0\].zbuf_top_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[31] sky130_fd_sc_hd__buf_2
XFILLER_0_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0869_ col\[7\].zbuf_bot_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[266] sky130_fd_sc_hd__buf_2
XFILLER_0_2_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput407 um_ow[8] vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__clkbuf_2
Xinput418 um_ow[9] vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_2
Xcol\[3\].zbuf_top_iw_I\[1\].genblk1.cell0_I net493 net426 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_2641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_2516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_sel_I\[3\].genblk1.cell0_I net29 net516 vssd1 vssd1 vccd1 vccd1 zbuf_bus_sel_I\[3\].genblk1.l
+ sky130_fd_sc_hd__and2_2
XFILLER_0_2_2549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0723_ col\[3\].zbuf_bot_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[120] sky130_fd_sc_hd__buf_2
X_0654_ col\[1\].zbuf_bot_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[51] sky130_fd_sc_hd__buf_2
XFILLER_0_0_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0585_ _0147_ _0148_ _0145_ _0153_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__and4b_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput226 um_ow[272] vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput204 um_ow[252] vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput215 um_ow[262] vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput237 um_ow[282] vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_2
Xinput248 um_ow[292] vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_1
Xinput259 um_ow[301] vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_2869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_top_iw_I\[14\].genblk1.cell0_I net502 net437 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0370_ zbuf_bus_sel_I\[4\].z vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_2714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0706_ col\[2\].zbuf_top_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[103] sky130_fd_sc_hd__buf_2
XFILLER_0_4_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0568_ net469 net455 _0192_ zbuf_bus_ena_I.z vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__or4b_4
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0499_ _0111_ _0108_ _0109_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__or3b_1
Xcol\[4\].zbuf_top_iw_I\[9\].genblk1.cell0_I net477 net423 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[6\].zbuf_top_iw_I\[4\].genblk1.cell0_I net488 net442 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_12_2819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0422_ _0042_ _0044_ _0066_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__or3_1
X_0353_ _0033_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_117 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_128 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_2896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_35 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_46 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_57 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_79 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_2605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0971_ col\[0\].genblk1.mux4_I\[0\].x _0191_ vssd1 vssd1 vccd1 vccd1 bus_ow\[0\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0405_ _0058_ _0059_ _0053_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__or3_1
X_0336_ _0001_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_8_2330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_2205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_2352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xzbuf_bus_iw_I\[9\].genblk1.cell0_I net18 net514 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[9\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_4_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout510 col\[0\].zbuf_bot_iw_I\[10\].a vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__clkbuf_4
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_2603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_2569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_17 col\[0\].zbuf_bot_iw_I\[6\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_2293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_39 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 zbuf_bus_ena_I.z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0954_ bus_ow\[7\] _0174_ vssd1 vssd1 vccd1 vccd1 spine_ow[8] sky130_fd_sc_hd__ebufn_8
XFILLER_0_10_2181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0885_ col\[7\].zbuf_top_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[282] sky130_fd_sc_hd__buf_2
XFILLER_0_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[18\].cell0_I net158 net184 net210 net237 net470 net457 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[18\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0319_ _0014_ vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_2013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_2834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput37 um_ow[101] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput26 spine_iw[29] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
Xinput15 spine_iw[19] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
X_0670_ col\[1\].zbuf_top_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[67] sky130_fd_sc_hd__buf_2
Xinput59 um_ow[121] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput48 um_ow[111] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[0\].zbuf_top_iw_I\[15\].genblk1.cell0_I net499 net435 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0937_ col\[0\].zbuf_top_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[30] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0868_ col\[7\].zbuf_bot_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[265] sky130_fd_sc_hd__buf_2
XFILLER_0_3_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0799_ col\[5\].zbuf_bot_iw_I\[16\].z vssd1 vssd1 vccd1 vccd1 um_iw[196] sky130_fd_sc_hd__buf_2
XFILLER_0_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput408 um_ow[90] vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[4\].zbuf_bot_iw_I\[17\].genblk1.cell0_I net495 net443 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_bot_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_2675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0722_ col\[3\].zbuf_bot_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[119] sky130_fd_sc_hd__buf_2
X_0653_ col\[1\].zbuf_bot_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[50] sky130_fd_sc_hd__buf_2
XFILLER_0_0_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0584_ _0154_ vssd1 vssd1 vccd1 vccd1 col\[2\].zbuf_top_ena_I.e sky130_fd_sc_hd__clkbuf_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[13\].genblk1.cell1_I zbuf_bus_iw_I\[13\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[13\].a sky130_fd_sc_hd__buf_6
XFILLER_0_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput227 um_ow[273] vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput216 um_ow[263] vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput205 um_ow[253] vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput238 um_ow[283] vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_2
Xinput249 um_ow[293] vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_1
Xcol\[2\].zbuf_top_iw_I\[14\].genblk1.cell0_I net501 net429 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_10_2725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_2572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_2748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_2603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0705_ col\[2\].zbuf_top_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[102] sky130_fd_sc_hd__buf_2
XFILLER_0_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0567_ _0143_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__clkbuf_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0498_ _0116_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[6\].zbuf_bot_iw_I\[16\].genblk1.cell0_I net498 net450 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_bot_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[0\].genblk1.cell1_I zbuf_bus_iw_I\[0\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[0\].a sky130_fd_sc_hd__buf_6
XFILLER_0_3_2601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[2\].zbuf_bot_iw_I\[7\].genblk1.cell0_I net481 net445 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_bot_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0421_ _0072_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__clkbuf_1
X_0352_ _0023_ _0024_ _0025_ _0026_ vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_2400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[4\].zbuf_bot_iw_I\[2\].genblk1.cell0_I net491 net444 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_bot_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_15_1732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_2177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[4\].zbuf_top_iw_I\[13\].genblk1.cell0_I net503 net423 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_118 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_129 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_2910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].genblk1.mux4_I\[13\].cell0_I net79 net345 net376 net402 net465 net452 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[13\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_9_2854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[0\].zbuf_top_iw_I\[6\].genblk1.cell0_I net483 net436 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[6\].z sky130_fd_sc_hd__and2_1
XTAP_36 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_47 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_58 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_69 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_2617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0970_ bus_ow\[23\] _0190_ vssd1 vssd1 vccd1 vccd1 spine_ow[24] sky130_fd_sc_hd__ebufn_8
XFILLER_0_3_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0404_ _0063_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__clkbuf_1
X_0335_ _0022_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__clkbuf_1
Xcol\[2\].zbuf_top_iw_I\[1\].genblk1.cell0_I net493 net430 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout511 col\[0\].zbuf_bot_iw_I\[0\].a vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__buf_6
Xfanout500 col\[0\].zbuf_bot_iw_I\[15\].a vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[6\].zbuf_top_iw_I\[12\].genblk1.cell0_I net506 net441 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_18 col\[0\].zbuf_bot_iw_I\[6\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_29 zbuf_bus_ena_I.z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0953_ bus_ow\[6\] _0173_ vssd1 vssd1 vccd1 vccd1 spine_ow[7] sky130_fd_sc_hd__ebufn_8
Xcol\[2\].genblk1.mux4_I\[23\].cell0_I net56 net83 net109 net136 net467 net456 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[23\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0884_ col\[7\].zbuf_top_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[281] sky130_fd_sc_hd__buf_2
XFILLER_0_10_2193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_bot_iw_I\[5\].genblk1.cell0_I net486 net440 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_bot_iw_I\[5\].z sky130_fd_sc_hd__and2_1
X_0318_ _0002_ _0006_ _0009_ _0013_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_2025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.mux4_I\[0\].cell0_I net243 net271 net297 net324 net473 net460 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[0\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_15_2071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_2813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput16 spine_iw[1] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput27 spine_iw[2] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
Xinput38 um_ow[102] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput49 um_ow[112] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__dlymetal6s2s_1
Xcol\[3\].zbuf_top_iw_I\[9\].genblk1.cell0_I net477 net425 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0936_ col\[0\].zbuf_top_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[29] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0867_ col\[7\].zbuf_bot_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[264] sky130_fd_sc_hd__buf_2
XFILLER_0_3_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0798_ col\[5\].zbuf_bot_iw_I\[15\].z vssd1 vssd1 vccd1 vccd1 um_iw[195] sky130_fd_sc_hd__buf_2
XFILLER_0_3_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput409 um_ow[91] vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[5\].zbuf_top_iw_I\[4\].genblk1.cell0_I net488 net420 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0721_ col\[3\].zbuf_bot_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[118] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0652_ col\[1\].zbuf_bot_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[49] sky130_fd_sc_hd__buf_2
XFILLER_0_12_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0583_ _0145_ _0153_ _0147_ _0148_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__and4b_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_2153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1066_ col\[6\].genblk1.mux4_I\[23\].x _0286_ vssd1 vssd1 vccd1 vccd1 bus_ow\[23\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_1_2017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0919_ col\[0\].zbuf_bot_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[12] sky130_fd_sc_hd__buf_2
XFILLER_0_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput217 um_ow[264] vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput206 um_ow[254] vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput239 um_ow[284] vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_2
Xinput228 um_ow[274] vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_2838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_2737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_2748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_2659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].genblk1.mux4_I\[10\].cell0_I net254 net282 net308 net335 net474 net461 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[10\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_6_2484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_2348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0704_ col\[2\].zbuf_top_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[101] sky130_fd_sc_hd__buf_2
XFILLER_0_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0566_ _0042_ _0044_ _0066_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__or3_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0497_ _0111_ _0108_ _0109_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__or3b_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[1\].zbuf_bot_iw_I\[16\].genblk1.cell0_I net497 net433 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_bot_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_7_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1049_ col\[6\].genblk1.mux4_I\[6\].x _0269_ vssd1 vssd1 vccd1 vccd1 bus_ow\[6\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_7_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[4\].genblk1.mux4_I\[1\].cell0_I net138 net165 net192 net218 net472 net459 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[1\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_10_1833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0420_ _0042_ _0044_ _0066_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__or3_1
X_0351_ _0032_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__clkbuf_1
Xcol\[1\].zbuf_top_ena_I.genblk1.cell0_I net539 net432 vssd1 vssd1 vccd1 vccd1 col\[1\].zbuf_top_ena_I.z
+ sky130_fd_sc_hd__and2_1
XFILLER_0_8_1801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0549_ _0137_ _0138_ _0139_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__nand3b_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_119 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_108 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_37 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_48 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_59 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[0\].genblk1.mux4_I\[17\].cell0_I net123 net354 net380 net406 net464 net451 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[17\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_12_2629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[3\].zbuf_bot_iw_I\[15\].genblk1.cell0_I net499 net427 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_bot_iw_I\[15\].z sky130_fd_sc_hd__and2_1
X_0403_ _0058_ _0059_ _0053_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__or3_1
X_0334_ _0002_ _0006_ _0009_ _0013_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_2253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout512 col\[0\].zbuf_bot_iw_I\[0\].a vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_4
Xfanout501 col\[0\].zbuf_bot_iw_I\[14\].a vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__buf_6
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[1\].zbuf_top_iw_I\[12\].genblk1.cell0_I net505 net431 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_sel_I\[2\].genblk1.cell1_I zbuf_bus_sel_I\[2\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 zbuf_bus_sel_I\[2\].z sky130_fd_sc_hd__buf_8
XFILLER_0_9_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_19 col\[0\].zbuf_bot_iw_I\[7\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0952_ bus_ow\[5\] _0172_ vssd1 vssd1 vccd1 vccd1 spine_ow[6] sky130_fd_sc_hd__ebufn_8
XFILLER_0_7_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0883_ col\[7\].zbuf_top_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[280] sky130_fd_sc_hd__buf_2
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0317_ _0002_ _0006_ _0009_ _0013_ vssd1 vssd1 vccd1 vccd1 zbuf_bus_ena_I.e sky130_fd_sc_hd__nor4_1
XFILLER_0_4_2037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].genblk1.mux4_I\[4\].cell0_I net248 net275 net302 net328 net473 net461 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[4\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_15_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[5\].zbuf_bot_iw_I\[14\].genblk1.cell0_I net502 net421 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_bot_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_2825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_2713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput17 spine_iw[20] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
Xinput28 spine_iw[3] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
Xinput39 um_ow[103] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_11_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_2267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0935_ col\[0\].zbuf_top_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[28] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0866_ col\[7\].zbuf_bot_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[263] sky130_fd_sc_hd__buf_2
Xcol\[2\].genblk1.mux4_I\[2\].cell0_I net416 net60 net86 net113 net469 net455 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[2\].x sky130_fd_sc_hd__mux4_1
Xcol\[3\].zbuf_top_iw_I\[11\].genblk1.cell0_I net507 net425 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[11\].z sky130_fd_sc_hd__and2_1
X_0797_ col\[5\].zbuf_bot_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[194] sky130_fd_sc_hd__buf_2
XFILLER_0_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[1\].zbuf_bot_iw_I\[7\].genblk1.cell0_I net481 net434 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_bot_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_1409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[3\].zbuf_bot_iw_I\[2\].genblk1.cell0_I net491 net428 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_bot_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0720_ col\[3\].zbuf_bot_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[117] sky130_fd_sc_hd__buf_2
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0651_ col\[1\].zbuf_bot_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[48] sky130_fd_sc_hd__buf_2
XFILLER_0_0_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0582_ _0216_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__inv_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[7\].zbuf_bot_iw_I\[13\].genblk1.cell0_I net504 net439 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_bot_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_2121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1065_ col\[6\].genblk1.mux4_I\[22\].x _0285_ vssd1 vssd1 vccd1 vccd1 bus_ow\[22\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_5_2165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0918_ col\[0\].zbuf_bot_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[11] sky130_fd_sc_hd__buf_2
X_0849_ col\[6\].zbuf_top_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[246] sky130_fd_sc_hd__buf_2
XFILLER_0_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput218 um_ow[265] vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_1
Xinput207 um_ow[255] vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput229 um_ow[275] vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_7_2920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[6\].zbuf_bot_ena_I.genblk1.cell0_I net548 net450 vssd1 vssd1 vccd1 vccd1 col\[6\].zbuf_bot_ena_I.z
+ sky130_fd_sc_hd__and2_1
XFILLER_0_14_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[5\].zbuf_top_iw_I\[10\].genblk1.cell0_I net510 net419 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[10\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_iw_I\[1\].genblk1.cell0_I net493 net432 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.mux4_I\[14\].cell0_I net260 net286 net313 net339 net474 net461 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[14\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_0_2073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0703_ col\[2\].zbuf_top_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[100] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0565_ _0142_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__clkbuf_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0496_ _0115_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__clkbuf_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xzbuf_bus_iw_I\[8\].genblk1.cell1_I zbuf_bus_iw_I\[8\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[8\].a sky130_fd_sc_hd__buf_6
XFILLER_0_7_2238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1048_ col\[6\].genblk1.mux4_I\[5\].x _0268_ vssd1 vssd1 vccd1 vccd1 bus_ow\[5\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[5\].cell0_I net142 net170 net196 net222 net472 net459 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[5\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_10_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0350_ _0023_ _0024_ _0025_ _0026_ vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__or4_1
Xcol\[6\].zbuf_bot_iw_I\[5\].genblk1.cell0_I net486 net449 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_bot_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_2157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_2168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0548_ _0137_ _0138_ _0139_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__nand3b_2
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0479_ _0105_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__clkbuf_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_2934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].genblk1.mux4_I\[3\].cell0_I net352 net234 net365 net391 net466 net453 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[3\].x sky130_fd_sc_hd__mux4_2
Xcol\[2\].zbuf_top_iw_I\[9\].genblk1.cell0_I net477 net429 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_38 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_49 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_2444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[4\].zbuf_top_iw_I\[4\].genblk1.cell0_I net487 net424 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[4\].z sky130_fd_sc_hd__and2_1
X_0402_ _0062_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__clkbuf_1
X_0333_ _0021_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__clkbuf_1
Xinput390 um_ow[74] vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout502 col\[0\].zbuf_bot_iw_I\[14\].a vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__clkbuf_4
Xfanout513 net514 vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_2617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xzbuf_bus_iw_I\[17\].genblk1.cell0_I net26 net513 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[17\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_0_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0951_ bus_ow\[4\] _0171_ vssd1 vssd1 vccd1 vccd1 spine_ow[5] sky130_fd_sc_hd__ebufn_8
XFILLER_0_12_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0882_ col\[7\].zbuf_top_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[279] sky130_fd_sc_hd__buf_2
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0316_ _0012_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_15_2073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[0\].zbuf_bot_iw_I\[14\].genblk1.cell0_I net501 net447 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_bot_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_11_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].genblk1.mux4_I\[8\].cell0_I net252 net280 net306 net332 net473 net460 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[8\].x sky130_fd_sc_hd__mux4_1
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_2725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_2414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_2561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput18 spine_iw[21] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput29 spine_iw[4] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
Xzbuf_bus_iw_I\[4\].genblk1.cell0_I net12 net514 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[4\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_9_1793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0934_ col\[0\].zbuf_top_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[27] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0865_ col\[7\].zbuf_bot_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[262] sky130_fd_sc_hd__buf_2
XFILLER_0_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[7\].zbuf_top_iw_I\[7\].genblk1.cell0_I net482 net438 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[7\].z sky130_fd_sc_hd__and2_1
X_0796_ col\[5\].zbuf_bot_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[193] sky130_fd_sc_hd__buf_2
Xcol\[2\].genblk1.mux4_I\[6\].cell0_I net38 net64 net91 net117 net469 net455 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[6\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_1_2712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_2909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0650_ col\[1\].zbuf_bot_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[47] sky130_fd_sc_hd__buf_2
XFILLER_0_0_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[2\].zbuf_bot_iw_I\[13\].genblk1.cell0_I net503 net445 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_bot_iw_I\[13\].z sky130_fd_sc_hd__and2_1
X_0581_ _0152_ vssd1 vssd1 vccd1 vccd1 col\[2\].zbuf_bot_ena_I.e sky130_fd_sc_hd__inv_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1064_ col\[6\].genblk1.mux4_I\[21\].x _0284_ vssd1 vssd1 vccd1 vccd1 bus_ow\[21\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_5_2177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0917_ col\[0\].zbuf_bot_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[10] sky130_fd_sc_hd__buf_2
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0848_ col\[6\].zbuf_top_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[245] sky130_fd_sc_hd__buf_2
XFILLER_0_12_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0779_ col\[4\].zbuf_top_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[176] sky130_fd_sc_hd__buf_2
Xinput208 um_ow[256] vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput219 um_ow[266] vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_10_2717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].zbuf_top_iw_I\[10\].genblk1.cell0_I net509 net435 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_2729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0702_ col\[2\].zbuf_top_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[99] sky130_fd_sc_hd__buf_2
Xcol\[6\].genblk1.mux4_I\[18\].cell0_I net264 net291 net317 net343 net475 net462 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[18\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0564_ _0043_ _0046_ _0097_ vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__or3b_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0495_ _0111_ _0108_ _0109_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__or3b_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1047_ col\[6\].genblk1.mux4_I\[4\].x _0267_ vssd1 vssd1 vccd1 vccd1 bus_ow\[4\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_14_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_2862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_bot_iw_I\[12\].genblk1.cell0_I net505 net443 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_bot_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[9\].cell0_I net148 net174 net200 net227 net471 net458 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[9\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_15_2425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0547_ _0137_ _0138_ _0139_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__nand3b_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0478_ zbuf_bus_sel_I\[4\].z zbuf_bus_sel_I\[2\].z zbuf_bus_sel_I\[3\].z vssd1 vssd1
+ vccd1 vccd1 _0105_ sky130_fd_sc_hd__or3b_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].genblk1.mux4_I\[7\].cell0_I net396 net279 net369 net395 net465 net452 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[7\].x sky130_fd_sc_hd__mux4_2
XTAP_39 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_2480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_2377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0401_ _0058_ _0059_ _0053_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__or3_1
X_0332_ _0002_ _0006_ _0009_ _0013_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__or4_1
Xinput380 um_ow[65] vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__clkbuf_1
Xinput391 um_ow[75] vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_2211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[0\].zbuf_bot_iw_I\[7\].genblk1.cell0_I net481 net447 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_bot_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_2288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].zbuf_bot_iw_I\[11\].genblk1.cell0_I net508 net450 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_bot_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout503 col\[0\].zbuf_bot_iw_I\[13\].a vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__buf_6
Xfanout514 net515 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__clkbuf_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_2109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].zbuf_bot_iw_I\[2\].genblk1.cell0_I net491 net446 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_bot_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_2710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_2631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_2253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0950_ bus_ow\[3\] _0170_ vssd1 vssd1 vccd1 vccd1 spine_ow[4] sky130_fd_sc_hd__ebufn_8
XFILLER_0_3_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0881_ col\[7\].zbuf_top_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[278] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0315_ net2 _0000_ _0010_ net7 _0011_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__a221o_2
XFILLER_0_8_1485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_top_iw_I\[1\].genblk1.cell0_I net493 net436 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[1\].z sky130_fd_sc_hd__and2_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_2737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_2573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput19 spine_iw[22] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_2326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0933_ col\[0\].zbuf_top_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[26] sky130_fd_sc_hd__buf_2
X_0864_ col\[7\].zbuf_bot_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[261] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0795_ col\[5\].zbuf_bot_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[192] sky130_fd_sc_hd__buf_2
XFILLER_0_5_2871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[5\].zbuf_bot_iw_I\[5\].genblk1.cell0_I net486 net422 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_bot_iw_I\[5\].z sky130_fd_sc_hd__and2_1
Xcol\[2\].genblk1.mux4_I\[13\].cell0_I net45 net72 net98 net125 net467 net454 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[13\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_6_1901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0580_ net468 net455 _0216_ zbuf_bus_ena_I.z vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__or4b_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[7\].zbuf_bot_iw_I\[0\].genblk1.cell0_I net512 net440 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_bot_iw_I\[0\].z sky130_fd_sc_hd__and2_1
X_1063_ col\[6\].genblk1.mux4_I\[20\].x _0283_ vssd1 vssd1 vccd1 vccd1 bus_ow\[20\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_5_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0916_ col\[0\].zbuf_bot_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[9] sky130_fd_sc_hd__buf_2
XFILLER_0_12_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0847_ col\[6\].zbuf_top_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[244] sky130_fd_sc_hd__buf_2
XFILLER_0_3_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0778_ col\[4\].zbuf_top_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[175] sky130_fd_sc_hd__buf_2
Xinput209 um_ow[257] vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__dlymetal6s2s_1
Xcol\[1\].zbuf_top_iw_I\[9\].genblk1.cell0_I net477 net431 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[9\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_2521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[3\].zbuf_top_iw_I\[4\].genblk1.cell0_I net487 net426 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_2353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[23\].cell0_I net163 net189 net216 net242 net471 net458 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[23\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_13_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0701_ col\[2\].zbuf_top_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[98] sky130_fd_sc_hd__buf_2
XFILLER_0_13_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0563_ _0141_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0494_ _0114_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__clkbuf_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_2117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1046_ col\[6\].genblk1.mux4_I\[3\].x _0266_ vssd1 vssd1 vccd1 vccd1 bus_ow\[3\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_2351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_2505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_top_iw_I\[17\].genblk1.cell0_I net496 net437 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_15_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_2295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0546_ _0047_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__clkbuf_4
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0477_ _0104_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__clkbuf_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_2903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1029_ col\[4\].genblk1.mux4_I\[10\].x _0249_ vssd1 vssd1 vccd1 vccd1 bus_ow\[10\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_7_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_2824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[6\].zbuf_top_iw_I\[7\].genblk1.cell0_I net482 net442 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0400_ _0061_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__clkbuf_1
X_0331_ _0020_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__clkbuf_1
Xcol\[1\].zbuf_bot_iw_I\[11\].genblk1.cell0_I net507 net433 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_bot_iw_I\[11\].z sky130_fd_sc_hd__and2_1
Xinput381 um_ow[66] vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__clkbuf_1
Xinput370 um_ow[56] vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__clkbuf_1
Xinput392 um_ow[76] vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_2234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_2368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout504 col\[0\].zbuf_bot_iw_I\[13\].a vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout515 net516 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__clkbuf_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0529_ _0133_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__clkbuf_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_2490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0880_ col\[7\].zbuf_top_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[277] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0314_ net4 net6 vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_2928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_2806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_2541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_2405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[3\].zbuf_bot_iw_I\[10\].genblk1.cell0_I net509 net427 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_bot_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_4_2585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_2338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0932_ col\[0\].zbuf_top_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[25] sky130_fd_sc_hd__buf_2
X_0863_ col\[7\].zbuf_bot_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[260] sky130_fd_sc_hd__buf_2
X_0794_ col\[5\].zbuf_bot_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[191] sky130_fd_sc_hd__buf_2
XFILLER_0_12_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_2894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[2\].genblk1.mux4_I\[17\].cell0_I net50 net76 net103 net129 net467 net456 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[17\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_6_2603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_2658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_2246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1062_ col\[6\].genblk1.mux4_I\[19\].x _0282_ vssd1 vssd1 vccd1 vccd1 bus_ow\[19\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_5_1401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0915_ col\[0\].zbuf_bot_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[8] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0846_ col\[6\].zbuf_top_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[243] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0777_ col\[4\].zbuf_top_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[174] sky130_fd_sc_hd__buf_2
XFILLER_0_3_2809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0700_ col\[2\].zbuf_top_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[97] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0562_ _0124_ _0045_ _0076_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__or3b_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0493_ _0111_ _0108_ _0109_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__or3b_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[1\].zbuf_bot_iw_I\[2\].genblk1.cell0_I net491 net434 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_bot_iw_I\[2\].z sky130_fd_sc_hd__and2_1
X_1045_ col\[6\].genblk1.mux4_I\[2\].x _0265_ vssd1 vssd1 vccd1 vccd1 bus_ow\[2\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_14_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0829_ col\[6\].zbuf_bot_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[226] sky130_fd_sc_hd__buf_2
Xzbuf_bus_iw_I\[16\].genblk1.cell1_I zbuf_bus_iw_I\[16\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[16\].a sky130_fd_sc_hd__buf_6
XFILLER_0_7_2720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_2742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_2505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].zbuf_top_iw_I\[17\].genblk1.cell0_I net495 net429 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_8_2517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_2263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0545_ _0077_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__clkbuf_4
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0476_ _0096_ _0046_ _0097_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__or3b_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1028_ col\[4\].genblk1.mux4_I\[9\].x _0248_ vssd1 vssd1 vccd1 vccd1 bus_ow\[9\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_8_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[2\].zbuf_bot_ena_I.genblk1.cell0_I net540 net446 vssd1 vssd1 vccd1 vccd1 col\[2\].zbuf_bot_ena_I.z
+ sky130_fd_sc_hd__and2_1
XFILLER_0_14_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xzbuf_bus_iw_I\[3\].genblk1.cell1_I zbuf_bus_iw_I\[3\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[3\].a sky130_fd_sc_hd__buf_6
X_0330_ _0002_ _0006_ _0009_ _0013_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__or4_1
Xinput360 um_ow[47] vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__clkbuf_2
Xinput371 um_ow[57] vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_1
Xinput393 um_ow[77] vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__clkbuf_1
Xinput382 um_ow[67] vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_2358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout505 col\[0\].zbuf_bot_iw_I\[12\].a vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__buf_6
XFILLER_0_1_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_bot_iw_I\[5\].genblk1.cell0_I net485 net444 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_bot_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0528_ _0124_ _0121_ _0122_ vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__or3b_1
Xfanout516 zbuf_bus_ena_I.e vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0459_ _0094_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__clkbuf_1
Xcol\[4\].zbuf_top_iw_I\[16\].genblk1.cell0_I net497 net423 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[6\].zbuf_bot_iw_I\[0\].genblk1.cell0_I net512 net449 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_bot_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_top_iw_I\[9\].genblk1.cell0_I net477 net435 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[9\].z sky130_fd_sc_hd__and2_1
X_0313_ net5 vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__inv_2
Xinput190 um_ow[23] vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_8_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_2043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[2\].zbuf_top_iw_I\[4\].genblk1.cell0_I net487 net430 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_2829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_2597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0931_ col\[0\].zbuf_top_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[24] sky130_fd_sc_hd__buf_2
XFILLER_0_3_2085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].zbuf_top_iw_I\[15\].genblk1.cell0_I net500 net441 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[15\].z sky130_fd_sc_hd__and2_1
X_0862_ col\[7\].zbuf_bot_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[259] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0793_ col\[5\].zbuf_bot_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[190] sky130_fd_sc_hd__buf_2
XFILLER_0_3_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xzbuf_bus_iw_I\[12\].genblk1.cell0_I net21 net515 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[12\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_8_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[7\].zbuf_bot_iw_I\[8\].genblk1.cell0_I net480 net439 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_bot_iw_I\[8\].z sky130_fd_sc_hd__and2_1
Xcol\[0\].genblk1.mux4_I\[22\].cell0_I net179 net359 net386 net412 net464 net451 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[22\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_6_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_2350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1061_ col\[6\].genblk1.mux4_I\[18\].x _0281_ vssd1 vssd1 vccd1 vccd1 bus_ow\[18\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_9_2272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0914_ col\[0\].zbuf_bot_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[7] sky130_fd_sc_hd__buf_2
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0845_ col\[6\].zbuf_top_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[242] sky130_fd_sc_hd__buf_2
XFILLER_0_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0776_ col\[4\].zbuf_top_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[173] sky130_fd_sc_hd__buf_2
XFILLER_0_3_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_2913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[5\].zbuf_top_iw_I\[7\].genblk1.cell0_I net482 net420 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[6\].zbuf_top_ena_I.genblk1.cell0_I net549 net441 vssd1 vssd1 vccd1 vccd1 col\[6\].zbuf_top_ena_I.z
+ sky130_fd_sc_hd__and2_1
XFILLER_0_6_2412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[7\].zbuf_top_iw_I\[2\].genblk1.cell0_I net492 net438 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_2099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[0\].zbuf_bot_ena_I.genblk1.cell0_I_536 vssd1 vssd1 vccd1 vccd1 net536 col\[0\].zbuf_bot_ena_I.genblk1.cell0_I_536/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_1_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0561_ _0075_ _0077_ _0047_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__nand3b_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0492_ _0113_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__clkbuf_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1044_ col\[6\].genblk1.mux4_I\[1\].x _0264_ vssd1 vssd1 vccd1 vccd1 bus_ow\[1\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_0_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0828_ col\[6\].zbuf_bot_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[225] sky130_fd_sc_hd__buf_2
XFILLER_0_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0759_ col\[4\].zbuf_bot_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[156] sky130_fd_sc_hd__buf_2
XFILLER_0_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_2620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_2529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0544_ _0075_ vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__clkbuf_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0475_ _0103_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__clkbuf_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1027_ col\[4\].genblk1.mux4_I\[8\].x _0247_ vssd1 vssd1 vccd1 vccd1 bus_ow\[8\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_5_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_2827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput350 um_ow[38] vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__clkbuf_2
Xinput372 um_ow[58] vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__clkbuf_1
Xinput361 um_ow[48] vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__clkbuf_1
Xinput394 um_ow[78] vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__clkbuf_1
Xinput383 um_ow[68] vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_2892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[1\].zbuf_bot_ena_I.genblk1.cell0_I_538 vssd1 vssd1 vccd1 vccd1 net538 col\[1\].zbuf_bot_ena_I.genblk1.cell0_I_538/LO
+ sky130_fd_sc_hd__conb_1
Xfanout506 col\[0\].zbuf_bot_iw_I\[12\].a vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__clkbuf_4
X_0527_ _0132_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__clkbuf_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0458_ _0083_ _0089_ _0084_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__or3b_1
X_0389_ _0043_ _0045_ _0053_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__or3_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_2601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0312_ _0008_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__clkbuf_2
Xinput180 um_ow[230] vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_2101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput191 um_ow[240] vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_15_2099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_bot_iw_I\[2\].genblk1.cell0_I net491 net448 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_bot_iw_I\[2\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_iw_I\[15\].genblk1.cell0_I net499 net431 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[15\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0930_ col\[0\].zbuf_top_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[23] sky130_fd_sc_hd__buf_2
XFILLER_0_3_2053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_2097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0861_ col\[7\].zbuf_bot_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[258] sky130_fd_sc_hd__buf_2
X_0792_ col\[5\].zbuf_bot_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[189] sky130_fd_sc_hd__buf_2
XFILLER_0_12_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_2773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_2226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[5\].zbuf_bot_iw_I\[17\].genblk1.cell0_I net496 net421 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_bot_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1060_ col\[6\].genblk1.mux4_I\[17\].x _0280_ vssd1 vssd1 vccd1 vccd1 bus_ow\[17\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_9_2284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_2025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_2069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0913_ col\[0\].zbuf_bot_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[6] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0844_ col\[6\].zbuf_top_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[241] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0775_ col\[4\].zbuf_top_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[172] sky130_fd_sc_hd__buf_2
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[3\].zbuf_top_iw_I\[14\].genblk1.cell0_I net501 net425 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_2546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_2345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_2389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_2181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0560_ _0140_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0491_ _0111_ _0108_ _0109_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__or3b_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[3\].zbuf_bot_iw_I\[5\].genblk1.cell0_I net485 net428 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_bot_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1043_ col\[6\].genblk1.mux4_I\[0\].x _0263_ vssd1 vssd1 vccd1 vccd1 bus_ow\[0\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_14_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_2890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0827_ col\[6\].zbuf_bot_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[224] sky130_fd_sc_hd__buf_2
X_0758_ col\[4\].zbuf_bot_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[155] sky130_fd_sc_hd__buf_2
Xcol\[5\].zbuf_bot_iw_I\[0\].genblk1.cell0_I net512 net422 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_bot_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0689_ col\[2\].zbuf_bot_iw_I\[14\].z vssd1 vssd1 vccd1 vccd1 um_iw[86] sky130_fd_sc_hd__buf_2
Xcol\[7\].zbuf_bot_iw_I\[16\].genblk1.cell0_I net498 net439 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_bot_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_2654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_2632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[5\].zbuf_top_iw_I\[13\].genblk1.cell0_I net504 net419 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[13\].z sky130_fd_sc_hd__and2_1
Xcol\[1\].zbuf_top_iw_I\[4\].genblk1.cell0_I net487 net432 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[4\].z sky130_fd_sc_hd__and2_1
X_0543_ _0134_ _0135_ _0136_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__nand3b_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0474_ _0096_ _0046_ _0097_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__or3b_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1026_ col\[4\].genblk1.mux4_I\[7\].x _0246_ vssd1 vssd1 vccd1 vccd1 bus_ow\[7\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[13\].cell0_I net152 net178 net205 net231 net470 net457 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[13\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_14_2462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_2337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xzbuf_bus_sel_I\[1\].genblk1.cell0_I net27 net516 vssd1 vssd1 vccd1 vccd1 zbuf_bus_sel_I\[1\].genblk1.l
+ sky130_fd_sc_hd__and2_1
Xinput340 um_ow[375] vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput351 um_ow[39] vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_2
Xinput362 um_ow[49] vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_1
Xinput395 um_ow[79] vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__clkbuf_1
Xinput384 um_ow[69] vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__clkbuf_1
Xinput373 um_ow[59] vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_2316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_2338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].zbuf_bot_iw_I\[8\].genblk1.cell0_I net480 net449 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_bot_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout507 col\[0\].zbuf_bot_iw_I\[11\].a vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__buf_6
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0526_ _0124_ _0121_ _0122_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__or3b_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0457_ _0093_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__clkbuf_1
X_0388_ _0054_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_2872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_2883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1009_ col\[2\].genblk1.mux4_I\[14\].x _0229_ vssd1 vssd1 vccd1 vccd1 bus_ow\[14\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_4_2747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_2613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[7\].zbuf_top_iw_I\[12\].genblk1.cell0_I net506 net437 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[12\].z sky130_fd_sc_hd__and2_1
Xcol\[2\].zbuf_top_ena_I.genblk1.cell0_I_541 vssd1 vssd1 vccd1 vccd1 net541 col\[2\].zbuf_top_ena_I.genblk1.cell0_I_541/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_9_2625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[6\].genblk1.mux4_I\[23\].cell0_I net270 net296 net322 net349 net475 net462 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[23\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_9_2669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_2235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0311_ _0003_ net34 net1 _0004_ _0007_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__o221ai_4
Xinput170 um_ow[221] vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_1
Xinput181 um_ow[231] vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_2113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput192 um_ow[241] vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_2001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_2909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_top_iw_I\[7\].genblk1.cell0_I net481 net424 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0509_ _0111_ _0121_ _0122_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__or3b_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[6\].zbuf_top_iw_I\[2\].genblk1.cell0_I net492 net442 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_11_1775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0860_ col\[7\].zbuf_bot_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[257] sky130_fd_sc_hd__buf_2
X_0791_ col\[5\].zbuf_bot_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[188] sky130_fd_sc_hd__buf_2
XFILLER_0_11_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_2741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0989_ col\[0\].genblk1.mux4_I\[18\].x _0209_ vssd1 vssd1 vccd1 vccd1 bus_ow\[18\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].zbuf_bot_iw_I\[17\].genblk1.cell0_I net495 net448 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_bot_iw_I\[17\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_2617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_2538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[3\].zbuf_top_ena_I.genblk1.cell0_I_543 vssd1 vssd1 vccd1 vccd1 net543 col\[3\].zbuf_top_ena_I.genblk1.cell0_I_543/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_9_2241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_2127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0912_ col\[0\].zbuf_bot_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[5] sky130_fd_sc_hd__buf_2
X_0843_ col\[6\].zbuf_top_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[240] sky130_fd_sc_hd__buf_2
XFILLER_0_4_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0774_ col\[4\].zbuf_top_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[171] sky130_fd_sc_hd__buf_2
Xzbuf_bus_iw_I\[7\].genblk1.cell0_I net15 net513 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[7\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_12_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_2193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_2035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_2068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0490_ _0112_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__clkbuf_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1042_ col\[4\].genblk1.mux4_I\[23\].x _0262_ vssd1 vssd1 vccd1 vccd1 bus_ow\[23\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_9_2071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_2856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].zbuf_bot_iw_I\[16\].genblk1.cell0_I net497 net445 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_bot_iw_I\[16\].z sky130_fd_sc_hd__and2_1
XFILLER_0_12_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0826_ col\[6\].zbuf_bot_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[223] sky130_fd_sc_hd__buf_2
X_0757_ col\[4\].zbuf_bot_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[154] sky130_fd_sc_hd__buf_2
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0688_ col\[2\].zbuf_bot_iw_I\[13\].z vssd1 vssd1 vccd1 vccd1 um_iw[85] sky130_fd_sc_hd__buf_2
XFILLER_0_7_2712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_2745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_2644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[0\].zbuf_top_iw_I\[13\].genblk1.cell0_I net503 net435 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0542_ _0134_ _0135_ _0136_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__nand3b_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0473_ _0102_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__clkbuf_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[4\].zbuf_top_ena_I.genblk1.cell0_I_545 vssd1 vssd1 vccd1 vccd1 net545 col\[4\].zbuf_top_ena_I.genblk1.cell0_I_545/LO
+ sky130_fd_sc_hd__conb_1
X_1025_ col\[4\].genblk1.mux4_I\[6\].x _0245_ vssd1 vssd1 vccd1 vccd1 bus_ow\[6\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_11_2828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0809_ col\[5\].zbuf_top_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[206] sky130_fd_sc_hd__buf_2
XFILLER_0_13_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[17\].cell0_I net156 net183 net209 net236 net470 net457 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[17\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_9_2818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_2575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[4\].zbuf_bot_iw_I\[15\].genblk1.cell0_I net499 net443 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_bot_iw_I\[15\].z sky130_fd_sc_hd__and2_1
Xinput330 um_ow[366] vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput341 um_ow[376] vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__clkbuf_2
Xinput352 um_ow[3] vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput363 um_ow[4] vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput374 um_ow[5] vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput396 um_ow[7] vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__clkbuf_2
Xinput385 um_ow[6] vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_15_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _0150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout508 col\[0\].zbuf_bot_iw_I\[11\].a vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_4
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0525_ _0131_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__clkbuf_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0456_ _0083_ _0089_ _0084_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__or3b_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xzbuf_bus_iw_I\[11\].genblk1.cell1_I zbuf_bus_iw_I\[11\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[11\].a sky130_fd_sc_hd__buf_6
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0387_ _0043_ _0045_ _0053_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_2840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1008_ col\[2\].genblk1.mux4_I\[13\].x _0228_ vssd1 vssd1 vccd1 vccd1 bus_ow\[13\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_14_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].zbuf_top_iw_I\[12\].genblk1.cell0_I net505 net429 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_2157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0310_ net7 net5 vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__or2b_1
Xinput171 um_ow[222] vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_1
Xinput160 um_ow[212] vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_1
Xinput182 um_ow[232] vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_1
Xinput193 um_ow[242] vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_8_2125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_2169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_2057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_2934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0508_ _0046_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0439_ _0042_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__clkbuf_2
Xcol\[6\].zbuf_bot_iw_I\[14\].genblk1.cell0_I net502 net450 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_bot_iw_I\[14\].z sky130_fd_sc_hd__and2_1
Xcol\[5\].zbuf_top_ena_I.genblk1.cell0_I_547 vssd1 vssd1 vccd1 vccd1 net547 col\[5\].zbuf_top_ena_I.genblk1.cell0_I_547/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_0_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].zbuf_bot_iw_I\[5\].genblk1.cell0_I net485 net446 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_bot_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_2489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0790_ col\[5\].zbuf_bot_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[187] sky130_fd_sc_hd__buf_2
XFILLER_0_3_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_bot_iw_I\[0\].genblk1.cell0_I net511 net444 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_bot_iw_I\[0\].z sky130_fd_sc_hd__and2_1
XFILLER_0_11_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_top_iw_I\[11\].genblk1.cell0_I net507 net423 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_2843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_2753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0988_ col\[0\].genblk1.mux4_I\[17\].x _0208_ vssd1 vssd1 vccd1 vccd1 bus_ow\[17\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_6_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_2629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_2206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_2386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_2241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[0\].zbuf_top_iw_I\[4\].genblk1.cell0_I net487 net436 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_top_iw_I\[4\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0911_ col\[0\].zbuf_bot_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[4] sky130_fd_sc_hd__buf_2
X_0842_ col\[6\].zbuf_top_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[239] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0773_ col\[4\].zbuf_top_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[170] sky130_fd_sc_hd__buf_2
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_2826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_2437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[6\].zbuf_top_ena_I.genblk1.cell0_I_549 vssd1 vssd1 vccd1 vccd1 net549 col\[6\].zbuf_top_ena_I.genblk1.cell0_I_549/LO
+ sky130_fd_sc_hd__conb_1
Xcol\[6\].zbuf_top_iw_I\[10\].genblk1.cell0_I net510 net441 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_top_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[5\].zbuf_bot_iw_I\[8\].genblk1.cell0_I net480 net421 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_bot_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1041_ col\[4\].genblk1.mux4_I\[22\].x _0261_ vssd1 vssd1 vccd1 vccd1 bus_ow\[22\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xcol\[0\].genblk1.mux4_I\[12\].cell0_I net68 net334 net375 net401 net465 net452 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[12\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_13_2881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_bot_iw_I\[3\].genblk1.cell0_I net490 net440 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_bot_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0825_ col\[6\].zbuf_bot_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[222] sky130_fd_sc_hd__buf_2
XFILLER_0_3_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0756_ col\[4\].zbuf_bot_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[153] sky130_fd_sc_hd__buf_2
XFILLER_0_12_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0687_ col\[2\].zbuf_bot_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[84] sky130_fd_sc_hd__buf_2
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_2667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_2345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[3\].zbuf_top_iw_I\[7\].genblk1.cell0_I net481 net426 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_top_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0541_ _0134_ _0135_ _0136_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__nand3b_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0472_ _0096_ _0046_ _0097_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__or3b_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_2009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1024_ col\[4\].genblk1.mux4_I\[5\].x _0244_ vssd1 vssd1 vccd1 vccd1 bus_ow\[5\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[5\].zbuf_top_iw_I\[2\].genblk1.cell0_I net492 net420 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_top_iw_I\[2\].z sky130_fd_sc_hd__and2_1
XFILLER_0_2_1986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0808_ col\[5\].zbuf_top_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[205] sky130_fd_sc_hd__buf_2
XFILLER_0_4_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].genblk1.mux4_I\[22\].cell0_I net55 net82 net108 net135 net467 net456 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[22\].x sky130_fd_sc_hd__mux4_1
X_0739_ col\[3\].zbuf_top_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[136] sky130_fd_sc_hd__buf_2
XFILLER_0_7_2521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_2407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].zbuf_top_ena_I.genblk1.cell0_I net541 net430 vssd1 vssd1 vccd1 vccd1 col\[2\].zbuf_top_ena_I.z
+ sky130_fd_sc_hd__and2_1
Xinput320 um_ow[357] vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput353 um_ow[40] vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__clkbuf_2
Xinput331 um_ow[367] vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput342 um_ow[377] vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_2
Xinput397 um_ow[80] vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__clkbuf_1
Xinput386 um_ow[70] vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_1
Xinput375 um_ow[60] vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__clkbuf_1
Xinput364 um_ow[50] vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_2 bus_ow\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout509 col\[0\].zbuf_bot_iw_I\[10\].a vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__buf_8
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0524_ _0124_ _0121_ _0122_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__or3b_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0455_ _0092_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__clkbuf_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0386_ _0046_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__clkbuf_2
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_2863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1007_ col\[2\].genblk1.mux4_I\[12\].x _0227_ vssd1 vssd1 vccd1 vccd1 bus_ow\[12\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_8_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_2773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_2451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_2261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_2125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_2169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput172 um_ow[223] vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_1
Xinput150 um_ow[203] vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_1
Xinput161 um_ow[213] vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__clkbuf_1
Xinput183 um_ow[233] vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_1
Xinput194 um_ow[243] vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_8_2137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_2782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[1\].zbuf_bot_iw_I\[14\].genblk1.cell0_I net501 net433 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_bot_iw_I\[14\].z sky130_fd_sc_hd__and2_1
XFILLER_0_1_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0507_ zbuf_bus_sel_I\[2\].z vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__clkbuf_2
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0438_ _0082_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__clkbuf_1
X_0369_ _0041_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_1801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_2489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_2402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_2209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_2911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_2067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_2765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0987_ col\[0\].genblk1.mux4_I\[16\].x _0207_ vssd1 vssd1 vccd1 vccd1 bus_ow\[16\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_6_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_2297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[3\].zbuf_bot_iw_I\[13\].genblk1.cell0_I net503 net427 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_bot_iw_I\[13\].z sky130_fd_sc_hd__and2_1
XFILLER_0_9_2221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0910_ col\[0\].zbuf_bot_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[3] sky130_fd_sc_hd__buf_2
XFILLER_0_3_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0841_ col\[6\].zbuf_top_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[238] sky130_fd_sc_hd__buf_2
XFILLER_0_0_2785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0772_ col\[4\].zbuf_top_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[169] sky130_fd_sc_hd__buf_2
XFILLER_0_3_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xcol\[4\].genblk1.mux4_I\[0\].cell0_I net137 net164 net191 net217 net472 net459 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[0\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_12_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[1\].zbuf_top_iw_I\[10\].genblk1.cell0_I net509 net431 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_top_iw_I\[10\].z sky130_fd_sc_hd__and2_1
XFILLER_0_13_1625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xzbuf_bus_sel_I\[0\].genblk1.cell1_I zbuf_bus_sel_I\[0\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 zbuf_bus_sel_I\[0\].z sky130_fd_sc_hd__buf_6
XFILLER_0_11_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1040_ col\[4\].genblk1.mux4_I\[21\].x _0260_ vssd1 vssd1 vccd1 vccd1 bus_ow\[21\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_9_2051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_2073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_2836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[0\].genblk1.mux4_I\[16\].cell0_I net112 net353 net379 net405 net464 net451 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[16\].x sky130_fd_sc_hd__mux4_2
XFILLER_0_0_2593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0824_ col\[6\].zbuf_bot_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[221] sky130_fd_sc_hd__buf_2
XFILLER_0_4_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0755_ col\[4\].zbuf_bot_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[152] sky130_fd_sc_hd__buf_2
XFILLER_0_3_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0686_ col\[2\].zbuf_bot_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[83] sky130_fd_sc_hd__buf_2
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[7\].zbuf_bot_ena_I.genblk1.cell0_I net550 net440 vssd1 vssd1 vccd1 vccd1 col\[7\].zbuf_bot_ena_I.z
+ sky130_fd_sc_hd__and2_1
XFILLER_0_14_1912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[5\].zbuf_bot_iw_I\[12\].genblk1.cell0_I net506 net421 vssd1 vssd1 vccd1 vccd1
+ col\[5\].zbuf_bot_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_1989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_2381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_2213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_2167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0540_ _0134_ _0135_ _0136_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_0_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0471_ _0101_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1023_ col\[4\].genblk1.mux4_I\[4\].x _0243_ vssd1 vssd1 vccd1 vccd1 bus_ow\[4\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_2_2600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_2819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_2633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_2644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0807_ col\[5\].zbuf_top_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[204] sky130_fd_sc_hd__buf_2
XFILLER_0_4_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0738_ col\[3\].zbuf_top_iw_I\[9\].z vssd1 vssd1 vccd1 vccd1 um_iw[135] sky130_fd_sc_hd__buf_2
XFILLER_0_13_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[1\].zbuf_bot_iw_I\[5\].genblk1.cell0_I net485 net434 vssd1 vssd1 vccd1 vccd1
+ col\[1\].zbuf_bot_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0669_ col\[1\].zbuf_top_iw_I\[12\].z vssd1 vssd1 vccd1 vccd1 um_iw[66] sky130_fd_sc_hd__buf_2
XFILLER_0_0_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_2533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_2577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[3\].zbuf_bot_iw_I\[0\].genblk1.cell0_I net511 net428 vssd1 vssd1 vccd1 vccd1
+ col\[3\].zbuf_bot_iw_I\[0\].z sky130_fd_sc_hd__and2_1
Xcol\[6\].genblk1.mux4_I\[3\].cell0_I net247 net274 net300 net327 net473 net460 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[3\].x sky130_fd_sc_hd__mux4_1
Xinput310 um_ow[348] vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput321 um_ow[358] vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput332 um_ow[368] vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput343 um_ow[378] vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_2
Xinput354 um_ow[41] vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_2
Xinput387 um_ow[71] vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__clkbuf_1
Xinput376 um_ow[61] vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__clkbuf_1
Xinput365 um_ow[51] vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_1
Xinput398 um_ow[81] vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_2043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_2841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_3 col\[0\].zbuf_bot_iw_I\[12\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[7\].zbuf_bot_iw_I\[11\].genblk1.cell0_I net508 net439 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_bot_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_10_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0523_ _0130_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__clkbuf_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0454_ _0083_ _0089_ _0084_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__or3b_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0385_ _0052_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_2853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1006_ col\[2\].genblk1.mux4_I\[11\].x _0226_ vssd1 vssd1 vccd1 vccd1 bus_ow\[11\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_4_2717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_2739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_2897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_2796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_2785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[2\].genblk1.mux4_I\[1\].cell0_I net415 net59 net85 net111 net468 net454 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[1\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput151 um_ow[204] vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__clkbuf_1
Xinput162 um_ow[214] vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_1
Xinput140 um_ow[195] vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_1
Xinput173 um_ow[224] vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_1
Xinput184 um_ow[234] vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_1
Xinput195 um_ow[244] vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_8_2149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xzbuf_bus_iw_I\[6\].genblk1.cell1_I zbuf_bus_iw_I\[6\].genblk1.l vssd1 vssd1 vccd1
+ vccd1 col\[0\].zbuf_bot_iw_I\[6\].a sky130_fd_sc_hd__buf_6
XFILLER_0_14_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0506_ _0120_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__clkbuf_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0437_ _0075_ _0076_ _0077_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__or3b_1
X_0368_ zbuf_bus_sel_I\[4\].z zbuf_bus_sel_I\[2\].z zbuf_bus_sel_I\[3\].z vssd1 vssd1
+ vccd1 vccd1 _0041_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_2661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_2547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_2593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_bot_iw_I\[8\].genblk1.cell0_I net479 net443 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_bot_iw_I\[8\].z sky130_fd_sc_hd__and2_1
XFILLER_0_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xcol\[6\].zbuf_bot_iw_I\[3\].genblk1.cell0_I net490 net449 vssd1 vssd1 vccd1 vccd1
+ col\[6\].zbuf_bot_iw_I\[3\].z sky130_fd_sc_hd__and2_1
XFILLER_0_10_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_2878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0986_ col\[0\].genblk1.mux4_I\[15\].x _0206_ vssd1 vssd1 vccd1 vccd1 bus_ow\[15\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_14_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[6\].genblk1.mux4_I\[13\].cell0_I net259 net285 net311 net338 net474 net461 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[13\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_1_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_2508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_2491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_2265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[2\].zbuf_top_iw_I\[7\].genblk1.cell0_I net481 net430 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_top_iw_I\[7\].z sky130_fd_sc_hd__and2_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_2233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].zbuf_top_iw_I\[2\].genblk1.cell0_I net491 net424 vssd1 vssd1 vccd1 vccd1
+ col\[4\].zbuf_top_iw_I\[2\].z sky130_fd_sc_hd__and2_1
X_0840_ col\[6\].zbuf_top_iw_I\[3\].z vssd1 vssd1 vccd1 vccd1 um_iw[237] sky130_fd_sc_hd__buf_2
XFILLER_0_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_2797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0771_ col\[4\].zbuf_top_iw_I\[6\].z vssd1 vssd1 vccd1 vccd1 um_iw[168] sky130_fd_sc_hd__buf_2
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xcol\[4\].genblk1.mux4_I\[4\].cell0_I net141 net169 net195 net221 net472 net459 vssd1
+ vssd1 vccd1 vccd1 col\[4\].genblk1.mux4_I\[4\].x sky130_fd_sc_hd__mux4_1
XFILLER_0_7_2929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_2817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_2631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_2528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_2517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_2686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0969_ bus_ow\[22\] _0189_ vssd1 vssd1 vccd1 vccd1 spine_ow[23] sky130_fd_sc_hd__ebufn_8
XFILLER_0_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xzbuf_bus_iw_I\[15\].genblk1.cell0_I net24 net513 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[15\].genblk1.l
+ sky130_fd_sc_hd__and2_1
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_2073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[0\].genblk1.mux4_I\[2\].cell0_I net257 net223 net364 net390 net466 net453 vssd1
+ vssd1 vccd1 vccd1 col\[0\].genblk1.mux4_I\[2\].x sky130_fd_sc_hd__mux4_2
Xfanout490 col\[0\].zbuf_bot_iw_I\[3\].a vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_2085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_2894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0823_ col\[6\].zbuf_bot_iw_I\[4\].z vssd1 vssd1 vccd1 vccd1 um_iw[220] sky130_fd_sc_hd__buf_2
XFILLER_0_4_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0754_ col\[4\].zbuf_bot_iw_I\[7\].z vssd1 vssd1 vccd1 vccd1 um_iw[151] sky130_fd_sc_hd__buf_2
XFILLER_0_4_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0685_ col\[2\].zbuf_bot_iw_I\[10\].z vssd1 vssd1 vccd1 vccd1 um_iw[82] sky130_fd_sc_hd__buf_2
XFILLER_0_12_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[0\].zbuf_bot_iw_I\[12\].genblk1.cell0_I net505 net447 vssd1 vssd1 vccd1 vccd1
+ col\[0\].zbuf_bot_iw_I\[12\].z sky130_fd_sc_hd__and2_1
XFILLER_0_14_1968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_2269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xzbuf_bus_iw_I\[2\].genblk1.cell0_I net10 net513 vssd1 vssd1 vccd1 vccd1 zbuf_bus_iw_I\[2\].genblk1.l
+ sky130_fd_sc_hd__and2_1
X_0470_ _0096_ _0089_ _0097_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__or3b_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1022_ col\[4\].genblk1.mux4_I\[3\].x _0242_ vssd1 vssd1 vccd1 vccd1 bus_ow\[3\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_15_2934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_2923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcol\[7\].zbuf_top_iw_I\[5\].genblk1.cell0_I net486 net437 vssd1 vssd1 vccd1 vccd1
+ col\[7\].zbuf_top_iw_I\[5\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_2770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0806_ col\[5\].zbuf_top_iw_I\[5\].z vssd1 vssd1 vccd1 vccd1 um_iw[203] sky130_fd_sc_hd__buf_2
XFILLER_0_4_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0737_ col\[3\].zbuf_top_iw_I\[8\].z vssd1 vssd1 vccd1 vccd1 um_iw[134] sky130_fd_sc_hd__buf_2
XFILLER_0_12_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0668_ col\[1\].zbuf_top_iw_I\[11\].z vssd1 vssd1 vccd1 vccd1 um_iw[65] sky130_fd_sc_hd__buf_2
X_0599_ _0162_ vssd1 vssd1 vccd1 vccd1 col\[6\].zbuf_bot_ena_I.e sky130_fd_sc_hd__inv_2
XFILLER_0_7_2501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_2444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_2589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xcol\[6\].genblk1.mux4_I\[7\].cell0_I net251 net278 net305 net331 net473 net460 vssd1
+ vssd1 vccd1 vccd1 col\[6\].genblk1.mux4_I\[7\].x sky130_fd_sc_hd__mux4_1
Xinput300 um_ow[339] vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput311 um_ow[349] vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput344 um_ow[379] vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__clkbuf_2
Xinput333 um_ow[369] vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__clkbuf_2
Xinput322 um_ow[359] vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput388 um_ow[72] vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__clkbuf_1
Xinput355 um_ow[42] vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__clkbuf_2
Xinput377 um_ow[62] vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__clkbuf_1
Xinput366 um_ow[52] vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_1
Xinput399 um_ow[82] vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_2910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcol\[2\].zbuf_bot_iw_I\[11\].genblk1.cell0_I net507 net445 vssd1 vssd1 vccd1 vccd1
+ col\[2\].zbuf_bot_iw_I\[11\].z sky130_fd_sc_hd__and2_1
XFILLER_0_6_2099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 col\[0\].zbuf_bot_iw_I\[12\].a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0522_ _0124_ _0121_ _0122_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__or3b_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0453_ _0091_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__clkbuf_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0384_ _0043_ _0045_ _0047_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__or3_1
X_1005_ col\[2\].genblk1.mux4_I\[10\].x _0225_ vssd1 vssd1 vccd1 vccd1 bus_ow\[10\]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_4_2729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xcol\[2\].genblk1.mux4_I\[5\].cell0_I net37 net63 net89 net116 net469 net455 vssd1
+ vssd1 vccd1 vccd1 col\[2\].genblk1.mux4_I\[5\].x sky130_fd_sc_hd__mux4_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_2342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_2353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_2239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_2149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput130 um_ow[186] vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__clkbuf_1
Xinput141 um_ow[196] vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__clkbuf_1
Xinput152 um_ow[205] vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__clkbuf_1
Xinput163 um_ow[215] vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_1
Xinput174 um_ow[225] vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_1
Xinput185 um_ow[235] vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_1
Xinput196 um_ow[245] vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_8_1405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_2915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_2661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0505_ _0111_ _0108_ _0109_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__or3b_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0436_ _0081_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__clkbuf_1
.ends

