// This is the unpowered netlist.
module tt_mux (k_one,
    k_zero,
    addr,
    spine_iw,
    spine_ow,
    um_ena,
    um_iw,
    um_k_zero,
    um_ow);
 output k_one;
 output k_zero;
 input [4:0] addr;
 input [30:0] spine_iw;
 output [25:0] spine_ow;
 output [15:0] um_ena;
 output [287:0] um_iw;
 output [15:0] um_k_zero;
 input [383:0] um_ow;

 wire net552;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire \bus_ow[0] ;
 wire \bus_ow[10] ;
 wire \bus_ow[11] ;
 wire \bus_ow[12] ;
 wire \bus_ow[13] ;
 wire \bus_ow[14] ;
 wire \bus_ow[15] ;
 wire \bus_ow[16] ;
 wire \bus_ow[17] ;
 wire \bus_ow[18] ;
 wire \bus_ow[19] ;
 wire \bus_ow[1] ;
 wire \bus_ow[20] ;
 wire \bus_ow[21] ;
 wire \bus_ow[22] ;
 wire \bus_ow[23] ;
 wire \bus_ow[2] ;
 wire \bus_ow[3] ;
 wire \bus_ow[4] ;
 wire \bus_ow[5] ;
 wire \bus_ow[6] ;
 wire \bus_ow[7] ;
 wire \bus_ow[8] ;
 wire \bus_ow[9] ;
 wire \col[0].genblk1.mux4_I[0].x ;
 wire \col[0].genblk1.mux4_I[10].x ;
 wire \col[0].genblk1.mux4_I[11].x ;
 wire \col[0].genblk1.mux4_I[12].x ;
 wire \col[0].genblk1.mux4_I[13].x ;
 wire \col[0].genblk1.mux4_I[14].x ;
 wire \col[0].genblk1.mux4_I[15].x ;
 wire \col[0].genblk1.mux4_I[16].x ;
 wire \col[0].genblk1.mux4_I[17].x ;
 wire \col[0].genblk1.mux4_I[18].x ;
 wire \col[0].genblk1.mux4_I[19].x ;
 wire \col[0].genblk1.mux4_I[1].x ;
 wire \col[0].genblk1.mux4_I[20].x ;
 wire \col[0].genblk1.mux4_I[21].x ;
 wire \col[0].genblk1.mux4_I[22].x ;
 wire \col[0].genblk1.mux4_I[23].x ;
 wire \col[0].genblk1.mux4_I[2].x ;
 wire \col[0].genblk1.mux4_I[3].x ;
 wire \col[0].genblk1.mux4_I[4].x ;
 wire \col[0].genblk1.mux4_I[5].x ;
 wire \col[0].genblk1.mux4_I[6].x ;
 wire \col[0].genblk1.mux4_I[7].x ;
 wire \col[0].genblk1.mux4_I[8].x ;
 wire \col[0].genblk1.mux4_I[9].x ;
 wire \col[0].zbuf_bot_ena_I.e ;
 wire \col[0].zbuf_bot_ena_I.z ;
 wire \col[0].zbuf_bot_iw_I[0].a ;
 wire \col[0].zbuf_bot_iw_I[0].z ;
 wire \col[0].zbuf_bot_iw_I[10].a ;
 wire \col[0].zbuf_bot_iw_I[10].z ;
 wire \col[0].zbuf_bot_iw_I[11].a ;
 wire \col[0].zbuf_bot_iw_I[11].z ;
 wire \col[0].zbuf_bot_iw_I[12].a ;
 wire \col[0].zbuf_bot_iw_I[12].z ;
 wire \col[0].zbuf_bot_iw_I[13].a ;
 wire \col[0].zbuf_bot_iw_I[13].z ;
 wire \col[0].zbuf_bot_iw_I[14].a ;
 wire \col[0].zbuf_bot_iw_I[14].z ;
 wire \col[0].zbuf_bot_iw_I[15].a ;
 wire \col[0].zbuf_bot_iw_I[15].z ;
 wire \col[0].zbuf_bot_iw_I[16].a ;
 wire \col[0].zbuf_bot_iw_I[16].z ;
 wire \col[0].zbuf_bot_iw_I[17].a ;
 wire \col[0].zbuf_bot_iw_I[17].z ;
 wire \col[0].zbuf_bot_iw_I[1].a ;
 wire \col[0].zbuf_bot_iw_I[1].z ;
 wire \col[0].zbuf_bot_iw_I[2].a ;
 wire \col[0].zbuf_bot_iw_I[2].z ;
 wire \col[0].zbuf_bot_iw_I[3].a ;
 wire \col[0].zbuf_bot_iw_I[3].z ;
 wire \col[0].zbuf_bot_iw_I[4].a ;
 wire \col[0].zbuf_bot_iw_I[4].z ;
 wire \col[0].zbuf_bot_iw_I[5].a ;
 wire \col[0].zbuf_bot_iw_I[5].z ;
 wire \col[0].zbuf_bot_iw_I[6].a ;
 wire \col[0].zbuf_bot_iw_I[6].z ;
 wire \col[0].zbuf_bot_iw_I[7].a ;
 wire \col[0].zbuf_bot_iw_I[7].z ;
 wire \col[0].zbuf_bot_iw_I[8].a ;
 wire \col[0].zbuf_bot_iw_I[8].z ;
 wire \col[0].zbuf_bot_iw_I[9].a ;
 wire \col[0].zbuf_bot_iw_I[9].z ;
 wire \col[0].zbuf_top_ena_I.e ;
 wire \col[0].zbuf_top_ena_I.z ;
 wire \col[0].zbuf_top_iw_I[0].z ;
 wire \col[0].zbuf_top_iw_I[10].z ;
 wire \col[0].zbuf_top_iw_I[11].z ;
 wire \col[0].zbuf_top_iw_I[12].z ;
 wire \col[0].zbuf_top_iw_I[13].z ;
 wire \col[0].zbuf_top_iw_I[14].z ;
 wire \col[0].zbuf_top_iw_I[15].z ;
 wire \col[0].zbuf_top_iw_I[16].z ;
 wire \col[0].zbuf_top_iw_I[17].z ;
 wire \col[0].zbuf_top_iw_I[1].z ;
 wire \col[0].zbuf_top_iw_I[2].z ;
 wire \col[0].zbuf_top_iw_I[3].z ;
 wire \col[0].zbuf_top_iw_I[4].z ;
 wire \col[0].zbuf_top_iw_I[5].z ;
 wire \col[0].zbuf_top_iw_I[6].z ;
 wire \col[0].zbuf_top_iw_I[7].z ;
 wire \col[0].zbuf_top_iw_I[8].z ;
 wire \col[0].zbuf_top_iw_I[9].z ;
 wire \col[1].zbuf_bot_ena_I.e ;
 wire \col[1].zbuf_bot_ena_I.z ;
 wire \col[1].zbuf_bot_iw_I[0].z ;
 wire \col[1].zbuf_bot_iw_I[10].z ;
 wire \col[1].zbuf_bot_iw_I[11].z ;
 wire \col[1].zbuf_bot_iw_I[12].z ;
 wire \col[1].zbuf_bot_iw_I[13].z ;
 wire \col[1].zbuf_bot_iw_I[14].z ;
 wire \col[1].zbuf_bot_iw_I[15].z ;
 wire \col[1].zbuf_bot_iw_I[16].z ;
 wire \col[1].zbuf_bot_iw_I[17].z ;
 wire \col[1].zbuf_bot_iw_I[1].z ;
 wire \col[1].zbuf_bot_iw_I[2].z ;
 wire \col[1].zbuf_bot_iw_I[3].z ;
 wire \col[1].zbuf_bot_iw_I[4].z ;
 wire \col[1].zbuf_bot_iw_I[5].z ;
 wire \col[1].zbuf_bot_iw_I[6].z ;
 wire \col[1].zbuf_bot_iw_I[7].z ;
 wire \col[1].zbuf_bot_iw_I[8].z ;
 wire \col[1].zbuf_bot_iw_I[9].z ;
 wire \col[1].zbuf_top_ena_I.e ;
 wire \col[1].zbuf_top_ena_I.z ;
 wire \col[1].zbuf_top_iw_I[0].z ;
 wire \col[1].zbuf_top_iw_I[10].z ;
 wire \col[1].zbuf_top_iw_I[11].z ;
 wire \col[1].zbuf_top_iw_I[12].z ;
 wire \col[1].zbuf_top_iw_I[13].z ;
 wire \col[1].zbuf_top_iw_I[14].z ;
 wire \col[1].zbuf_top_iw_I[15].z ;
 wire \col[1].zbuf_top_iw_I[16].z ;
 wire \col[1].zbuf_top_iw_I[17].z ;
 wire \col[1].zbuf_top_iw_I[1].z ;
 wire \col[1].zbuf_top_iw_I[2].z ;
 wire \col[1].zbuf_top_iw_I[3].z ;
 wire \col[1].zbuf_top_iw_I[4].z ;
 wire \col[1].zbuf_top_iw_I[5].z ;
 wire \col[1].zbuf_top_iw_I[6].z ;
 wire \col[1].zbuf_top_iw_I[7].z ;
 wire \col[1].zbuf_top_iw_I[8].z ;
 wire \col[1].zbuf_top_iw_I[9].z ;
 wire \col[2].genblk1.mux4_I[0].x ;
 wire \col[2].genblk1.mux4_I[10].x ;
 wire \col[2].genblk1.mux4_I[11].x ;
 wire \col[2].genblk1.mux4_I[12].x ;
 wire \col[2].genblk1.mux4_I[13].x ;
 wire \col[2].genblk1.mux4_I[14].x ;
 wire \col[2].genblk1.mux4_I[15].x ;
 wire \col[2].genblk1.mux4_I[16].x ;
 wire \col[2].genblk1.mux4_I[17].x ;
 wire \col[2].genblk1.mux4_I[18].x ;
 wire \col[2].genblk1.mux4_I[19].x ;
 wire \col[2].genblk1.mux4_I[1].x ;
 wire \col[2].genblk1.mux4_I[20].x ;
 wire \col[2].genblk1.mux4_I[21].x ;
 wire \col[2].genblk1.mux4_I[22].x ;
 wire \col[2].genblk1.mux4_I[23].x ;
 wire \col[2].genblk1.mux4_I[2].x ;
 wire \col[2].genblk1.mux4_I[3].x ;
 wire \col[2].genblk1.mux4_I[4].x ;
 wire \col[2].genblk1.mux4_I[5].x ;
 wire \col[2].genblk1.mux4_I[6].x ;
 wire \col[2].genblk1.mux4_I[7].x ;
 wire \col[2].genblk1.mux4_I[8].x ;
 wire \col[2].genblk1.mux4_I[9].x ;
 wire \col[2].zbuf_bot_ena_I.e ;
 wire \col[2].zbuf_bot_ena_I.z ;
 wire \col[2].zbuf_bot_iw_I[0].z ;
 wire \col[2].zbuf_bot_iw_I[10].z ;
 wire \col[2].zbuf_bot_iw_I[11].z ;
 wire \col[2].zbuf_bot_iw_I[12].z ;
 wire \col[2].zbuf_bot_iw_I[13].z ;
 wire \col[2].zbuf_bot_iw_I[14].z ;
 wire \col[2].zbuf_bot_iw_I[15].z ;
 wire \col[2].zbuf_bot_iw_I[16].z ;
 wire \col[2].zbuf_bot_iw_I[17].z ;
 wire \col[2].zbuf_bot_iw_I[1].z ;
 wire \col[2].zbuf_bot_iw_I[2].z ;
 wire \col[2].zbuf_bot_iw_I[3].z ;
 wire \col[2].zbuf_bot_iw_I[4].z ;
 wire \col[2].zbuf_bot_iw_I[5].z ;
 wire \col[2].zbuf_bot_iw_I[6].z ;
 wire \col[2].zbuf_bot_iw_I[7].z ;
 wire \col[2].zbuf_bot_iw_I[8].z ;
 wire \col[2].zbuf_bot_iw_I[9].z ;
 wire \col[2].zbuf_top_ena_I.e ;
 wire \col[2].zbuf_top_ena_I.z ;
 wire \col[2].zbuf_top_iw_I[0].z ;
 wire \col[2].zbuf_top_iw_I[10].z ;
 wire \col[2].zbuf_top_iw_I[11].z ;
 wire \col[2].zbuf_top_iw_I[12].z ;
 wire \col[2].zbuf_top_iw_I[13].z ;
 wire \col[2].zbuf_top_iw_I[14].z ;
 wire \col[2].zbuf_top_iw_I[15].z ;
 wire \col[2].zbuf_top_iw_I[16].z ;
 wire \col[2].zbuf_top_iw_I[17].z ;
 wire \col[2].zbuf_top_iw_I[1].z ;
 wire \col[2].zbuf_top_iw_I[2].z ;
 wire \col[2].zbuf_top_iw_I[3].z ;
 wire \col[2].zbuf_top_iw_I[4].z ;
 wire \col[2].zbuf_top_iw_I[5].z ;
 wire \col[2].zbuf_top_iw_I[6].z ;
 wire \col[2].zbuf_top_iw_I[7].z ;
 wire \col[2].zbuf_top_iw_I[8].z ;
 wire \col[2].zbuf_top_iw_I[9].z ;
 wire \col[3].zbuf_bot_ena_I.e ;
 wire \col[3].zbuf_bot_ena_I.z ;
 wire \col[3].zbuf_bot_iw_I[0].z ;
 wire \col[3].zbuf_bot_iw_I[10].z ;
 wire \col[3].zbuf_bot_iw_I[11].z ;
 wire \col[3].zbuf_bot_iw_I[12].z ;
 wire \col[3].zbuf_bot_iw_I[13].z ;
 wire \col[3].zbuf_bot_iw_I[14].z ;
 wire \col[3].zbuf_bot_iw_I[15].z ;
 wire \col[3].zbuf_bot_iw_I[16].z ;
 wire \col[3].zbuf_bot_iw_I[17].z ;
 wire \col[3].zbuf_bot_iw_I[1].z ;
 wire \col[3].zbuf_bot_iw_I[2].z ;
 wire \col[3].zbuf_bot_iw_I[3].z ;
 wire \col[3].zbuf_bot_iw_I[4].z ;
 wire \col[3].zbuf_bot_iw_I[5].z ;
 wire \col[3].zbuf_bot_iw_I[6].z ;
 wire \col[3].zbuf_bot_iw_I[7].z ;
 wire \col[3].zbuf_bot_iw_I[8].z ;
 wire \col[3].zbuf_bot_iw_I[9].z ;
 wire \col[3].zbuf_top_ena_I.e ;
 wire \col[3].zbuf_top_ena_I.z ;
 wire \col[3].zbuf_top_iw_I[0].z ;
 wire \col[3].zbuf_top_iw_I[10].z ;
 wire \col[3].zbuf_top_iw_I[11].z ;
 wire \col[3].zbuf_top_iw_I[12].z ;
 wire \col[3].zbuf_top_iw_I[13].z ;
 wire \col[3].zbuf_top_iw_I[14].z ;
 wire \col[3].zbuf_top_iw_I[15].z ;
 wire \col[3].zbuf_top_iw_I[16].z ;
 wire \col[3].zbuf_top_iw_I[17].z ;
 wire \col[3].zbuf_top_iw_I[1].z ;
 wire \col[3].zbuf_top_iw_I[2].z ;
 wire \col[3].zbuf_top_iw_I[3].z ;
 wire \col[3].zbuf_top_iw_I[4].z ;
 wire \col[3].zbuf_top_iw_I[5].z ;
 wire \col[3].zbuf_top_iw_I[6].z ;
 wire \col[3].zbuf_top_iw_I[7].z ;
 wire \col[3].zbuf_top_iw_I[8].z ;
 wire \col[3].zbuf_top_iw_I[9].z ;
 wire \col[4].genblk1.mux4_I[0].x ;
 wire \col[4].genblk1.mux4_I[10].x ;
 wire \col[4].genblk1.mux4_I[11].x ;
 wire \col[4].genblk1.mux4_I[12].x ;
 wire \col[4].genblk1.mux4_I[13].x ;
 wire \col[4].genblk1.mux4_I[14].x ;
 wire \col[4].genblk1.mux4_I[15].x ;
 wire \col[4].genblk1.mux4_I[16].x ;
 wire \col[4].genblk1.mux4_I[17].x ;
 wire \col[4].genblk1.mux4_I[18].x ;
 wire \col[4].genblk1.mux4_I[19].x ;
 wire \col[4].genblk1.mux4_I[1].x ;
 wire \col[4].genblk1.mux4_I[20].x ;
 wire \col[4].genblk1.mux4_I[21].x ;
 wire \col[4].genblk1.mux4_I[22].x ;
 wire \col[4].genblk1.mux4_I[23].x ;
 wire \col[4].genblk1.mux4_I[2].x ;
 wire \col[4].genblk1.mux4_I[3].x ;
 wire \col[4].genblk1.mux4_I[4].x ;
 wire \col[4].genblk1.mux4_I[5].x ;
 wire \col[4].genblk1.mux4_I[6].x ;
 wire \col[4].genblk1.mux4_I[7].x ;
 wire \col[4].genblk1.mux4_I[8].x ;
 wire \col[4].genblk1.mux4_I[9].x ;
 wire \col[4].zbuf_bot_ena_I.e ;
 wire \col[4].zbuf_bot_ena_I.z ;
 wire \col[4].zbuf_bot_iw_I[0].z ;
 wire \col[4].zbuf_bot_iw_I[10].z ;
 wire \col[4].zbuf_bot_iw_I[11].z ;
 wire \col[4].zbuf_bot_iw_I[12].z ;
 wire \col[4].zbuf_bot_iw_I[13].z ;
 wire \col[4].zbuf_bot_iw_I[14].z ;
 wire \col[4].zbuf_bot_iw_I[15].z ;
 wire \col[4].zbuf_bot_iw_I[16].z ;
 wire \col[4].zbuf_bot_iw_I[17].z ;
 wire \col[4].zbuf_bot_iw_I[1].z ;
 wire \col[4].zbuf_bot_iw_I[2].z ;
 wire \col[4].zbuf_bot_iw_I[3].z ;
 wire \col[4].zbuf_bot_iw_I[4].z ;
 wire \col[4].zbuf_bot_iw_I[5].z ;
 wire \col[4].zbuf_bot_iw_I[6].z ;
 wire \col[4].zbuf_bot_iw_I[7].z ;
 wire \col[4].zbuf_bot_iw_I[8].z ;
 wire \col[4].zbuf_bot_iw_I[9].z ;
 wire \col[4].zbuf_top_ena_I.e ;
 wire \col[4].zbuf_top_ena_I.z ;
 wire \col[4].zbuf_top_iw_I[0].z ;
 wire \col[4].zbuf_top_iw_I[10].z ;
 wire \col[4].zbuf_top_iw_I[11].z ;
 wire \col[4].zbuf_top_iw_I[12].z ;
 wire \col[4].zbuf_top_iw_I[13].z ;
 wire \col[4].zbuf_top_iw_I[14].z ;
 wire \col[4].zbuf_top_iw_I[15].z ;
 wire \col[4].zbuf_top_iw_I[16].z ;
 wire \col[4].zbuf_top_iw_I[17].z ;
 wire \col[4].zbuf_top_iw_I[1].z ;
 wire \col[4].zbuf_top_iw_I[2].z ;
 wire \col[4].zbuf_top_iw_I[3].z ;
 wire \col[4].zbuf_top_iw_I[4].z ;
 wire \col[4].zbuf_top_iw_I[5].z ;
 wire \col[4].zbuf_top_iw_I[6].z ;
 wire \col[4].zbuf_top_iw_I[7].z ;
 wire \col[4].zbuf_top_iw_I[8].z ;
 wire \col[4].zbuf_top_iw_I[9].z ;
 wire \col[5].zbuf_bot_ena_I.e ;
 wire \col[5].zbuf_bot_ena_I.z ;
 wire \col[5].zbuf_bot_iw_I[0].z ;
 wire \col[5].zbuf_bot_iw_I[10].z ;
 wire \col[5].zbuf_bot_iw_I[11].z ;
 wire \col[5].zbuf_bot_iw_I[12].z ;
 wire \col[5].zbuf_bot_iw_I[13].z ;
 wire \col[5].zbuf_bot_iw_I[14].z ;
 wire \col[5].zbuf_bot_iw_I[15].z ;
 wire \col[5].zbuf_bot_iw_I[16].z ;
 wire \col[5].zbuf_bot_iw_I[17].z ;
 wire \col[5].zbuf_bot_iw_I[1].z ;
 wire \col[5].zbuf_bot_iw_I[2].z ;
 wire \col[5].zbuf_bot_iw_I[3].z ;
 wire \col[5].zbuf_bot_iw_I[4].z ;
 wire \col[5].zbuf_bot_iw_I[5].z ;
 wire \col[5].zbuf_bot_iw_I[6].z ;
 wire \col[5].zbuf_bot_iw_I[7].z ;
 wire \col[5].zbuf_bot_iw_I[8].z ;
 wire \col[5].zbuf_bot_iw_I[9].z ;
 wire \col[5].zbuf_top_ena_I.e ;
 wire \col[5].zbuf_top_ena_I.z ;
 wire \col[5].zbuf_top_iw_I[0].z ;
 wire \col[5].zbuf_top_iw_I[10].z ;
 wire \col[5].zbuf_top_iw_I[11].z ;
 wire \col[5].zbuf_top_iw_I[12].z ;
 wire \col[5].zbuf_top_iw_I[13].z ;
 wire \col[5].zbuf_top_iw_I[14].z ;
 wire \col[5].zbuf_top_iw_I[15].z ;
 wire \col[5].zbuf_top_iw_I[16].z ;
 wire \col[5].zbuf_top_iw_I[17].z ;
 wire \col[5].zbuf_top_iw_I[1].z ;
 wire \col[5].zbuf_top_iw_I[2].z ;
 wire \col[5].zbuf_top_iw_I[3].z ;
 wire \col[5].zbuf_top_iw_I[4].z ;
 wire \col[5].zbuf_top_iw_I[5].z ;
 wire \col[5].zbuf_top_iw_I[6].z ;
 wire \col[5].zbuf_top_iw_I[7].z ;
 wire \col[5].zbuf_top_iw_I[8].z ;
 wire \col[5].zbuf_top_iw_I[9].z ;
 wire \col[6].genblk1.mux4_I[0].x ;
 wire \col[6].genblk1.mux4_I[10].x ;
 wire \col[6].genblk1.mux4_I[11].x ;
 wire \col[6].genblk1.mux4_I[12].x ;
 wire \col[6].genblk1.mux4_I[13].x ;
 wire \col[6].genblk1.mux4_I[14].x ;
 wire \col[6].genblk1.mux4_I[15].x ;
 wire \col[6].genblk1.mux4_I[16].x ;
 wire \col[6].genblk1.mux4_I[17].x ;
 wire \col[6].genblk1.mux4_I[18].x ;
 wire \col[6].genblk1.mux4_I[19].x ;
 wire \col[6].genblk1.mux4_I[1].x ;
 wire \col[6].genblk1.mux4_I[20].x ;
 wire \col[6].genblk1.mux4_I[21].x ;
 wire \col[6].genblk1.mux4_I[22].x ;
 wire \col[6].genblk1.mux4_I[23].x ;
 wire \col[6].genblk1.mux4_I[2].x ;
 wire \col[6].genblk1.mux4_I[3].x ;
 wire \col[6].genblk1.mux4_I[4].x ;
 wire \col[6].genblk1.mux4_I[5].x ;
 wire \col[6].genblk1.mux4_I[6].x ;
 wire \col[6].genblk1.mux4_I[7].x ;
 wire \col[6].genblk1.mux4_I[8].x ;
 wire \col[6].genblk1.mux4_I[9].x ;
 wire \col[6].zbuf_bot_ena_I.e ;
 wire \col[6].zbuf_bot_ena_I.z ;
 wire \col[6].zbuf_bot_iw_I[0].z ;
 wire \col[6].zbuf_bot_iw_I[10].z ;
 wire \col[6].zbuf_bot_iw_I[11].z ;
 wire \col[6].zbuf_bot_iw_I[12].z ;
 wire \col[6].zbuf_bot_iw_I[13].z ;
 wire \col[6].zbuf_bot_iw_I[14].z ;
 wire \col[6].zbuf_bot_iw_I[15].z ;
 wire \col[6].zbuf_bot_iw_I[16].z ;
 wire \col[6].zbuf_bot_iw_I[17].z ;
 wire \col[6].zbuf_bot_iw_I[1].z ;
 wire \col[6].zbuf_bot_iw_I[2].z ;
 wire \col[6].zbuf_bot_iw_I[3].z ;
 wire \col[6].zbuf_bot_iw_I[4].z ;
 wire \col[6].zbuf_bot_iw_I[5].z ;
 wire \col[6].zbuf_bot_iw_I[6].z ;
 wire \col[6].zbuf_bot_iw_I[7].z ;
 wire \col[6].zbuf_bot_iw_I[8].z ;
 wire \col[6].zbuf_bot_iw_I[9].z ;
 wire \col[6].zbuf_top_ena_I.e ;
 wire \col[6].zbuf_top_ena_I.z ;
 wire \col[6].zbuf_top_iw_I[0].z ;
 wire \col[6].zbuf_top_iw_I[10].z ;
 wire \col[6].zbuf_top_iw_I[11].z ;
 wire \col[6].zbuf_top_iw_I[12].z ;
 wire \col[6].zbuf_top_iw_I[13].z ;
 wire \col[6].zbuf_top_iw_I[14].z ;
 wire \col[6].zbuf_top_iw_I[15].z ;
 wire \col[6].zbuf_top_iw_I[16].z ;
 wire \col[6].zbuf_top_iw_I[17].z ;
 wire \col[6].zbuf_top_iw_I[1].z ;
 wire \col[6].zbuf_top_iw_I[2].z ;
 wire \col[6].zbuf_top_iw_I[3].z ;
 wire \col[6].zbuf_top_iw_I[4].z ;
 wire \col[6].zbuf_top_iw_I[5].z ;
 wire \col[6].zbuf_top_iw_I[6].z ;
 wire \col[6].zbuf_top_iw_I[7].z ;
 wire \col[6].zbuf_top_iw_I[8].z ;
 wire \col[6].zbuf_top_iw_I[9].z ;
 wire \col[7].zbuf_bot_ena_I.e ;
 wire \col[7].zbuf_bot_ena_I.z ;
 wire \col[7].zbuf_bot_iw_I[0].z ;
 wire \col[7].zbuf_bot_iw_I[10].z ;
 wire \col[7].zbuf_bot_iw_I[11].z ;
 wire \col[7].zbuf_bot_iw_I[12].z ;
 wire \col[7].zbuf_bot_iw_I[13].z ;
 wire \col[7].zbuf_bot_iw_I[14].z ;
 wire \col[7].zbuf_bot_iw_I[15].z ;
 wire \col[7].zbuf_bot_iw_I[16].z ;
 wire \col[7].zbuf_bot_iw_I[17].z ;
 wire \col[7].zbuf_bot_iw_I[1].z ;
 wire \col[7].zbuf_bot_iw_I[2].z ;
 wire \col[7].zbuf_bot_iw_I[3].z ;
 wire \col[7].zbuf_bot_iw_I[4].z ;
 wire \col[7].zbuf_bot_iw_I[5].z ;
 wire \col[7].zbuf_bot_iw_I[6].z ;
 wire \col[7].zbuf_bot_iw_I[7].z ;
 wire \col[7].zbuf_bot_iw_I[8].z ;
 wire \col[7].zbuf_bot_iw_I[9].z ;
 wire \col[7].zbuf_top_ena_I.e ;
 wire \col[7].zbuf_top_ena_I.z ;
 wire \col[7].zbuf_top_iw_I[0].z ;
 wire \col[7].zbuf_top_iw_I[10].z ;
 wire \col[7].zbuf_top_iw_I[11].z ;
 wire \col[7].zbuf_top_iw_I[12].z ;
 wire \col[7].zbuf_top_iw_I[13].z ;
 wire \col[7].zbuf_top_iw_I[14].z ;
 wire \col[7].zbuf_top_iw_I[15].z ;
 wire \col[7].zbuf_top_iw_I[16].z ;
 wire \col[7].zbuf_top_iw_I[17].z ;
 wire \col[7].zbuf_top_iw_I[1].z ;
 wire \col[7].zbuf_top_iw_I[2].z ;
 wire \col[7].zbuf_top_iw_I[3].z ;
 wire \col[7].zbuf_top_iw_I[4].z ;
 wire \col[7].zbuf_top_iw_I[5].z ;
 wire \col[7].zbuf_top_iw_I[6].z ;
 wire \col[7].zbuf_top_iw_I[7].z ;
 wire \col[7].zbuf_top_iw_I[8].z ;
 wire \col[7].zbuf_top_iw_I[9].z ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net52;
 wire net53;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \zbuf_bus_ena_I.e ;
 wire \zbuf_bus_ena_I.genblk1.l ;
 wire \zbuf_bus_ena_I.z ;
 wire \zbuf_bus_iw_I[0].genblk1.l ;
 wire \zbuf_bus_iw_I[10].genblk1.l ;
 wire \zbuf_bus_iw_I[11].genblk1.l ;
 wire \zbuf_bus_iw_I[12].genblk1.l ;
 wire \zbuf_bus_iw_I[13].genblk1.l ;
 wire \zbuf_bus_iw_I[14].genblk1.l ;
 wire \zbuf_bus_iw_I[15].genblk1.l ;
 wire \zbuf_bus_iw_I[16].genblk1.l ;
 wire \zbuf_bus_iw_I[17].genblk1.l ;
 wire \zbuf_bus_iw_I[1].genblk1.l ;
 wire \zbuf_bus_iw_I[2].genblk1.l ;
 wire \zbuf_bus_iw_I[3].genblk1.l ;
 wire \zbuf_bus_iw_I[4].genblk1.l ;
 wire \zbuf_bus_iw_I[5].genblk1.l ;
 wire \zbuf_bus_iw_I[6].genblk1.l ;
 wire \zbuf_bus_iw_I[7].genblk1.l ;
 wire \zbuf_bus_iw_I[8].genblk1.l ;
 wire \zbuf_bus_iw_I[9].genblk1.l ;
 wire \zbuf_bus_sel_I[0].genblk1.l ;
 wire \zbuf_bus_sel_I[0].z ;
 wire \zbuf_bus_sel_I[1].genblk1.l ;
 wire \zbuf_bus_sel_I[1].z ;
 wire \zbuf_bus_sel_I[2].genblk1.l ;
 wire \zbuf_bus_sel_I[2].z ;
 wire \zbuf_bus_sel_I[3].genblk1.l ;
 wire \zbuf_bus_sel_I[3].z ;
 wire \zbuf_bus_sel_I[4].genblk1.l ;
 wire \zbuf_bus_sel_I[4].z ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0150_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\col[0].zbuf_bot_iw_I[1].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\col[0].zbuf_bot_iw_I[1].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(\col[0].zbuf_bot_iw_I[13].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\col[0].zbuf_bot_iw_I[3].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\col[0].zbuf_bot_iw_I[4].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\col[0].zbuf_bot_iw_I[4].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\col[0].zbuf_bot_iw_I[5].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\col[0].zbuf_bot_iw_I[5].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(\col[0].zbuf_bot_iw_I[6].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\col[0].zbuf_bot_iw_I[6].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\col[0].zbuf_bot_iw_I[7].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\bus_ow[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\col[0].zbuf_bot_iw_I[8].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\col[0].zbuf_bot_iw_I[8].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(\col[0].zbuf_bot_iw_I[9].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(\col[0].zbuf_bot_iw_I[9].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(spine_iw[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(spine_iw[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(spine_iw[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(spine_iw[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(\zbuf_bus_ena_I.z ));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(\zbuf_bus_ena_I.z ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\col[0].zbuf_bot_iw_I[12].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(\zbuf_bus_ena_I.z ));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\col[0].zbuf_bot_iw_I[12].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\col[0].zbuf_bot_iw_I[13].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\col[0].zbuf_bot_iw_I[16].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\col[0].zbuf_bot_iw_I[16].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\col[0].zbuf_bot_iw_I[17].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(_0145_));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(_0145_));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(_0145_));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(_0145_));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(_0147_));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(_0147_));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(_0147_));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(_0147_));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(\bus_ow[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(\bus_ow[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\col[0].zbuf_bot_iw_I[17].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(spine_iw[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(net477));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1672 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1807 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1827 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1859 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_2029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2039 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2068 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_2073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_2206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_2234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_2465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_2521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2527 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_2597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2736 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_2785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_2822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2844 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2863 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2871 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2891 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2928 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2070 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_2346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_2419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_2685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_2692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_2711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2802 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2826 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_2829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2850 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_2857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_2909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_2350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_2390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_2406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_2417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_2423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_2439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_2701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_2710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_2720 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_2730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_2740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_2813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_2819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_2824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_2828 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_2833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_2840 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_2847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_2854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_2857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2863 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_2875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_2896 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_2913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_2927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_2934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1723 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1731 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1779 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_2209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_2537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_2602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_2805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_2810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_2814 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_2826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_2829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2835 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2870 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2879 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2883 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2915 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_2934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1723 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1815 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1831 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2015 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2042 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_2054 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_2069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2083 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2099 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_2107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_2129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_2185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_2465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_2518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_2797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_2801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_2815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_2821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_2825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_2857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_2865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_2869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_2873 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_2910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_2913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2932 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1690 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1802 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1883 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1896 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2001 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_2041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2057 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2066 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2084 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_2489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2532 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2644 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_2933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1672 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1702 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1790 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1802 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1827 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1859 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1919 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1945 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1971 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_2013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2039 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2057 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_2181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_2461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_2535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2639 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_2769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2934 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1700 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1818 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1826 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1878 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1973 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_2013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2057 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2082 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2098 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_2125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_2293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_2517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2842 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2873 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2882 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2891 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2900 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_2909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2928 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_1649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1730 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_1779 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_1817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1907 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1930 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1986 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2018 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2042 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_2097 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_2381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_2713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2844 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2891 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2900 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_2933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_952 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1828 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_2061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_2193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_2241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_2253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_2257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_2293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_2297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2631 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2639 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2646 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_2685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_2745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_2801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_2809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2822 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2850 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_2877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2882 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2889 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2896 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_2910 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_2934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1676 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_2269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_2321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_2381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_2437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_2460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_2658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_2661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_2670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_2683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_2687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_2717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_2747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_2770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_2773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2814 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2822 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_2877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_2882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2903 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2910 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_2934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1704 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1818 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1830 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_2053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_2221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_2641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2756 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2855 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_2865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2871 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2878 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2919 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1676 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1744 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1827 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2675 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_2825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2846 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2868 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2915 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2924 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2932 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_2229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_2238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_2294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_2306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_2349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_2377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_2409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_2686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_2742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_2809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2820 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2842 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2899 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_2913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2920 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2935 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1579 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1650 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_2037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_2042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_2045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_2055 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2059 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_2338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_2342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_2381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_2434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_2714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_2770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_2773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_2804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_2826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_2829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2840 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2863 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2883 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2903 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2922 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1816 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_2037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_2042 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_2051 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_2249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_2335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_2345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_2349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_2353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_2430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_2434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_2681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_2686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_2733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_2753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2759 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2779 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_2798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2818 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_2854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_2857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2868 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_2913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_2933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_977 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__inv_2 _0303_ (.A(net33),
    .Y(_0000_));
 sky130_fd_sc_hd__nor2_2 _0304_ (.A(net2),
    .B(_0000_),
    .Y(_0001_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0305_ (.A(_0001_),
    .X(_0002_));
 sky130_fd_sc_hd__inv_2 _0306_ (.A(net3),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _0307_ (.A(net31),
    .Y(_0004_));
 sky130_fd_sc_hd__a22o_2 _0308_ (.A1(_0003_),
    .A2(net34),
    .B1(net1),
    .B2(_0004_),
    .X(_0005_));
 sky130_fd_sc_hd__clkbuf_2 _0309_ (.A(_0005_),
    .X(_0006_));
 sky130_fd_sc_hd__or2b_1 _0310_ (.A(net7),
    .B_N(net5),
    .X(_0007_));
 sky130_fd_sc_hd__o221ai_4 _0311_ (.A1(_0003_),
    .A2(net34),
    .B1(net1),
    .B2(_0004_),
    .C1(_0007_),
    .Y(_0008_));
 sky130_fd_sc_hd__clkbuf_2 _0312_ (.A(_0008_),
    .X(_0009_));
 sky130_fd_sc_hd__inv_2 _0313_ (.A(net5),
    .Y(_0010_));
 sky130_fd_sc_hd__xor2_1 _0314_ (.A(net4),
    .B(net6),
    .X(_0011_));
 sky130_fd_sc_hd__a221o_2 _0315_ (.A1(net2),
    .A2(_0000_),
    .B1(_0010_),
    .B2(net7),
    .C1(_0011_),
    .X(_0012_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0316_ (.A(_0012_),
    .X(_0013_));
 sky130_fd_sc_hd__nor4_1 _0317_ (.A(_0002_),
    .B(_0006_),
    .C(_0009_),
    .D(_0013_),
    .Y(\zbuf_bus_ena_I.e ));
 sky130_fd_sc_hd__or4_1 _0318_ (.A(_0002_),
    .B(_0006_),
    .C(_0009_),
    .D(_0013_),
    .X(_0014_));
 sky130_fd_sc_hd__clkbuf_1 _0319_ (.A(_0014_),
    .X(_0168_));
 sky130_fd_sc_hd__or4_1 _0320_ (.A(_0002_),
    .B(_0006_),
    .C(_0009_),
    .D(_0013_),
    .X(_0015_));
 sky130_fd_sc_hd__clkbuf_1 _0321_ (.A(_0015_),
    .X(_0169_));
 sky130_fd_sc_hd__or4_1 _0322_ (.A(_0002_),
    .B(_0006_),
    .C(_0009_),
    .D(_0013_),
    .X(_0016_));
 sky130_fd_sc_hd__clkbuf_1 _0323_ (.A(_0016_),
    .X(_0170_));
 sky130_fd_sc_hd__or4_1 _0324_ (.A(_0002_),
    .B(_0006_),
    .C(_0009_),
    .D(_0013_),
    .X(_0017_));
 sky130_fd_sc_hd__clkbuf_1 _0325_ (.A(_0017_),
    .X(_0171_));
 sky130_fd_sc_hd__or4_1 _0326_ (.A(_0002_),
    .B(_0006_),
    .C(_0009_),
    .D(_0013_),
    .X(_0018_));
 sky130_fd_sc_hd__clkbuf_1 _0327_ (.A(_0018_),
    .X(_0172_));
 sky130_fd_sc_hd__or4_1 _0328_ (.A(_0002_),
    .B(_0006_),
    .C(_0009_),
    .D(_0013_),
    .X(_0019_));
 sky130_fd_sc_hd__clkbuf_1 _0329_ (.A(_0019_),
    .X(_0173_));
 sky130_fd_sc_hd__or4_1 _0330_ (.A(_0002_),
    .B(_0006_),
    .C(_0009_),
    .D(_0013_),
    .X(_0020_));
 sky130_fd_sc_hd__clkbuf_1 _0331_ (.A(_0020_),
    .X(_0174_));
 sky130_fd_sc_hd__or4_1 _0332_ (.A(_0002_),
    .B(_0006_),
    .C(_0009_),
    .D(_0013_),
    .X(_0021_));
 sky130_fd_sc_hd__clkbuf_1 _0333_ (.A(_0021_),
    .X(_0175_));
 sky130_fd_sc_hd__or4_1 _0334_ (.A(_0002_),
    .B(_0006_),
    .C(_0009_),
    .D(_0013_),
    .X(_0022_));
 sky130_fd_sc_hd__clkbuf_1 _0335_ (.A(_0022_),
    .X(_0176_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0336_ (.A(_0001_),
    .X(_0023_));
 sky130_fd_sc_hd__clkbuf_2 _0337_ (.A(_0005_),
    .X(_0024_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0338_ (.A(_0008_),
    .X(_0025_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0339_ (.A(_0012_),
    .X(_0026_));
 sky130_fd_sc_hd__or4_1 _0340_ (.A(_0023_),
    .B(_0024_),
    .C(_0025_),
    .D(_0026_),
    .X(_0027_));
 sky130_fd_sc_hd__clkbuf_1 _0341_ (.A(_0027_),
    .X(_0177_));
 sky130_fd_sc_hd__or4_1 _0342_ (.A(_0023_),
    .B(_0024_),
    .C(_0025_),
    .D(_0026_),
    .X(_0028_));
 sky130_fd_sc_hd__clkbuf_1 _0343_ (.A(_0028_),
    .X(_0178_));
 sky130_fd_sc_hd__or4_1 _0344_ (.A(_0023_),
    .B(_0024_),
    .C(_0025_),
    .D(_0026_),
    .X(_0029_));
 sky130_fd_sc_hd__clkbuf_1 _0345_ (.A(_0029_),
    .X(_0179_));
 sky130_fd_sc_hd__or4_1 _0346_ (.A(_0023_),
    .B(_0024_),
    .C(_0025_),
    .D(_0026_),
    .X(_0030_));
 sky130_fd_sc_hd__clkbuf_1 _0347_ (.A(_0030_),
    .X(_0180_));
 sky130_fd_sc_hd__or4_1 _0348_ (.A(_0023_),
    .B(_0024_),
    .C(_0025_),
    .D(_0026_),
    .X(_0031_));
 sky130_fd_sc_hd__clkbuf_1 _0349_ (.A(_0031_),
    .X(_0181_));
 sky130_fd_sc_hd__or4_1 _0350_ (.A(_0023_),
    .B(_0024_),
    .C(_0025_),
    .D(_0026_),
    .X(_0032_));
 sky130_fd_sc_hd__clkbuf_1 _0351_ (.A(_0032_),
    .X(_0182_));
 sky130_fd_sc_hd__or4_1 _0352_ (.A(_0023_),
    .B(_0024_),
    .C(_0025_),
    .D(_0026_),
    .X(_0033_));
 sky130_fd_sc_hd__clkbuf_1 _0353_ (.A(_0033_),
    .X(_0183_));
 sky130_fd_sc_hd__or4_1 _0354_ (.A(_0023_),
    .B(_0024_),
    .C(_0025_),
    .D(_0026_),
    .X(_0034_));
 sky130_fd_sc_hd__clkbuf_1 _0355_ (.A(_0034_),
    .X(_0184_));
 sky130_fd_sc_hd__or4_1 _0356_ (.A(_0023_),
    .B(_0024_),
    .C(_0025_),
    .D(_0026_),
    .X(_0035_));
 sky130_fd_sc_hd__clkbuf_1 _0357_ (.A(_0035_),
    .X(_0185_));
 sky130_fd_sc_hd__or4_1 _0358_ (.A(_0023_),
    .B(_0024_),
    .C(_0025_),
    .D(_0026_),
    .X(_0036_));
 sky130_fd_sc_hd__clkbuf_1 _0359_ (.A(_0036_),
    .X(_0186_));
 sky130_fd_sc_hd__or4_1 _0360_ (.A(_0001_),
    .B(_0005_),
    .C(_0008_),
    .D(_0012_),
    .X(_0037_));
 sky130_fd_sc_hd__clkbuf_1 _0361_ (.A(_0037_),
    .X(_0187_));
 sky130_fd_sc_hd__or4_1 _0362_ (.A(_0001_),
    .B(_0005_),
    .C(_0008_),
    .D(_0012_),
    .X(_0038_));
 sky130_fd_sc_hd__clkbuf_1 _0363_ (.A(_0038_),
    .X(_0188_));
 sky130_fd_sc_hd__or4_1 _0364_ (.A(_0001_),
    .B(_0005_),
    .C(_0008_),
    .D(_0012_),
    .X(_0039_));
 sky130_fd_sc_hd__clkbuf_1 _0365_ (.A(_0039_),
    .X(_0189_));
 sky130_fd_sc_hd__or4_1 _0366_ (.A(_0001_),
    .B(_0005_),
    .C(_0008_),
    .D(_0012_),
    .X(_0040_));
 sky130_fd_sc_hd__clkbuf_1 _0367_ (.A(_0040_),
    .X(_0190_));
 sky130_fd_sc_hd__or3_1 _0368_ (.A(\zbuf_bus_sel_I[4].z ),
    .B(\zbuf_bus_sel_I[2].z ),
    .C(\zbuf_bus_sel_I[3].z ),
    .X(_0041_));
 sky130_fd_sc_hd__clkbuf_2 _0369_ (.A(_0041_),
    .X(_0192_));
 sky130_fd_sc_hd__clkbuf_4 _0370_ (.A(\zbuf_bus_sel_I[4].z ),
    .X(_0042_));
 sky130_fd_sc_hd__clkbuf_2 _0371_ (.A(_0042_),
    .X(_0043_));
 sky130_fd_sc_hd__clkbuf_4 _0372_ (.A(\zbuf_bus_sel_I[2].z ),
    .X(_0044_));
 sky130_fd_sc_hd__buf_2 _0373_ (.A(_0044_),
    .X(_0045_));
 sky130_fd_sc_hd__clkbuf_4 _0374_ (.A(\zbuf_bus_sel_I[3].z ),
    .X(_0046_));
 sky130_fd_sc_hd__clkbuf_8 _0375_ (.A(_0046_),
    .X(_0047_));
 sky130_fd_sc_hd__or3_1 _0376_ (.A(_0043_),
    .B(_0045_),
    .C(_0047_),
    .X(_0048_));
 sky130_fd_sc_hd__clkbuf_1 _0377_ (.A(_0048_),
    .X(_0193_));
 sky130_fd_sc_hd__or3_1 _0378_ (.A(_0043_),
    .B(_0045_),
    .C(_0047_),
    .X(_0049_));
 sky130_fd_sc_hd__clkbuf_1 _0379_ (.A(_0049_),
    .X(_0194_));
 sky130_fd_sc_hd__or3_1 _0380_ (.A(_0043_),
    .B(_0045_),
    .C(_0047_),
    .X(_0050_));
 sky130_fd_sc_hd__clkbuf_1 _0381_ (.A(_0050_),
    .X(_0195_));
 sky130_fd_sc_hd__or3_1 _0382_ (.A(_0043_),
    .B(_0045_),
    .C(_0047_),
    .X(_0051_));
 sky130_fd_sc_hd__clkbuf_1 _0383_ (.A(_0051_),
    .X(_0196_));
 sky130_fd_sc_hd__or3_1 _0384_ (.A(_0043_),
    .B(_0045_),
    .C(_0047_),
    .X(_0052_));
 sky130_fd_sc_hd__clkbuf_1 _0385_ (.A(_0052_),
    .X(_0197_));
 sky130_fd_sc_hd__clkbuf_2 _0386_ (.A(_0046_),
    .X(_0053_));
 sky130_fd_sc_hd__or3_1 _0387_ (.A(_0043_),
    .B(_0045_),
    .C(_0053_),
    .X(_0054_));
 sky130_fd_sc_hd__clkbuf_1 _0388_ (.A(_0054_),
    .X(_0198_));
 sky130_fd_sc_hd__or3_1 _0389_ (.A(_0043_),
    .B(_0045_),
    .C(_0053_),
    .X(_0055_));
 sky130_fd_sc_hd__clkbuf_1 _0390_ (.A(_0055_),
    .X(_0199_));
 sky130_fd_sc_hd__or3_1 _0391_ (.A(_0043_),
    .B(_0045_),
    .C(_0053_),
    .X(_0056_));
 sky130_fd_sc_hd__clkbuf_1 _0392_ (.A(_0056_),
    .X(_0200_));
 sky130_fd_sc_hd__or3_1 _0393_ (.A(_0043_),
    .B(_0045_),
    .C(_0053_),
    .X(_0057_));
 sky130_fd_sc_hd__clkbuf_1 _0394_ (.A(_0057_),
    .X(_0201_));
 sky130_fd_sc_hd__clkbuf_2 _0395_ (.A(\zbuf_bus_sel_I[4].z ),
    .X(_0058_));
 sky130_fd_sc_hd__clkbuf_2 _0396_ (.A(_0044_),
    .X(_0059_));
 sky130_fd_sc_hd__or3_1 _0397_ (.A(_0058_),
    .B(_0059_),
    .C(_0053_),
    .X(_0060_));
 sky130_fd_sc_hd__clkbuf_1 _0398_ (.A(_0060_),
    .X(_0202_));
 sky130_fd_sc_hd__or3_1 _0399_ (.A(_0058_),
    .B(_0059_),
    .C(_0053_),
    .X(_0061_));
 sky130_fd_sc_hd__clkbuf_1 _0400_ (.A(_0061_),
    .X(_0203_));
 sky130_fd_sc_hd__or3_1 _0401_ (.A(_0058_),
    .B(_0059_),
    .C(_0053_),
    .X(_0062_));
 sky130_fd_sc_hd__clkbuf_1 _0402_ (.A(_0062_),
    .X(_0204_));
 sky130_fd_sc_hd__or3_1 _0403_ (.A(_0058_),
    .B(_0059_),
    .C(_0053_),
    .X(_0063_));
 sky130_fd_sc_hd__clkbuf_1 _0404_ (.A(_0063_),
    .X(_0205_));
 sky130_fd_sc_hd__or3_1 _0405_ (.A(_0058_),
    .B(_0059_),
    .C(_0053_),
    .X(_0064_));
 sky130_fd_sc_hd__clkbuf_1 _0406_ (.A(_0064_),
    .X(_0206_));
 sky130_fd_sc_hd__or3_1 _0407_ (.A(_0058_),
    .B(_0059_),
    .C(_0053_),
    .X(_0065_));
 sky130_fd_sc_hd__clkbuf_1 _0408_ (.A(_0065_),
    .X(_0207_));
 sky130_fd_sc_hd__clkbuf_4 _0409_ (.A(_0046_),
    .X(_0066_));
 sky130_fd_sc_hd__or3_1 _0410_ (.A(_0058_),
    .B(_0059_),
    .C(_0066_),
    .X(_0067_));
 sky130_fd_sc_hd__clkbuf_1 _0411_ (.A(_0067_),
    .X(_0208_));
 sky130_fd_sc_hd__or3_1 _0412_ (.A(_0058_),
    .B(_0059_),
    .C(_0066_),
    .X(_0068_));
 sky130_fd_sc_hd__clkbuf_1 _0413_ (.A(_0068_),
    .X(_0209_));
 sky130_fd_sc_hd__or3_1 _0414_ (.A(_0058_),
    .B(_0059_),
    .C(_0066_),
    .X(_0069_));
 sky130_fd_sc_hd__clkbuf_1 _0415_ (.A(_0069_),
    .X(_0210_));
 sky130_fd_sc_hd__or3_1 _0416_ (.A(_0058_),
    .B(_0059_),
    .C(_0066_),
    .X(_0070_));
 sky130_fd_sc_hd__clkbuf_1 _0417_ (.A(_0070_),
    .X(_0211_));
 sky130_fd_sc_hd__or3_1 _0418_ (.A(_0042_),
    .B(_0044_),
    .C(_0066_),
    .X(_0071_));
 sky130_fd_sc_hd__clkbuf_1 _0419_ (.A(_0071_),
    .X(_0212_));
 sky130_fd_sc_hd__or3_1 _0420_ (.A(_0042_),
    .B(_0044_),
    .C(_0066_),
    .X(_0072_));
 sky130_fd_sc_hd__clkbuf_1 _0421_ (.A(_0072_),
    .X(_0213_));
 sky130_fd_sc_hd__or3_1 _0422_ (.A(_0042_),
    .B(_0044_),
    .C(_0066_),
    .X(_0073_));
 sky130_fd_sc_hd__clkbuf_1 _0423_ (.A(_0073_),
    .X(_0214_));
 sky130_fd_sc_hd__or3b_1 _0424_ (.A(\zbuf_bus_sel_I[4].z ),
    .B(\zbuf_bus_sel_I[3].z ),
    .C_N(\zbuf_bus_sel_I[2].z ),
    .X(_0074_));
 sky130_fd_sc_hd__clkbuf_2 _0425_ (.A(_0074_),
    .X(_0216_));
 sky130_fd_sc_hd__buf_4 _0426_ (.A(_0042_),
    .X(_0075_));
 sky130_fd_sc_hd__buf_2 _0427_ (.A(_0046_),
    .X(_0076_));
 sky130_fd_sc_hd__buf_4 _0428_ (.A(_0044_),
    .X(_0077_));
 sky130_fd_sc_hd__or3b_1 _0429_ (.A(_0075_),
    .B(_0076_),
    .C_N(_0077_),
    .X(_0078_));
 sky130_fd_sc_hd__clkbuf_1 _0430_ (.A(_0078_),
    .X(_0217_));
 sky130_fd_sc_hd__or3b_1 _0431_ (.A(_0075_),
    .B(_0076_),
    .C_N(_0077_),
    .X(_0079_));
 sky130_fd_sc_hd__clkbuf_1 _0432_ (.A(_0079_),
    .X(_0218_));
 sky130_fd_sc_hd__or3b_1 _0433_ (.A(_0075_),
    .B(_0076_),
    .C_N(_0077_),
    .X(_0080_));
 sky130_fd_sc_hd__clkbuf_1 _0434_ (.A(_0080_),
    .X(_0219_));
 sky130_fd_sc_hd__or3b_1 _0435_ (.A(_0075_),
    .B(_0076_),
    .C_N(_0077_),
    .X(_0081_));
 sky130_fd_sc_hd__clkbuf_1 _0436_ (.A(_0081_),
    .X(_0220_));
 sky130_fd_sc_hd__or3b_1 _0437_ (.A(_0075_),
    .B(_0076_),
    .C_N(_0077_),
    .X(_0082_));
 sky130_fd_sc_hd__clkbuf_1 _0438_ (.A(_0082_),
    .X(_0221_));
 sky130_fd_sc_hd__clkbuf_2 _0439_ (.A(_0042_),
    .X(_0083_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0440_ (.A(_0044_),
    .X(_0084_));
 sky130_fd_sc_hd__or3b_1 _0441_ (.A(_0083_),
    .B(_0076_),
    .C_N(_0084_),
    .X(_0085_));
 sky130_fd_sc_hd__clkbuf_1 _0442_ (.A(_0085_),
    .X(_0222_));
 sky130_fd_sc_hd__or3b_1 _0443_ (.A(_0083_),
    .B(_0076_),
    .C_N(_0084_),
    .X(_0086_));
 sky130_fd_sc_hd__clkbuf_1 _0444_ (.A(_0086_),
    .X(_0223_));
 sky130_fd_sc_hd__or3b_1 _0445_ (.A(_0083_),
    .B(_0076_),
    .C_N(_0084_),
    .X(_0087_));
 sky130_fd_sc_hd__clkbuf_1 _0446_ (.A(_0087_),
    .X(_0224_));
 sky130_fd_sc_hd__or3b_1 _0447_ (.A(_0083_),
    .B(_0076_),
    .C_N(_0084_),
    .X(_0088_));
 sky130_fd_sc_hd__clkbuf_1 _0448_ (.A(_0088_),
    .X(_0225_));
 sky130_fd_sc_hd__clkbuf_2 _0449_ (.A(\zbuf_bus_sel_I[3].z ),
    .X(_0089_));
 sky130_fd_sc_hd__or3b_1 _0450_ (.A(_0083_),
    .B(_0089_),
    .C_N(_0084_),
    .X(_0090_));
 sky130_fd_sc_hd__clkbuf_1 _0451_ (.A(_0090_),
    .X(_0226_));
 sky130_fd_sc_hd__or3b_1 _0452_ (.A(_0083_),
    .B(_0089_),
    .C_N(_0084_),
    .X(_0091_));
 sky130_fd_sc_hd__clkbuf_1 _0453_ (.A(_0091_),
    .X(_0227_));
 sky130_fd_sc_hd__or3b_1 _0454_ (.A(_0083_),
    .B(_0089_),
    .C_N(_0084_),
    .X(_0092_));
 sky130_fd_sc_hd__clkbuf_1 _0455_ (.A(_0092_),
    .X(_0228_));
 sky130_fd_sc_hd__or3b_1 _0456_ (.A(_0083_),
    .B(_0089_),
    .C_N(_0084_),
    .X(_0093_));
 sky130_fd_sc_hd__clkbuf_1 _0457_ (.A(_0093_),
    .X(_0229_));
 sky130_fd_sc_hd__or3b_1 _0458_ (.A(_0083_),
    .B(_0089_),
    .C_N(_0084_),
    .X(_0094_));
 sky130_fd_sc_hd__clkbuf_1 _0459_ (.A(_0094_),
    .X(_0230_));
 sky130_fd_sc_hd__or3b_1 _0460_ (.A(_0083_),
    .B(_0089_),
    .C_N(_0084_),
    .X(_0095_));
 sky130_fd_sc_hd__clkbuf_1 _0461_ (.A(_0095_),
    .X(_0231_));
 sky130_fd_sc_hd__clkbuf_4 _0462_ (.A(_0042_),
    .X(_0096_));
 sky130_fd_sc_hd__clkbuf_4 _0463_ (.A(_0044_),
    .X(_0097_));
 sky130_fd_sc_hd__or3b_1 _0464_ (.A(_0096_),
    .B(_0089_),
    .C_N(_0097_),
    .X(_0098_));
 sky130_fd_sc_hd__clkbuf_1 _0465_ (.A(_0098_),
    .X(_0232_));
 sky130_fd_sc_hd__or3b_1 _0466_ (.A(_0096_),
    .B(_0089_),
    .C_N(_0097_),
    .X(_0099_));
 sky130_fd_sc_hd__clkbuf_1 _0467_ (.A(_0099_),
    .X(_0233_));
 sky130_fd_sc_hd__or3b_1 _0468_ (.A(_0096_),
    .B(_0089_),
    .C_N(_0097_),
    .X(_0100_));
 sky130_fd_sc_hd__clkbuf_1 _0469_ (.A(_0100_),
    .X(_0234_));
 sky130_fd_sc_hd__or3b_1 _0470_ (.A(_0096_),
    .B(_0089_),
    .C_N(_0097_),
    .X(_0101_));
 sky130_fd_sc_hd__clkbuf_1 _0471_ (.A(_0101_),
    .X(_0235_));
 sky130_fd_sc_hd__or3b_1 _0472_ (.A(_0096_),
    .B(_0046_),
    .C_N(_0097_),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_1 _0473_ (.A(_0102_),
    .X(_0236_));
 sky130_fd_sc_hd__or3b_1 _0474_ (.A(_0096_),
    .B(_0046_),
    .C_N(_0097_),
    .X(_0103_));
 sky130_fd_sc_hd__clkbuf_1 _0475_ (.A(_0103_),
    .X(_0237_));
 sky130_fd_sc_hd__or3b_1 _0476_ (.A(_0096_),
    .B(_0046_),
    .C_N(_0097_),
    .X(_0104_));
 sky130_fd_sc_hd__clkbuf_1 _0477_ (.A(_0104_),
    .X(_0238_));
 sky130_fd_sc_hd__or3b_1 _0478_ (.A(\zbuf_bus_sel_I[4].z ),
    .B(\zbuf_bus_sel_I[2].z ),
    .C_N(\zbuf_bus_sel_I[3].z ),
    .X(_0105_));
 sky130_fd_sc_hd__clkbuf_2 _0479_ (.A(_0105_),
    .X(_0240_));
 sky130_fd_sc_hd__or3b_1 _0480_ (.A(_0096_),
    .B(_0097_),
    .C_N(_0066_),
    .X(_0106_));
 sky130_fd_sc_hd__clkbuf_1 _0481_ (.A(_0106_),
    .X(_0241_));
 sky130_fd_sc_hd__or3b_1 _0482_ (.A(_0096_),
    .B(_0097_),
    .C_N(_0066_),
    .X(_0107_));
 sky130_fd_sc_hd__clkbuf_1 _0483_ (.A(_0107_),
    .X(_0242_));
 sky130_fd_sc_hd__clkbuf_2 _0484_ (.A(_0044_),
    .X(_0108_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0485_ (.A(_0046_),
    .X(_0109_));
 sky130_fd_sc_hd__or3b_1 _0486_ (.A(_0096_),
    .B(_0108_),
    .C_N(_0109_),
    .X(_0110_));
 sky130_fd_sc_hd__clkbuf_1 _0487_ (.A(_0110_),
    .X(_0243_));
 sky130_fd_sc_hd__clkbuf_2 _0488_ (.A(_0042_),
    .X(_0111_));
 sky130_fd_sc_hd__or3b_1 _0489_ (.A(_0111_),
    .B(_0108_),
    .C_N(_0109_),
    .X(_0112_));
 sky130_fd_sc_hd__clkbuf_1 _0490_ (.A(_0112_),
    .X(_0244_));
 sky130_fd_sc_hd__or3b_1 _0491_ (.A(_0111_),
    .B(_0108_),
    .C_N(_0109_),
    .X(_0113_));
 sky130_fd_sc_hd__clkbuf_1 _0492_ (.A(_0113_),
    .X(_0245_));
 sky130_fd_sc_hd__or3b_1 _0493_ (.A(_0111_),
    .B(_0108_),
    .C_N(_0109_),
    .X(_0114_));
 sky130_fd_sc_hd__clkbuf_1 _0494_ (.A(_0114_),
    .X(_0246_));
 sky130_fd_sc_hd__or3b_1 _0495_ (.A(_0111_),
    .B(_0108_),
    .C_N(_0109_),
    .X(_0115_));
 sky130_fd_sc_hd__clkbuf_1 _0496_ (.A(_0115_),
    .X(_0247_));
 sky130_fd_sc_hd__or3b_1 _0497_ (.A(_0111_),
    .B(_0108_),
    .C_N(_0109_),
    .X(_0116_));
 sky130_fd_sc_hd__clkbuf_1 _0498_ (.A(_0116_),
    .X(_0248_));
 sky130_fd_sc_hd__or3b_1 _0499_ (.A(_0111_),
    .B(_0108_),
    .C_N(_0109_),
    .X(_0117_));
 sky130_fd_sc_hd__clkbuf_1 _0500_ (.A(_0117_),
    .X(_0249_));
 sky130_fd_sc_hd__or3b_1 _0501_ (.A(_0111_),
    .B(_0108_),
    .C_N(_0109_),
    .X(_0118_));
 sky130_fd_sc_hd__clkbuf_1 _0502_ (.A(_0118_),
    .X(_0250_));
 sky130_fd_sc_hd__or3b_1 _0503_ (.A(_0111_),
    .B(_0108_),
    .C_N(_0109_),
    .X(_0119_));
 sky130_fd_sc_hd__clkbuf_1 _0504_ (.A(_0119_),
    .X(_0251_));
 sky130_fd_sc_hd__or3b_1 _0505_ (.A(_0111_),
    .B(_0108_),
    .C_N(_0109_),
    .X(_0120_));
 sky130_fd_sc_hd__clkbuf_1 _0506_ (.A(_0120_),
    .X(_0252_));
 sky130_fd_sc_hd__clkbuf_2 _0507_ (.A(\zbuf_bus_sel_I[2].z ),
    .X(_0121_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0508_ (.A(_0046_),
    .X(_0122_));
 sky130_fd_sc_hd__or3b_1 _0509_ (.A(_0111_),
    .B(_0121_),
    .C_N(_0122_),
    .X(_0123_));
 sky130_fd_sc_hd__clkbuf_1 _0510_ (.A(_0123_),
    .X(_0253_));
 sky130_fd_sc_hd__clkbuf_2 _0511_ (.A(_0042_),
    .X(_0124_));
 sky130_fd_sc_hd__or3b_1 _0512_ (.A(_0124_),
    .B(_0121_),
    .C_N(_0122_),
    .X(_0125_));
 sky130_fd_sc_hd__clkbuf_1 _0513_ (.A(_0125_),
    .X(_0254_));
 sky130_fd_sc_hd__or3b_1 _0514_ (.A(_0124_),
    .B(_0121_),
    .C_N(_0122_),
    .X(_0126_));
 sky130_fd_sc_hd__clkbuf_1 _0515_ (.A(_0126_),
    .X(_0255_));
 sky130_fd_sc_hd__or3b_1 _0516_ (.A(_0124_),
    .B(_0121_),
    .C_N(_0122_),
    .X(_0127_));
 sky130_fd_sc_hd__clkbuf_1 _0517_ (.A(_0127_),
    .X(_0256_));
 sky130_fd_sc_hd__or3b_1 _0518_ (.A(_0124_),
    .B(_0121_),
    .C_N(_0122_),
    .X(_0128_));
 sky130_fd_sc_hd__clkbuf_1 _0519_ (.A(_0128_),
    .X(_0257_));
 sky130_fd_sc_hd__or3b_1 _0520_ (.A(_0124_),
    .B(_0121_),
    .C_N(_0122_),
    .X(_0129_));
 sky130_fd_sc_hd__clkbuf_1 _0521_ (.A(_0129_),
    .X(_0258_));
 sky130_fd_sc_hd__or3b_1 _0522_ (.A(_0124_),
    .B(_0121_),
    .C_N(_0122_),
    .X(_0130_));
 sky130_fd_sc_hd__clkbuf_1 _0523_ (.A(_0130_),
    .X(_0259_));
 sky130_fd_sc_hd__or3b_1 _0524_ (.A(_0124_),
    .B(_0121_),
    .C_N(_0122_),
    .X(_0131_));
 sky130_fd_sc_hd__clkbuf_1 _0525_ (.A(_0131_),
    .X(_0260_));
 sky130_fd_sc_hd__or3b_1 _0526_ (.A(_0124_),
    .B(_0121_),
    .C_N(_0122_),
    .X(_0132_));
 sky130_fd_sc_hd__clkbuf_1 _0527_ (.A(_0132_),
    .X(_0261_));
 sky130_fd_sc_hd__or3b_1 _0528_ (.A(_0124_),
    .B(_0121_),
    .C_N(_0122_),
    .X(_0133_));
 sky130_fd_sc_hd__clkbuf_1 _0529_ (.A(_0133_),
    .X(_0262_));
 sky130_fd_sc_hd__nand3b_4 _0530_ (.A_N(\zbuf_bus_sel_I[4].z ),
    .B(\zbuf_bus_sel_I[2].z ),
    .C(\zbuf_bus_sel_I[3].z ),
    .Y(_0264_));
 sky130_fd_sc_hd__clkbuf_2 _0531_ (.A(_0075_),
    .X(_0134_));
 sky130_fd_sc_hd__clkbuf_4 _0532_ (.A(_0077_),
    .X(_0135_));
 sky130_fd_sc_hd__clkbuf_4 _0533_ (.A(_0047_),
    .X(_0136_));
 sky130_fd_sc_hd__nand3b_2 _0534_ (.A_N(_0134_),
    .B(_0135_),
    .C(_0136_),
    .Y(_0265_));
 sky130_fd_sc_hd__nand3b_2 _0535_ (.A_N(_0134_),
    .B(_0135_),
    .C(_0136_),
    .Y(_0266_));
 sky130_fd_sc_hd__nand3b_2 _0536_ (.A_N(_0134_),
    .B(_0135_),
    .C(_0136_),
    .Y(_0267_));
 sky130_fd_sc_hd__nand3b_1 _0537_ (.A_N(_0134_),
    .B(_0135_),
    .C(_0136_),
    .Y(_0268_));
 sky130_fd_sc_hd__nand3b_1 _0538_ (.A_N(_0134_),
    .B(_0135_),
    .C(_0136_),
    .Y(_0269_));
 sky130_fd_sc_hd__nand3b_2 _0539_ (.A_N(_0134_),
    .B(_0135_),
    .C(_0136_),
    .Y(_0270_));
 sky130_fd_sc_hd__nand3b_1 _0540_ (.A_N(_0134_),
    .B(_0135_),
    .C(_0136_),
    .Y(_0271_));
 sky130_fd_sc_hd__nand3b_1 _0541_ (.A_N(_0134_),
    .B(_0135_),
    .C(_0136_),
    .Y(_0272_));
 sky130_fd_sc_hd__nand3b_1 _0542_ (.A_N(_0134_),
    .B(_0135_),
    .C(_0136_),
    .Y(_0273_));
 sky130_fd_sc_hd__nand3b_1 _0543_ (.A_N(_0134_),
    .B(_0135_),
    .C(_0136_),
    .Y(_0274_));
 sky130_fd_sc_hd__clkbuf_2 _0544_ (.A(_0075_),
    .X(_0137_));
 sky130_fd_sc_hd__clkbuf_4 _0545_ (.A(_0077_),
    .X(_0138_));
 sky130_fd_sc_hd__clkbuf_4 _0546_ (.A(_0047_),
    .X(_0139_));
 sky130_fd_sc_hd__nand3b_2 _0547_ (.A_N(_0137_),
    .B(_0138_),
    .C(_0139_),
    .Y(_0275_));
 sky130_fd_sc_hd__nand3b_2 _0548_ (.A_N(_0137_),
    .B(_0138_),
    .C(_0139_),
    .Y(_0276_));
 sky130_fd_sc_hd__nand3b_2 _0549_ (.A_N(_0137_),
    .B(_0138_),
    .C(_0139_),
    .Y(_0277_));
 sky130_fd_sc_hd__nand3b_2 _0550_ (.A_N(_0137_),
    .B(_0138_),
    .C(_0139_),
    .Y(_0278_));
 sky130_fd_sc_hd__nand3b_2 _0551_ (.A_N(_0137_),
    .B(_0138_),
    .C(_0139_),
    .Y(_0279_));
 sky130_fd_sc_hd__nand3b_2 _0552_ (.A_N(_0137_),
    .B(_0138_),
    .C(_0139_),
    .Y(_0280_));
 sky130_fd_sc_hd__nand3b_2 _0553_ (.A_N(_0137_),
    .B(_0138_),
    .C(_0139_),
    .Y(_0281_));
 sky130_fd_sc_hd__nand3b_2 _0554_ (.A_N(_0137_),
    .B(_0138_),
    .C(_0139_),
    .Y(_0282_));
 sky130_fd_sc_hd__nand3b_1 _0555_ (.A_N(_0137_),
    .B(_0138_),
    .C(_0139_),
    .Y(_0283_));
 sky130_fd_sc_hd__nand3b_1 _0556_ (.A_N(_0137_),
    .B(_0138_),
    .C(_0139_),
    .Y(_0284_));
 sky130_fd_sc_hd__nand3b_1 _0557_ (.A_N(_0075_),
    .B(_0077_),
    .C(_0047_),
    .Y(_0285_));
 sky130_fd_sc_hd__nand3b_1 _0558_ (.A_N(_0075_),
    .B(_0077_),
    .C(_0047_),
    .Y(_0286_));
 sky130_fd_sc_hd__or4_1 _0559_ (.A(_0001_),
    .B(_0005_),
    .C(_0008_),
    .D(_0012_),
    .X(_0140_));
 sky130_fd_sc_hd__clkbuf_1 _0560_ (.A(_0140_),
    .X(_0167_));
 sky130_fd_sc_hd__nand3b_2 _0561_ (.A_N(_0075_),
    .B(_0077_),
    .C(_0047_),
    .Y(_0263_));
 sky130_fd_sc_hd__or3b_1 _0562_ (.A(_0124_),
    .B(_0045_),
    .C_N(_0076_),
    .X(_0141_));
 sky130_fd_sc_hd__clkbuf_1 _0563_ (.A(_0141_),
    .X(_0239_));
 sky130_fd_sc_hd__or3b_1 _0564_ (.A(_0043_),
    .B(_0046_),
    .C_N(_0097_),
    .X(_0142_));
 sky130_fd_sc_hd__clkbuf_1 _0565_ (.A(_0142_),
    .X(_0215_));
 sky130_fd_sc_hd__or3_1 _0566_ (.A(_0042_),
    .B(_0044_),
    .C(_0066_),
    .X(_0143_));
 sky130_fd_sc_hd__clkbuf_1 _0567_ (.A(_0143_),
    .X(_0191_));
 sky130_fd_sc_hd__or4b_4 _0568_ (.A(net469),
    .B(net455),
    .C(_0192_),
    .D_N(\zbuf_bus_ena_I.z ),
    .X(_0144_));
 sky130_fd_sc_hd__inv_2 _0569_ (.A(_0144_),
    .Y(\col[0].zbuf_bot_ena_I.e ));
 sky130_fd_sc_hd__buf_4 _0570_ (.A(net458),
    .X(_0145_));
 sky130_fd_sc_hd__inv_2 _0571_ (.A(_0192_),
    .Y(_0146_));
 sky130_fd_sc_hd__buf_4 _0572_ (.A(net471),
    .X(_0147_));
 sky130_fd_sc_hd__buf_4 _0573_ (.A(\zbuf_bus_ena_I.z ),
    .X(_0148_));
 sky130_fd_sc_hd__and4b_2 _0574_ (.A_N(_0145_),
    .B(_0146_),
    .C(_0147_),
    .D(_0148_),
    .X(_0149_));
 sky130_fd_sc_hd__clkbuf_2 _0575_ (.A(_0149_),
    .X(\col[0].zbuf_top_ena_I.e ));
 sky130_fd_sc_hd__and4b_2 _0576_ (.A_N(_0147_),
    .B(_0148_),
    .C(_0145_),
    .D(_0146_),
    .X(_0150_));
 sky130_fd_sc_hd__clkbuf_1 _0577_ (.A(_0150_),
    .X(\col[1].zbuf_bot_ena_I.e ));
 sky130_fd_sc_hd__and4_2 _0578_ (.A(_0147_),
    .B(_0148_),
    .C(_0145_),
    .D(_0146_),
    .X(_0151_));
 sky130_fd_sc_hd__clkbuf_1 _0579_ (.A(_0151_),
    .X(\col[1].zbuf_top_ena_I.e ));
 sky130_fd_sc_hd__or4b_2 _0580_ (.A(net468),
    .B(net455),
    .C(_0216_),
    .D_N(\zbuf_bus_ena_I.z ),
    .X(_0152_));
 sky130_fd_sc_hd__inv_2 _0581_ (.A(_0152_),
    .Y(\col[2].zbuf_bot_ena_I.e ));
 sky130_fd_sc_hd__inv_2 _0582_ (.A(_0216_),
    .Y(_0153_));
 sky130_fd_sc_hd__and4b_1 _0583_ (.A_N(_0145_),
    .B(_0153_),
    .C(_0147_),
    .D(_0148_),
    .X(_0154_));
 sky130_fd_sc_hd__clkbuf_1 _0584_ (.A(_0154_),
    .X(\col[2].zbuf_top_ena_I.e ));
 sky130_fd_sc_hd__and4b_1 _0585_ (.A_N(_0147_),
    .B(_0148_),
    .C(_0145_),
    .D(_0153_),
    .X(_0155_));
 sky130_fd_sc_hd__clkbuf_1 _0586_ (.A(_0155_),
    .X(\col[3].zbuf_bot_ena_I.e ));
 sky130_fd_sc_hd__and4_1 _0587_ (.A(_0147_),
    .B(_0148_),
    .C(_0145_),
    .D(_0153_),
    .X(_0156_));
 sky130_fd_sc_hd__clkbuf_1 _0588_ (.A(_0156_),
    .X(\col[3].zbuf_top_ena_I.e ));
 sky130_fd_sc_hd__or4b_1 _0589_ (.A(net472),
    .B(net459),
    .C(_0240_),
    .D_N(\zbuf_bus_ena_I.z ),
    .X(_0157_));
 sky130_fd_sc_hd__inv_2 _0590_ (.A(_0157_),
    .Y(\col[4].zbuf_bot_ena_I.e ));
 sky130_fd_sc_hd__inv_2 _0591_ (.A(_0240_),
    .Y(_0158_));
 sky130_fd_sc_hd__and4b_1 _0592_ (.A_N(_0145_),
    .B(_0158_),
    .C(net472),
    .D(\zbuf_bus_ena_I.z ),
    .X(_0159_));
 sky130_fd_sc_hd__clkbuf_1 _0593_ (.A(_0159_),
    .X(\col[4].zbuf_top_ena_I.e ));
 sky130_fd_sc_hd__and4b_1 _0594_ (.A_N(_0147_),
    .B(_0148_),
    .C(_0145_),
    .D(_0158_),
    .X(_0160_));
 sky130_fd_sc_hd__clkbuf_1 _0595_ (.A(_0160_),
    .X(\col[5].zbuf_bot_ena_I.e ));
 sky130_fd_sc_hd__and4_1 _0596_ (.A(_0147_),
    .B(_0148_),
    .C(net463),
    .D(_0158_),
    .X(_0161_));
 sky130_fd_sc_hd__clkbuf_1 _0597_ (.A(_0161_),
    .X(\col[5].zbuf_top_ena_I.e ));
 sky130_fd_sc_hd__or4b_1 _0598_ (.A(net474),
    .B(net460),
    .C(_0264_),
    .D_N(\zbuf_bus_ena_I.z ),
    .X(_0162_));
 sky130_fd_sc_hd__inv_2 _0599_ (.A(_0162_),
    .Y(\col[6].zbuf_bot_ena_I.e ));
 sky130_fd_sc_hd__inv_2 _0600_ (.A(_0264_),
    .Y(_0163_));
 sky130_fd_sc_hd__and4b_1 _0601_ (.A_N(_0145_),
    .B(_0163_),
    .C(net474),
    .D(\zbuf_bus_ena_I.z ),
    .X(_0164_));
 sky130_fd_sc_hd__clkbuf_1 _0602_ (.A(_0164_),
    .X(\col[6].zbuf_top_ena_I.e ));
 sky130_fd_sc_hd__and4b_1 _0603_ (.A_N(_0147_),
    .B(_0148_),
    .C(_0145_),
    .D(_0163_),
    .X(_0165_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0604_ (.A(_0165_),
    .X(\col[7].zbuf_bot_ena_I.e ));
 sky130_fd_sc_hd__and4_1 _0605_ (.A(_0147_),
    .B(_0148_),
    .C(net461),
    .D(_0163_),
    .X(_0166_));
 sky130_fd_sc_hd__clkbuf_2 _0606_ (.A(_0166_),
    .X(\col[7].zbuf_top_ena_I.e ));
 sky130_fd_sc_hd__buf_2 _0643_ (.A(\col[1].zbuf_bot_iw_I[4].z ),
    .X(um_iw[40]));
 sky130_fd_sc_hd__buf_2 _0644_ (.A(\col[1].zbuf_bot_iw_I[5].z ),
    .X(um_iw[41]));
 sky130_fd_sc_hd__buf_2 _0645_ (.A(\col[1].zbuf_bot_iw_I[6].z ),
    .X(um_iw[42]));
 sky130_fd_sc_hd__buf_2 _0646_ (.A(\col[1].zbuf_bot_iw_I[7].z ),
    .X(um_iw[43]));
 sky130_fd_sc_hd__buf_2 _0647_ (.A(\col[1].zbuf_bot_iw_I[8].z ),
    .X(um_iw[44]));
 sky130_fd_sc_hd__buf_2 _0648_ (.A(\col[1].zbuf_bot_iw_I[9].z ),
    .X(um_iw[45]));
 sky130_fd_sc_hd__buf_2 _0649_ (.A(\col[1].zbuf_bot_iw_I[10].z ),
    .X(um_iw[46]));
 sky130_fd_sc_hd__buf_2 _0650_ (.A(\col[1].zbuf_bot_iw_I[11].z ),
    .X(um_iw[47]));
 sky130_fd_sc_hd__buf_2 _0651_ (.A(\col[1].zbuf_bot_iw_I[12].z ),
    .X(um_iw[48]));
 sky130_fd_sc_hd__buf_2 _0652_ (.A(\col[1].zbuf_bot_iw_I[13].z ),
    .X(um_iw[49]));
 sky130_fd_sc_hd__buf_2 _0653_ (.A(\col[1].zbuf_bot_iw_I[14].z ),
    .X(um_iw[50]));
 sky130_fd_sc_hd__buf_2 _0654_ (.A(\col[1].zbuf_bot_iw_I[15].z ),
    .X(um_iw[51]));
 sky130_fd_sc_hd__buf_2 _0655_ (.A(\col[1].zbuf_bot_iw_I[16].z ),
    .X(um_iw[52]));
 sky130_fd_sc_hd__buf_2 _0656_ (.A(\col[1].zbuf_bot_iw_I[17].z ),
    .X(um_iw[53]));
 sky130_fd_sc_hd__buf_2 _0657_ (.A(\col[1].zbuf_top_iw_I[0].z ),
    .X(um_iw[54]));
 sky130_fd_sc_hd__buf_2 _0658_ (.A(\col[1].zbuf_top_iw_I[1].z ),
    .X(um_iw[55]));
 sky130_fd_sc_hd__buf_2 _0659_ (.A(\col[1].zbuf_top_iw_I[2].z ),
    .X(um_iw[56]));
 sky130_fd_sc_hd__buf_2 _0660_ (.A(\col[1].zbuf_top_iw_I[3].z ),
    .X(um_iw[57]));
 sky130_fd_sc_hd__buf_2 _0661_ (.A(\col[1].zbuf_top_iw_I[4].z ),
    .X(um_iw[58]));
 sky130_fd_sc_hd__buf_2 _0662_ (.A(\col[1].zbuf_top_iw_I[5].z ),
    .X(um_iw[59]));
 sky130_fd_sc_hd__buf_2 _0663_ (.A(\col[1].zbuf_top_iw_I[6].z ),
    .X(um_iw[60]));
 sky130_fd_sc_hd__buf_2 _0664_ (.A(\col[1].zbuf_top_iw_I[7].z ),
    .X(um_iw[61]));
 sky130_fd_sc_hd__buf_2 _0665_ (.A(\col[1].zbuf_top_iw_I[8].z ),
    .X(um_iw[62]));
 sky130_fd_sc_hd__buf_2 _0666_ (.A(\col[1].zbuf_top_iw_I[9].z ),
    .X(um_iw[63]));
 sky130_fd_sc_hd__buf_2 _0667_ (.A(\col[1].zbuf_top_iw_I[10].z ),
    .X(um_iw[64]));
 sky130_fd_sc_hd__buf_2 _0668_ (.A(\col[1].zbuf_top_iw_I[11].z ),
    .X(um_iw[65]));
 sky130_fd_sc_hd__buf_2 _0669_ (.A(\col[1].zbuf_top_iw_I[12].z ),
    .X(um_iw[66]));
 sky130_fd_sc_hd__buf_2 _0670_ (.A(\col[1].zbuf_top_iw_I[13].z ),
    .X(um_iw[67]));
 sky130_fd_sc_hd__buf_2 _0671_ (.A(\col[1].zbuf_top_iw_I[14].z ),
    .X(um_iw[68]));
 sky130_fd_sc_hd__buf_2 _0672_ (.A(\col[1].zbuf_top_iw_I[15].z ),
    .X(um_iw[69]));
 sky130_fd_sc_hd__buf_2 _0673_ (.A(\col[1].zbuf_top_iw_I[16].z ),
    .X(um_iw[70]));
 sky130_fd_sc_hd__buf_2 _0674_ (.A(\col[1].zbuf_top_iw_I[17].z ),
    .X(um_iw[71]));
 sky130_fd_sc_hd__buf_2 _0675_ (.A(\col[2].zbuf_bot_iw_I[0].z ),
    .X(um_iw[72]));
 sky130_fd_sc_hd__buf_2 _0676_ (.A(\col[2].zbuf_bot_iw_I[1].z ),
    .X(um_iw[73]));
 sky130_fd_sc_hd__buf_2 _0677_ (.A(\col[2].zbuf_bot_iw_I[2].z ),
    .X(um_iw[74]));
 sky130_fd_sc_hd__buf_2 _0678_ (.A(\col[2].zbuf_bot_iw_I[3].z ),
    .X(um_iw[75]));
 sky130_fd_sc_hd__buf_2 _0679_ (.A(\col[2].zbuf_bot_iw_I[4].z ),
    .X(um_iw[76]));
 sky130_fd_sc_hd__buf_2 _0680_ (.A(\col[2].zbuf_bot_iw_I[5].z ),
    .X(um_iw[77]));
 sky130_fd_sc_hd__buf_2 _0681_ (.A(\col[2].zbuf_bot_iw_I[6].z ),
    .X(um_iw[78]));
 sky130_fd_sc_hd__buf_2 _0682_ (.A(\col[2].zbuf_bot_iw_I[7].z ),
    .X(um_iw[79]));
 sky130_fd_sc_hd__buf_2 _0683_ (.A(\col[2].zbuf_bot_iw_I[8].z ),
    .X(um_iw[80]));
 sky130_fd_sc_hd__buf_2 _0684_ (.A(\col[2].zbuf_bot_iw_I[9].z ),
    .X(um_iw[81]));
 sky130_fd_sc_hd__buf_2 _0685_ (.A(\col[2].zbuf_bot_iw_I[10].z ),
    .X(um_iw[82]));
 sky130_fd_sc_hd__buf_2 _0686_ (.A(\col[2].zbuf_bot_iw_I[11].z ),
    .X(um_iw[83]));
 sky130_fd_sc_hd__buf_2 _0687_ (.A(\col[2].zbuf_bot_iw_I[12].z ),
    .X(um_iw[84]));
 sky130_fd_sc_hd__buf_2 _0688_ (.A(\col[2].zbuf_bot_iw_I[13].z ),
    .X(um_iw[85]));
 sky130_fd_sc_hd__buf_2 _0689_ (.A(\col[2].zbuf_bot_iw_I[14].z ),
    .X(um_iw[86]));
 sky130_fd_sc_hd__buf_2 _0690_ (.A(\col[2].zbuf_bot_iw_I[15].z ),
    .X(um_iw[87]));
 sky130_fd_sc_hd__buf_2 _0691_ (.A(\col[2].zbuf_bot_iw_I[16].z ),
    .X(um_iw[88]));
 sky130_fd_sc_hd__buf_2 _0692_ (.A(\col[2].zbuf_bot_iw_I[17].z ),
    .X(um_iw[89]));
 sky130_fd_sc_hd__buf_2 _0693_ (.A(\col[2].zbuf_top_iw_I[0].z ),
    .X(um_iw[90]));
 sky130_fd_sc_hd__buf_2 _0694_ (.A(\col[2].zbuf_top_iw_I[1].z ),
    .X(um_iw[91]));
 sky130_fd_sc_hd__buf_2 _0695_ (.A(\col[2].zbuf_top_iw_I[2].z ),
    .X(um_iw[92]));
 sky130_fd_sc_hd__buf_2 _0696_ (.A(\col[2].zbuf_top_iw_I[3].z ),
    .X(um_iw[93]));
 sky130_fd_sc_hd__buf_2 _0697_ (.A(\col[2].zbuf_top_iw_I[4].z ),
    .X(um_iw[94]));
 sky130_fd_sc_hd__buf_2 _0698_ (.A(\col[2].zbuf_top_iw_I[5].z ),
    .X(um_iw[95]));
 sky130_fd_sc_hd__buf_2 _0699_ (.A(\col[2].zbuf_top_iw_I[6].z ),
    .X(um_iw[96]));
 sky130_fd_sc_hd__buf_2 _0700_ (.A(\col[2].zbuf_top_iw_I[7].z ),
    .X(um_iw[97]));
 sky130_fd_sc_hd__buf_2 _0701_ (.A(\col[2].zbuf_top_iw_I[8].z ),
    .X(um_iw[98]));
 sky130_fd_sc_hd__buf_2 _0702_ (.A(\col[2].zbuf_top_iw_I[9].z ),
    .X(um_iw[99]));
 sky130_fd_sc_hd__buf_2 _0703_ (.A(\col[2].zbuf_top_iw_I[10].z ),
    .X(um_iw[100]));
 sky130_fd_sc_hd__buf_2 _0704_ (.A(\col[2].zbuf_top_iw_I[11].z ),
    .X(um_iw[101]));
 sky130_fd_sc_hd__buf_2 _0705_ (.A(\col[2].zbuf_top_iw_I[12].z ),
    .X(um_iw[102]));
 sky130_fd_sc_hd__buf_2 _0706_ (.A(\col[2].zbuf_top_iw_I[13].z ),
    .X(um_iw[103]));
 sky130_fd_sc_hd__buf_2 _0707_ (.A(\col[2].zbuf_top_iw_I[14].z ),
    .X(um_iw[104]));
 sky130_fd_sc_hd__buf_2 _0708_ (.A(\col[2].zbuf_top_iw_I[15].z ),
    .X(um_iw[105]));
 sky130_fd_sc_hd__buf_2 _0709_ (.A(\col[2].zbuf_top_iw_I[16].z ),
    .X(um_iw[106]));
 sky130_fd_sc_hd__buf_2 _0710_ (.A(\col[2].zbuf_top_iw_I[17].z ),
    .X(um_iw[107]));
 sky130_fd_sc_hd__buf_2 _0711_ (.A(\col[3].zbuf_bot_iw_I[0].z ),
    .X(um_iw[108]));
 sky130_fd_sc_hd__buf_2 _0712_ (.A(\col[3].zbuf_bot_iw_I[1].z ),
    .X(um_iw[109]));
 sky130_fd_sc_hd__buf_2 _0713_ (.A(\col[3].zbuf_bot_iw_I[2].z ),
    .X(um_iw[110]));
 sky130_fd_sc_hd__buf_2 _0714_ (.A(\col[3].zbuf_bot_iw_I[3].z ),
    .X(um_iw[111]));
 sky130_fd_sc_hd__buf_2 _0715_ (.A(\col[3].zbuf_bot_iw_I[4].z ),
    .X(um_iw[112]));
 sky130_fd_sc_hd__buf_2 _0716_ (.A(\col[3].zbuf_bot_iw_I[5].z ),
    .X(um_iw[113]));
 sky130_fd_sc_hd__buf_2 _0717_ (.A(\col[3].zbuf_bot_iw_I[6].z ),
    .X(um_iw[114]));
 sky130_fd_sc_hd__buf_2 _0718_ (.A(\col[3].zbuf_bot_iw_I[7].z ),
    .X(um_iw[115]));
 sky130_fd_sc_hd__buf_2 _0719_ (.A(\col[3].zbuf_bot_iw_I[8].z ),
    .X(um_iw[116]));
 sky130_fd_sc_hd__buf_2 _0720_ (.A(\col[3].zbuf_bot_iw_I[9].z ),
    .X(um_iw[117]));
 sky130_fd_sc_hd__buf_2 _0721_ (.A(\col[3].zbuf_bot_iw_I[10].z ),
    .X(um_iw[118]));
 sky130_fd_sc_hd__buf_2 _0722_ (.A(\col[3].zbuf_bot_iw_I[11].z ),
    .X(um_iw[119]));
 sky130_fd_sc_hd__buf_2 _0723_ (.A(\col[3].zbuf_bot_iw_I[12].z ),
    .X(um_iw[120]));
 sky130_fd_sc_hd__buf_2 _0724_ (.A(\col[3].zbuf_bot_iw_I[13].z ),
    .X(um_iw[121]));
 sky130_fd_sc_hd__buf_2 _0725_ (.A(\col[3].zbuf_bot_iw_I[14].z ),
    .X(um_iw[122]));
 sky130_fd_sc_hd__buf_2 _0726_ (.A(\col[3].zbuf_bot_iw_I[15].z ),
    .X(um_iw[123]));
 sky130_fd_sc_hd__buf_2 _0727_ (.A(\col[3].zbuf_bot_iw_I[16].z ),
    .X(um_iw[124]));
 sky130_fd_sc_hd__buf_2 _0728_ (.A(\col[3].zbuf_bot_iw_I[17].z ),
    .X(um_iw[125]));
 sky130_fd_sc_hd__buf_2 _0729_ (.A(\col[3].zbuf_top_iw_I[0].z ),
    .X(um_iw[126]));
 sky130_fd_sc_hd__buf_2 _0730_ (.A(\col[3].zbuf_top_iw_I[1].z ),
    .X(um_iw[127]));
 sky130_fd_sc_hd__buf_2 _0731_ (.A(\col[3].zbuf_top_iw_I[2].z ),
    .X(um_iw[128]));
 sky130_fd_sc_hd__buf_2 _0732_ (.A(\col[3].zbuf_top_iw_I[3].z ),
    .X(um_iw[129]));
 sky130_fd_sc_hd__buf_2 _0733_ (.A(\col[3].zbuf_top_iw_I[4].z ),
    .X(um_iw[130]));
 sky130_fd_sc_hd__buf_2 _0734_ (.A(\col[3].zbuf_top_iw_I[5].z ),
    .X(um_iw[131]));
 sky130_fd_sc_hd__buf_2 _0735_ (.A(\col[3].zbuf_top_iw_I[6].z ),
    .X(um_iw[132]));
 sky130_fd_sc_hd__buf_2 _0736_ (.A(\col[3].zbuf_top_iw_I[7].z ),
    .X(um_iw[133]));
 sky130_fd_sc_hd__buf_2 _0737_ (.A(\col[3].zbuf_top_iw_I[8].z ),
    .X(um_iw[134]));
 sky130_fd_sc_hd__buf_2 _0738_ (.A(\col[3].zbuf_top_iw_I[9].z ),
    .X(um_iw[135]));
 sky130_fd_sc_hd__buf_2 _0739_ (.A(\col[3].zbuf_top_iw_I[10].z ),
    .X(um_iw[136]));
 sky130_fd_sc_hd__buf_2 _0740_ (.A(\col[3].zbuf_top_iw_I[11].z ),
    .X(um_iw[137]));
 sky130_fd_sc_hd__buf_2 _0741_ (.A(\col[3].zbuf_top_iw_I[12].z ),
    .X(um_iw[138]));
 sky130_fd_sc_hd__buf_2 _0742_ (.A(\col[3].zbuf_top_iw_I[13].z ),
    .X(um_iw[139]));
 sky130_fd_sc_hd__buf_2 _0743_ (.A(\col[3].zbuf_top_iw_I[14].z ),
    .X(um_iw[140]));
 sky130_fd_sc_hd__buf_2 _0744_ (.A(\col[3].zbuf_top_iw_I[15].z ),
    .X(um_iw[141]));
 sky130_fd_sc_hd__buf_2 _0745_ (.A(\col[3].zbuf_top_iw_I[16].z ),
    .X(um_iw[142]));
 sky130_fd_sc_hd__buf_2 _0746_ (.A(\col[3].zbuf_top_iw_I[17].z ),
    .X(um_iw[143]));
 sky130_fd_sc_hd__buf_2 _0747_ (.A(\col[4].zbuf_bot_iw_I[0].z ),
    .X(um_iw[144]));
 sky130_fd_sc_hd__buf_2 _0748_ (.A(\col[4].zbuf_bot_iw_I[1].z ),
    .X(um_iw[145]));
 sky130_fd_sc_hd__buf_2 _0749_ (.A(\col[4].zbuf_bot_iw_I[2].z ),
    .X(um_iw[146]));
 sky130_fd_sc_hd__buf_2 _0750_ (.A(\col[4].zbuf_bot_iw_I[3].z ),
    .X(um_iw[147]));
 sky130_fd_sc_hd__buf_2 _0751_ (.A(\col[4].zbuf_bot_iw_I[4].z ),
    .X(um_iw[148]));
 sky130_fd_sc_hd__buf_2 _0752_ (.A(\col[4].zbuf_bot_iw_I[5].z ),
    .X(um_iw[149]));
 sky130_fd_sc_hd__buf_2 _0753_ (.A(\col[4].zbuf_bot_iw_I[6].z ),
    .X(um_iw[150]));
 sky130_fd_sc_hd__buf_2 _0754_ (.A(\col[4].zbuf_bot_iw_I[7].z ),
    .X(um_iw[151]));
 sky130_fd_sc_hd__buf_2 _0755_ (.A(\col[4].zbuf_bot_iw_I[8].z ),
    .X(um_iw[152]));
 sky130_fd_sc_hd__buf_2 _0756_ (.A(\col[4].zbuf_bot_iw_I[9].z ),
    .X(um_iw[153]));
 sky130_fd_sc_hd__buf_2 _0757_ (.A(\col[4].zbuf_bot_iw_I[10].z ),
    .X(um_iw[154]));
 sky130_fd_sc_hd__buf_2 _0758_ (.A(\col[4].zbuf_bot_iw_I[11].z ),
    .X(um_iw[155]));
 sky130_fd_sc_hd__buf_2 _0759_ (.A(\col[4].zbuf_bot_iw_I[12].z ),
    .X(um_iw[156]));
 sky130_fd_sc_hd__buf_2 _0760_ (.A(\col[4].zbuf_bot_iw_I[13].z ),
    .X(um_iw[157]));
 sky130_fd_sc_hd__buf_2 _0761_ (.A(\col[4].zbuf_bot_iw_I[14].z ),
    .X(um_iw[158]));
 sky130_fd_sc_hd__buf_2 _0762_ (.A(\col[4].zbuf_bot_iw_I[15].z ),
    .X(um_iw[159]));
 sky130_fd_sc_hd__buf_2 _0763_ (.A(\col[4].zbuf_bot_iw_I[16].z ),
    .X(um_iw[160]));
 sky130_fd_sc_hd__buf_2 _0764_ (.A(\col[4].zbuf_bot_iw_I[17].z ),
    .X(um_iw[161]));
 sky130_fd_sc_hd__buf_2 _0765_ (.A(\col[4].zbuf_top_iw_I[0].z ),
    .X(um_iw[162]));
 sky130_fd_sc_hd__buf_2 _0766_ (.A(\col[4].zbuf_top_iw_I[1].z ),
    .X(um_iw[163]));
 sky130_fd_sc_hd__buf_2 _0767_ (.A(\col[4].zbuf_top_iw_I[2].z ),
    .X(um_iw[164]));
 sky130_fd_sc_hd__buf_2 _0768_ (.A(\col[4].zbuf_top_iw_I[3].z ),
    .X(um_iw[165]));
 sky130_fd_sc_hd__buf_2 _0769_ (.A(\col[4].zbuf_top_iw_I[4].z ),
    .X(um_iw[166]));
 sky130_fd_sc_hd__buf_2 _0770_ (.A(\col[4].zbuf_top_iw_I[5].z ),
    .X(um_iw[167]));
 sky130_fd_sc_hd__buf_2 _0771_ (.A(\col[4].zbuf_top_iw_I[6].z ),
    .X(um_iw[168]));
 sky130_fd_sc_hd__buf_2 _0772_ (.A(\col[4].zbuf_top_iw_I[7].z ),
    .X(um_iw[169]));
 sky130_fd_sc_hd__buf_2 _0773_ (.A(\col[4].zbuf_top_iw_I[8].z ),
    .X(um_iw[170]));
 sky130_fd_sc_hd__buf_2 _0774_ (.A(\col[4].zbuf_top_iw_I[9].z ),
    .X(um_iw[171]));
 sky130_fd_sc_hd__buf_2 _0775_ (.A(\col[4].zbuf_top_iw_I[10].z ),
    .X(um_iw[172]));
 sky130_fd_sc_hd__buf_2 _0776_ (.A(\col[4].zbuf_top_iw_I[11].z ),
    .X(um_iw[173]));
 sky130_fd_sc_hd__buf_2 _0777_ (.A(\col[4].zbuf_top_iw_I[12].z ),
    .X(um_iw[174]));
 sky130_fd_sc_hd__buf_2 _0778_ (.A(\col[4].zbuf_top_iw_I[13].z ),
    .X(um_iw[175]));
 sky130_fd_sc_hd__buf_2 _0779_ (.A(\col[4].zbuf_top_iw_I[14].z ),
    .X(um_iw[176]));
 sky130_fd_sc_hd__buf_2 _0780_ (.A(\col[4].zbuf_top_iw_I[15].z ),
    .X(um_iw[177]));
 sky130_fd_sc_hd__buf_2 _0781_ (.A(\col[4].zbuf_top_iw_I[16].z ),
    .X(um_iw[178]));
 sky130_fd_sc_hd__buf_2 _0782_ (.A(\col[4].zbuf_top_iw_I[17].z ),
    .X(um_iw[179]));
 sky130_fd_sc_hd__buf_2 _0783_ (.A(\col[5].zbuf_bot_iw_I[0].z ),
    .X(um_iw[180]));
 sky130_fd_sc_hd__buf_2 _0784_ (.A(\col[5].zbuf_bot_iw_I[1].z ),
    .X(um_iw[181]));
 sky130_fd_sc_hd__buf_2 _0785_ (.A(\col[5].zbuf_bot_iw_I[2].z ),
    .X(um_iw[182]));
 sky130_fd_sc_hd__buf_2 _0786_ (.A(\col[5].zbuf_bot_iw_I[3].z ),
    .X(um_iw[183]));
 sky130_fd_sc_hd__buf_2 _0787_ (.A(\col[5].zbuf_bot_iw_I[4].z ),
    .X(um_iw[184]));
 sky130_fd_sc_hd__buf_2 _0788_ (.A(\col[5].zbuf_bot_iw_I[5].z ),
    .X(um_iw[185]));
 sky130_fd_sc_hd__buf_2 _0789_ (.A(\col[5].zbuf_bot_iw_I[6].z ),
    .X(um_iw[186]));
 sky130_fd_sc_hd__buf_2 _0790_ (.A(\col[5].zbuf_bot_iw_I[7].z ),
    .X(um_iw[187]));
 sky130_fd_sc_hd__buf_2 _0791_ (.A(\col[5].zbuf_bot_iw_I[8].z ),
    .X(um_iw[188]));
 sky130_fd_sc_hd__buf_2 _0792_ (.A(\col[5].zbuf_bot_iw_I[9].z ),
    .X(um_iw[189]));
 sky130_fd_sc_hd__buf_2 _0793_ (.A(\col[5].zbuf_bot_iw_I[10].z ),
    .X(um_iw[190]));
 sky130_fd_sc_hd__buf_2 _0794_ (.A(\col[5].zbuf_bot_iw_I[11].z ),
    .X(um_iw[191]));
 sky130_fd_sc_hd__buf_2 _0795_ (.A(\col[5].zbuf_bot_iw_I[12].z ),
    .X(um_iw[192]));
 sky130_fd_sc_hd__buf_2 _0796_ (.A(\col[5].zbuf_bot_iw_I[13].z ),
    .X(um_iw[193]));
 sky130_fd_sc_hd__buf_2 _0797_ (.A(\col[5].zbuf_bot_iw_I[14].z ),
    .X(um_iw[194]));
 sky130_fd_sc_hd__buf_2 _0798_ (.A(\col[5].zbuf_bot_iw_I[15].z ),
    .X(um_iw[195]));
 sky130_fd_sc_hd__buf_2 _0799_ (.A(\col[5].zbuf_bot_iw_I[16].z ),
    .X(um_iw[196]));
 sky130_fd_sc_hd__buf_2 _0800_ (.A(\col[5].zbuf_bot_iw_I[17].z ),
    .X(um_iw[197]));
 sky130_fd_sc_hd__buf_2 _0801_ (.A(\col[5].zbuf_top_iw_I[0].z ),
    .X(um_iw[198]));
 sky130_fd_sc_hd__buf_2 _0802_ (.A(\col[5].zbuf_top_iw_I[1].z ),
    .X(um_iw[199]));
 sky130_fd_sc_hd__buf_2 _0803_ (.A(\col[5].zbuf_top_iw_I[2].z ),
    .X(um_iw[200]));
 sky130_fd_sc_hd__buf_2 _0804_ (.A(\col[5].zbuf_top_iw_I[3].z ),
    .X(um_iw[201]));
 sky130_fd_sc_hd__buf_2 _0805_ (.A(\col[5].zbuf_top_iw_I[4].z ),
    .X(um_iw[202]));
 sky130_fd_sc_hd__buf_2 _0806_ (.A(\col[5].zbuf_top_iw_I[5].z ),
    .X(um_iw[203]));
 sky130_fd_sc_hd__buf_2 _0807_ (.A(\col[5].zbuf_top_iw_I[6].z ),
    .X(um_iw[204]));
 sky130_fd_sc_hd__buf_2 _0808_ (.A(\col[5].zbuf_top_iw_I[7].z ),
    .X(um_iw[205]));
 sky130_fd_sc_hd__buf_2 _0809_ (.A(\col[5].zbuf_top_iw_I[8].z ),
    .X(um_iw[206]));
 sky130_fd_sc_hd__buf_2 _0810_ (.A(\col[5].zbuf_top_iw_I[9].z ),
    .X(um_iw[207]));
 sky130_fd_sc_hd__buf_2 _0811_ (.A(\col[5].zbuf_top_iw_I[10].z ),
    .X(um_iw[208]));
 sky130_fd_sc_hd__buf_2 _0812_ (.A(\col[5].zbuf_top_iw_I[11].z ),
    .X(um_iw[209]));
 sky130_fd_sc_hd__buf_2 _0813_ (.A(\col[5].zbuf_top_iw_I[12].z ),
    .X(um_iw[210]));
 sky130_fd_sc_hd__buf_2 _0814_ (.A(\col[5].zbuf_top_iw_I[13].z ),
    .X(um_iw[211]));
 sky130_fd_sc_hd__buf_2 _0815_ (.A(\col[5].zbuf_top_iw_I[14].z ),
    .X(um_iw[212]));
 sky130_fd_sc_hd__buf_2 _0816_ (.A(\col[5].zbuf_top_iw_I[15].z ),
    .X(um_iw[213]));
 sky130_fd_sc_hd__buf_2 _0817_ (.A(\col[5].zbuf_top_iw_I[16].z ),
    .X(um_iw[214]));
 sky130_fd_sc_hd__buf_2 _0818_ (.A(\col[5].zbuf_top_iw_I[17].z ),
    .X(um_iw[215]));
 sky130_fd_sc_hd__buf_2 _0819_ (.A(\col[6].zbuf_bot_iw_I[0].z ),
    .X(um_iw[216]));
 sky130_fd_sc_hd__buf_2 _0820_ (.A(\col[6].zbuf_bot_iw_I[1].z ),
    .X(um_iw[217]));
 sky130_fd_sc_hd__buf_2 _0821_ (.A(\col[6].zbuf_bot_iw_I[2].z ),
    .X(um_iw[218]));
 sky130_fd_sc_hd__buf_2 _0822_ (.A(\col[6].zbuf_bot_iw_I[3].z ),
    .X(um_iw[219]));
 sky130_fd_sc_hd__buf_2 _0823_ (.A(\col[6].zbuf_bot_iw_I[4].z ),
    .X(um_iw[220]));
 sky130_fd_sc_hd__buf_2 _0824_ (.A(\col[6].zbuf_bot_iw_I[5].z ),
    .X(um_iw[221]));
 sky130_fd_sc_hd__buf_2 _0825_ (.A(\col[6].zbuf_bot_iw_I[6].z ),
    .X(um_iw[222]));
 sky130_fd_sc_hd__buf_2 _0826_ (.A(\col[6].zbuf_bot_iw_I[7].z ),
    .X(um_iw[223]));
 sky130_fd_sc_hd__buf_2 _0827_ (.A(\col[6].zbuf_bot_iw_I[8].z ),
    .X(um_iw[224]));
 sky130_fd_sc_hd__buf_2 _0828_ (.A(\col[6].zbuf_bot_iw_I[9].z ),
    .X(um_iw[225]));
 sky130_fd_sc_hd__buf_2 _0829_ (.A(\col[6].zbuf_bot_iw_I[10].z ),
    .X(um_iw[226]));
 sky130_fd_sc_hd__buf_2 _0830_ (.A(\col[6].zbuf_bot_iw_I[11].z ),
    .X(um_iw[227]));
 sky130_fd_sc_hd__buf_2 _0831_ (.A(\col[6].zbuf_bot_iw_I[12].z ),
    .X(um_iw[228]));
 sky130_fd_sc_hd__buf_2 _0832_ (.A(\col[6].zbuf_bot_iw_I[13].z ),
    .X(um_iw[229]));
 sky130_fd_sc_hd__buf_2 _0833_ (.A(\col[6].zbuf_bot_iw_I[14].z ),
    .X(um_iw[230]));
 sky130_fd_sc_hd__buf_2 _0834_ (.A(\col[6].zbuf_bot_iw_I[15].z ),
    .X(um_iw[231]));
 sky130_fd_sc_hd__buf_2 _0835_ (.A(\col[6].zbuf_bot_iw_I[16].z ),
    .X(um_iw[232]));
 sky130_fd_sc_hd__buf_2 _0836_ (.A(\col[6].zbuf_bot_iw_I[17].z ),
    .X(um_iw[233]));
 sky130_fd_sc_hd__buf_2 _0837_ (.A(\col[6].zbuf_top_iw_I[0].z ),
    .X(um_iw[234]));
 sky130_fd_sc_hd__buf_2 _0838_ (.A(\col[6].zbuf_top_iw_I[1].z ),
    .X(um_iw[235]));
 sky130_fd_sc_hd__buf_2 _0839_ (.A(\col[6].zbuf_top_iw_I[2].z ),
    .X(um_iw[236]));
 sky130_fd_sc_hd__buf_2 _0840_ (.A(\col[6].zbuf_top_iw_I[3].z ),
    .X(um_iw[237]));
 sky130_fd_sc_hd__buf_2 _0841_ (.A(\col[6].zbuf_top_iw_I[4].z ),
    .X(um_iw[238]));
 sky130_fd_sc_hd__buf_2 _0842_ (.A(\col[6].zbuf_top_iw_I[5].z ),
    .X(um_iw[239]));
 sky130_fd_sc_hd__buf_2 _0843_ (.A(\col[6].zbuf_top_iw_I[6].z ),
    .X(um_iw[240]));
 sky130_fd_sc_hd__buf_2 _0844_ (.A(\col[6].zbuf_top_iw_I[7].z ),
    .X(um_iw[241]));
 sky130_fd_sc_hd__buf_2 _0845_ (.A(\col[6].zbuf_top_iw_I[8].z ),
    .X(um_iw[242]));
 sky130_fd_sc_hd__buf_2 _0846_ (.A(\col[6].zbuf_top_iw_I[9].z ),
    .X(um_iw[243]));
 sky130_fd_sc_hd__buf_2 _0847_ (.A(\col[6].zbuf_top_iw_I[10].z ),
    .X(um_iw[244]));
 sky130_fd_sc_hd__buf_2 _0848_ (.A(\col[6].zbuf_top_iw_I[11].z ),
    .X(um_iw[245]));
 sky130_fd_sc_hd__buf_2 _0849_ (.A(\col[6].zbuf_top_iw_I[12].z ),
    .X(um_iw[246]));
 sky130_fd_sc_hd__buf_2 _0850_ (.A(\col[6].zbuf_top_iw_I[13].z ),
    .X(um_iw[247]));
 sky130_fd_sc_hd__buf_2 _0851_ (.A(\col[6].zbuf_top_iw_I[14].z ),
    .X(um_iw[248]));
 sky130_fd_sc_hd__buf_2 _0852_ (.A(\col[6].zbuf_top_iw_I[15].z ),
    .X(um_iw[249]));
 sky130_fd_sc_hd__buf_2 _0853_ (.A(\col[6].zbuf_top_iw_I[16].z ),
    .X(um_iw[250]));
 sky130_fd_sc_hd__buf_2 _0854_ (.A(\col[6].zbuf_top_iw_I[17].z ),
    .X(um_iw[251]));
 sky130_fd_sc_hd__buf_2 _0855_ (.A(\col[7].zbuf_bot_iw_I[0].z ),
    .X(um_iw[252]));
 sky130_fd_sc_hd__buf_2 _0856_ (.A(\col[7].zbuf_bot_iw_I[1].z ),
    .X(um_iw[253]));
 sky130_fd_sc_hd__buf_2 _0857_ (.A(\col[7].zbuf_bot_iw_I[2].z ),
    .X(um_iw[254]));
 sky130_fd_sc_hd__buf_2 _0858_ (.A(\col[7].zbuf_bot_iw_I[3].z ),
    .X(um_iw[255]));
 sky130_fd_sc_hd__buf_2 _0859_ (.A(\col[7].zbuf_bot_iw_I[4].z ),
    .X(um_iw[256]));
 sky130_fd_sc_hd__buf_2 _0860_ (.A(\col[7].zbuf_bot_iw_I[5].z ),
    .X(um_iw[257]));
 sky130_fd_sc_hd__buf_2 _0861_ (.A(\col[7].zbuf_bot_iw_I[6].z ),
    .X(um_iw[258]));
 sky130_fd_sc_hd__buf_2 _0862_ (.A(\col[7].zbuf_bot_iw_I[7].z ),
    .X(um_iw[259]));
 sky130_fd_sc_hd__buf_2 _0863_ (.A(\col[7].zbuf_bot_iw_I[8].z ),
    .X(um_iw[260]));
 sky130_fd_sc_hd__buf_2 _0864_ (.A(\col[7].zbuf_bot_iw_I[9].z ),
    .X(um_iw[261]));
 sky130_fd_sc_hd__buf_2 _0865_ (.A(\col[7].zbuf_bot_iw_I[10].z ),
    .X(um_iw[262]));
 sky130_fd_sc_hd__buf_2 _0866_ (.A(\col[7].zbuf_bot_iw_I[11].z ),
    .X(um_iw[263]));
 sky130_fd_sc_hd__buf_2 _0867_ (.A(\col[7].zbuf_bot_iw_I[12].z ),
    .X(um_iw[264]));
 sky130_fd_sc_hd__buf_2 _0868_ (.A(\col[7].zbuf_bot_iw_I[13].z ),
    .X(um_iw[265]));
 sky130_fd_sc_hd__buf_2 _0869_ (.A(\col[7].zbuf_bot_iw_I[14].z ),
    .X(um_iw[266]));
 sky130_fd_sc_hd__buf_2 _0870_ (.A(\col[7].zbuf_bot_iw_I[15].z ),
    .X(um_iw[267]));
 sky130_fd_sc_hd__buf_2 _0871_ (.A(\col[7].zbuf_bot_iw_I[16].z ),
    .X(um_iw[268]));
 sky130_fd_sc_hd__buf_2 _0872_ (.A(\col[7].zbuf_bot_iw_I[17].z ),
    .X(um_iw[269]));
 sky130_fd_sc_hd__buf_2 _0873_ (.A(\col[7].zbuf_top_iw_I[0].z ),
    .X(um_iw[270]));
 sky130_fd_sc_hd__buf_2 _0874_ (.A(\col[7].zbuf_top_iw_I[1].z ),
    .X(um_iw[271]));
 sky130_fd_sc_hd__buf_2 _0875_ (.A(\col[7].zbuf_top_iw_I[2].z ),
    .X(um_iw[272]));
 sky130_fd_sc_hd__buf_2 _0876_ (.A(\col[7].zbuf_top_iw_I[3].z ),
    .X(um_iw[273]));
 sky130_fd_sc_hd__buf_2 _0877_ (.A(\col[7].zbuf_top_iw_I[4].z ),
    .X(um_iw[274]));
 sky130_fd_sc_hd__buf_2 _0878_ (.A(\col[7].zbuf_top_iw_I[5].z ),
    .X(um_iw[275]));
 sky130_fd_sc_hd__buf_2 _0879_ (.A(\col[7].zbuf_top_iw_I[6].z ),
    .X(um_iw[276]));
 sky130_fd_sc_hd__buf_2 _0880_ (.A(\col[7].zbuf_top_iw_I[7].z ),
    .X(um_iw[277]));
 sky130_fd_sc_hd__buf_2 _0881_ (.A(\col[7].zbuf_top_iw_I[8].z ),
    .X(um_iw[278]));
 sky130_fd_sc_hd__buf_2 _0882_ (.A(\col[7].zbuf_top_iw_I[9].z ),
    .X(um_iw[279]));
 sky130_fd_sc_hd__buf_2 _0883_ (.A(\col[7].zbuf_top_iw_I[10].z ),
    .X(um_iw[280]));
 sky130_fd_sc_hd__buf_2 _0884_ (.A(\col[7].zbuf_top_iw_I[11].z ),
    .X(um_iw[281]));
 sky130_fd_sc_hd__buf_2 _0885_ (.A(\col[7].zbuf_top_iw_I[12].z ),
    .X(um_iw[282]));
 sky130_fd_sc_hd__buf_2 _0886_ (.A(\col[7].zbuf_top_iw_I[13].z ),
    .X(um_iw[283]));
 sky130_fd_sc_hd__buf_2 _0887_ (.A(\col[7].zbuf_top_iw_I[14].z ),
    .X(um_iw[284]));
 sky130_fd_sc_hd__buf_2 _0888_ (.A(\col[7].zbuf_top_iw_I[15].z ),
    .X(um_iw[285]));
 sky130_fd_sc_hd__buf_2 _0889_ (.A(\col[7].zbuf_top_iw_I[16].z ),
    .X(um_iw[286]));
 sky130_fd_sc_hd__buf_2 _0890_ (.A(\col[7].zbuf_top_iw_I[17].z ),
    .X(um_iw[287]));
 sky130_fd_sc_hd__buf_2 _0891_ (.A(\col[0].zbuf_bot_ena_I.z ),
    .X(um_ena[0]));
 sky130_fd_sc_hd__buf_2 _0892_ (.A(\col[0].zbuf_top_ena_I.z ),
    .X(um_ena[1]));
 sky130_fd_sc_hd__buf_2 _0893_ (.A(\col[1].zbuf_bot_ena_I.z ),
    .X(um_ena[2]));
 sky130_fd_sc_hd__buf_2 _0894_ (.A(\col[1].zbuf_top_ena_I.z ),
    .X(um_ena[3]));
 sky130_fd_sc_hd__buf_2 _0895_ (.A(\col[2].zbuf_bot_ena_I.z ),
    .X(um_ena[4]));
 sky130_fd_sc_hd__buf_2 _0896_ (.A(\col[2].zbuf_top_ena_I.z ),
    .X(um_ena[5]));
 sky130_fd_sc_hd__buf_2 _0897_ (.A(\col[3].zbuf_bot_ena_I.z ),
    .X(um_ena[6]));
 sky130_fd_sc_hd__buf_2 _0898_ (.A(\col[3].zbuf_top_ena_I.z ),
    .X(um_ena[7]));
 sky130_fd_sc_hd__buf_2 _0899_ (.A(\col[4].zbuf_bot_ena_I.z ),
    .X(um_ena[8]));
 sky130_fd_sc_hd__buf_2 _0900_ (.A(\col[4].zbuf_top_ena_I.z ),
    .X(um_ena[9]));
 sky130_fd_sc_hd__buf_2 _0901_ (.A(\col[5].zbuf_bot_ena_I.z ),
    .X(um_ena[10]));
 sky130_fd_sc_hd__buf_2 _0902_ (.A(\col[5].zbuf_top_ena_I.z ),
    .X(um_ena[11]));
 sky130_fd_sc_hd__buf_2 _0903_ (.A(\col[6].zbuf_bot_ena_I.z ),
    .X(um_ena[12]));
 sky130_fd_sc_hd__buf_2 _0904_ (.A(\col[6].zbuf_top_ena_I.z ),
    .X(um_ena[13]));
 sky130_fd_sc_hd__buf_2 _0905_ (.A(\col[7].zbuf_bot_ena_I.z ),
    .X(um_ena[14]));
 sky130_fd_sc_hd__buf_2 _0906_ (.A(\col[7].zbuf_top_ena_I.z ),
    .X(um_ena[15]));
 sky130_fd_sc_hd__buf_2 _0907_ (.A(\col[0].zbuf_bot_iw_I[0].z ),
    .X(um_iw[0]));
 sky130_fd_sc_hd__buf_2 _0908_ (.A(\col[0].zbuf_bot_iw_I[1].z ),
    .X(um_iw[1]));
 sky130_fd_sc_hd__buf_2 _0909_ (.A(\col[0].zbuf_bot_iw_I[2].z ),
    .X(um_iw[2]));
 sky130_fd_sc_hd__buf_2 _0910_ (.A(\col[0].zbuf_bot_iw_I[3].z ),
    .X(um_iw[3]));
 sky130_fd_sc_hd__buf_2 _0911_ (.A(\col[0].zbuf_bot_iw_I[4].z ),
    .X(um_iw[4]));
 sky130_fd_sc_hd__buf_2 _0912_ (.A(\col[0].zbuf_bot_iw_I[5].z ),
    .X(um_iw[5]));
 sky130_fd_sc_hd__buf_2 _0913_ (.A(\col[0].zbuf_bot_iw_I[6].z ),
    .X(um_iw[6]));
 sky130_fd_sc_hd__buf_2 _0914_ (.A(\col[0].zbuf_bot_iw_I[7].z ),
    .X(um_iw[7]));
 sky130_fd_sc_hd__buf_2 _0915_ (.A(\col[0].zbuf_bot_iw_I[8].z ),
    .X(um_iw[8]));
 sky130_fd_sc_hd__buf_2 _0916_ (.A(\col[0].zbuf_bot_iw_I[9].z ),
    .X(um_iw[9]));
 sky130_fd_sc_hd__buf_2 _0917_ (.A(\col[0].zbuf_bot_iw_I[10].z ),
    .X(um_iw[10]));
 sky130_fd_sc_hd__buf_2 _0918_ (.A(\col[0].zbuf_bot_iw_I[11].z ),
    .X(um_iw[11]));
 sky130_fd_sc_hd__buf_2 _0919_ (.A(\col[0].zbuf_bot_iw_I[12].z ),
    .X(um_iw[12]));
 sky130_fd_sc_hd__buf_2 _0920_ (.A(\col[0].zbuf_bot_iw_I[13].z ),
    .X(um_iw[13]));
 sky130_fd_sc_hd__buf_2 _0921_ (.A(\col[0].zbuf_bot_iw_I[14].z ),
    .X(um_iw[14]));
 sky130_fd_sc_hd__clkbuf_4 _0922_ (.A(\col[0].zbuf_bot_iw_I[15].z ),
    .X(um_iw[15]));
 sky130_fd_sc_hd__clkbuf_4 _0923_ (.A(\col[0].zbuf_bot_iw_I[16].z ),
    .X(um_iw[16]));
 sky130_fd_sc_hd__clkbuf_4 _0924_ (.A(\col[0].zbuf_bot_iw_I[17].z ),
    .X(um_iw[17]));
 sky130_fd_sc_hd__buf_2 _0925_ (.A(\col[0].zbuf_top_iw_I[0].z ),
    .X(um_iw[18]));
 sky130_fd_sc_hd__buf_2 _0926_ (.A(\col[0].zbuf_top_iw_I[1].z ),
    .X(um_iw[19]));
 sky130_fd_sc_hd__buf_2 _0927_ (.A(\col[0].zbuf_top_iw_I[2].z ),
    .X(um_iw[20]));
 sky130_fd_sc_hd__buf_2 _0928_ (.A(\col[0].zbuf_top_iw_I[3].z ),
    .X(um_iw[21]));
 sky130_fd_sc_hd__buf_2 _0929_ (.A(\col[0].zbuf_top_iw_I[4].z ),
    .X(um_iw[22]));
 sky130_fd_sc_hd__buf_2 _0930_ (.A(\col[0].zbuf_top_iw_I[5].z ),
    .X(um_iw[23]));
 sky130_fd_sc_hd__buf_2 _0931_ (.A(\col[0].zbuf_top_iw_I[6].z ),
    .X(um_iw[24]));
 sky130_fd_sc_hd__buf_2 _0932_ (.A(\col[0].zbuf_top_iw_I[7].z ),
    .X(um_iw[25]));
 sky130_fd_sc_hd__buf_2 _0933_ (.A(\col[0].zbuf_top_iw_I[8].z ),
    .X(um_iw[26]));
 sky130_fd_sc_hd__buf_2 _0934_ (.A(\col[0].zbuf_top_iw_I[9].z ),
    .X(um_iw[27]));
 sky130_fd_sc_hd__buf_2 _0935_ (.A(\col[0].zbuf_top_iw_I[10].z ),
    .X(um_iw[28]));
 sky130_fd_sc_hd__buf_2 _0936_ (.A(\col[0].zbuf_top_iw_I[11].z ),
    .X(um_iw[29]));
 sky130_fd_sc_hd__buf_2 _0937_ (.A(\col[0].zbuf_top_iw_I[12].z ),
    .X(um_iw[30]));
 sky130_fd_sc_hd__buf_2 _0938_ (.A(\col[0].zbuf_top_iw_I[13].z ),
    .X(um_iw[31]));
 sky130_fd_sc_hd__buf_2 _0939_ (.A(\col[0].zbuf_top_iw_I[14].z ),
    .X(um_iw[32]));
 sky130_fd_sc_hd__buf_2 _0940_ (.A(\col[0].zbuf_top_iw_I[15].z ),
    .X(um_iw[33]));
 sky130_fd_sc_hd__clkbuf_4 _0941_ (.A(\col[0].zbuf_top_iw_I[16].z ),
    .X(um_iw[34]));
 sky130_fd_sc_hd__clkbuf_4 _0942_ (.A(\col[0].zbuf_top_iw_I[17].z ),
    .X(um_iw[35]));
 sky130_fd_sc_hd__buf_2 _0943_ (.A(\col[1].zbuf_bot_iw_I[0].z ),
    .X(um_iw[36]));
 sky130_fd_sc_hd__buf_2 _0944_ (.A(\col[1].zbuf_bot_iw_I[1].z ),
    .X(um_iw[37]));
 sky130_fd_sc_hd__buf_2 _0945_ (.A(\col[1].zbuf_bot_iw_I[2].z ),
    .X(um_iw[38]));
 sky130_fd_sc_hd__buf_2 _0946_ (.A(\col[1].zbuf_bot_iw_I[3].z ),
    .X(um_iw[39]));
 sky130_fd_sc_hd__ebufn_8 _0947_ (.A(\bus_ow[0] ),
    .TE_B(_0167_),
    .Z(spine_ow[1]));
 sky130_fd_sc_hd__ebufn_8 _0948_ (.A(\bus_ow[1] ),
    .TE_B(_0168_),
    .Z(spine_ow[2]));
 sky130_fd_sc_hd__ebufn_8 _0949_ (.A(\bus_ow[2] ),
    .TE_B(_0169_),
    .Z(spine_ow[3]));
 sky130_fd_sc_hd__ebufn_8 _0950_ (.A(\bus_ow[3] ),
    .TE_B(_0170_),
    .Z(spine_ow[4]));
 sky130_fd_sc_hd__ebufn_8 _0951_ (.A(\bus_ow[4] ),
    .TE_B(_0171_),
    .Z(spine_ow[5]));
 sky130_fd_sc_hd__ebufn_8 _0952_ (.A(\bus_ow[5] ),
    .TE_B(_0172_),
    .Z(spine_ow[6]));
 sky130_fd_sc_hd__ebufn_8 _0953_ (.A(\bus_ow[6] ),
    .TE_B(_0173_),
    .Z(spine_ow[7]));
 sky130_fd_sc_hd__ebufn_8 _0954_ (.A(\bus_ow[7] ),
    .TE_B(_0174_),
    .Z(spine_ow[8]));
 sky130_fd_sc_hd__ebufn_8 _0955_ (.A(\bus_ow[8] ),
    .TE_B(_0175_),
    .Z(spine_ow[9]));
 sky130_fd_sc_hd__ebufn_8 _0956_ (.A(\bus_ow[9] ),
    .TE_B(_0176_),
    .Z(spine_ow[10]));
 sky130_fd_sc_hd__ebufn_8 _0957_ (.A(\bus_ow[10] ),
    .TE_B(_0177_),
    .Z(spine_ow[11]));
 sky130_fd_sc_hd__ebufn_8 _0958_ (.A(\bus_ow[11] ),
    .TE_B(_0178_),
    .Z(spine_ow[12]));
 sky130_fd_sc_hd__ebufn_8 _0959_ (.A(\bus_ow[12] ),
    .TE_B(_0179_),
    .Z(spine_ow[13]));
 sky130_fd_sc_hd__ebufn_8 _0960_ (.A(\bus_ow[13] ),
    .TE_B(_0180_),
    .Z(spine_ow[14]));
 sky130_fd_sc_hd__ebufn_8 _0961_ (.A(\bus_ow[14] ),
    .TE_B(_0181_),
    .Z(spine_ow[15]));
 sky130_fd_sc_hd__ebufn_8 _0962_ (.A(\bus_ow[15] ),
    .TE_B(_0182_),
    .Z(spine_ow[16]));
 sky130_fd_sc_hd__ebufn_8 _0963_ (.A(\bus_ow[16] ),
    .TE_B(_0183_),
    .Z(spine_ow[17]));
 sky130_fd_sc_hd__ebufn_8 _0964_ (.A(\bus_ow[17] ),
    .TE_B(_0184_),
    .Z(spine_ow[18]));
 sky130_fd_sc_hd__ebufn_8 _0965_ (.A(\bus_ow[18] ),
    .TE_B(_0185_),
    .Z(spine_ow[19]));
 sky130_fd_sc_hd__ebufn_8 _0966_ (.A(\bus_ow[19] ),
    .TE_B(_0186_),
    .Z(spine_ow[20]));
 sky130_fd_sc_hd__ebufn_8 _0967_ (.A(\bus_ow[20] ),
    .TE_B(_0187_),
    .Z(spine_ow[21]));
 sky130_fd_sc_hd__ebufn_8 _0968_ (.A(\bus_ow[21] ),
    .TE_B(_0188_),
    .Z(spine_ow[22]));
 sky130_fd_sc_hd__ebufn_8 _0969_ (.A(\bus_ow[22] ),
    .TE_B(_0189_),
    .Z(spine_ow[23]));
 sky130_fd_sc_hd__ebufn_8 _0970_ (.A(\bus_ow[23] ),
    .TE_B(_0190_),
    .Z(spine_ow[24]));
 sky130_fd_sc_hd__ebufn_8 _0971_ (.A(\col[0].genblk1.mux4_I[0].x ),
    .TE_B(_0191_),
    .Z(\bus_ow[0] ));
 sky130_fd_sc_hd__ebufn_8 _0972_ (.A(\col[0].genblk1.mux4_I[1].x ),
    .TE_B(_0192_),
    .Z(\bus_ow[1] ));
 sky130_fd_sc_hd__ebufn_8 _0973_ (.A(\col[0].genblk1.mux4_I[2].x ),
    .TE_B(_0193_),
    .Z(\bus_ow[2] ));
 sky130_fd_sc_hd__ebufn_8 _0974_ (.A(\col[0].genblk1.mux4_I[3].x ),
    .TE_B(_0194_),
    .Z(\bus_ow[3] ));
 sky130_fd_sc_hd__ebufn_8 _0975_ (.A(\col[0].genblk1.mux4_I[4].x ),
    .TE_B(_0195_),
    .Z(\bus_ow[4] ));
 sky130_fd_sc_hd__ebufn_8 _0976_ (.A(\col[0].genblk1.mux4_I[5].x ),
    .TE_B(_0196_),
    .Z(\bus_ow[5] ));
 sky130_fd_sc_hd__ebufn_8 _0977_ (.A(\col[0].genblk1.mux4_I[6].x ),
    .TE_B(_0197_),
    .Z(\bus_ow[6] ));
 sky130_fd_sc_hd__ebufn_8 _0978_ (.A(\col[0].genblk1.mux4_I[7].x ),
    .TE_B(_0198_),
    .Z(\bus_ow[7] ));
 sky130_fd_sc_hd__ebufn_8 _0979_ (.A(\col[0].genblk1.mux4_I[8].x ),
    .TE_B(_0199_),
    .Z(\bus_ow[8] ));
 sky130_fd_sc_hd__ebufn_8 _0980_ (.A(\col[0].genblk1.mux4_I[9].x ),
    .TE_B(_0200_),
    .Z(\bus_ow[9] ));
 sky130_fd_sc_hd__ebufn_8 _0981_ (.A(\col[0].genblk1.mux4_I[10].x ),
    .TE_B(_0201_),
    .Z(\bus_ow[10] ));
 sky130_fd_sc_hd__ebufn_8 _0982_ (.A(\col[0].genblk1.mux4_I[11].x ),
    .TE_B(_0202_),
    .Z(\bus_ow[11] ));
 sky130_fd_sc_hd__ebufn_8 _0983_ (.A(\col[0].genblk1.mux4_I[12].x ),
    .TE_B(_0203_),
    .Z(\bus_ow[12] ));
 sky130_fd_sc_hd__ebufn_8 _0984_ (.A(\col[0].genblk1.mux4_I[13].x ),
    .TE_B(_0204_),
    .Z(\bus_ow[13] ));
 sky130_fd_sc_hd__ebufn_8 _0985_ (.A(\col[0].genblk1.mux4_I[14].x ),
    .TE_B(_0205_),
    .Z(\bus_ow[14] ));
 sky130_fd_sc_hd__ebufn_8 _0986_ (.A(\col[0].genblk1.mux4_I[15].x ),
    .TE_B(_0206_),
    .Z(\bus_ow[15] ));
 sky130_fd_sc_hd__ebufn_8 _0987_ (.A(\col[0].genblk1.mux4_I[16].x ),
    .TE_B(_0207_),
    .Z(\bus_ow[16] ));
 sky130_fd_sc_hd__ebufn_8 _0988_ (.A(\col[0].genblk1.mux4_I[17].x ),
    .TE_B(_0208_),
    .Z(\bus_ow[17] ));
 sky130_fd_sc_hd__ebufn_8 _0989_ (.A(\col[0].genblk1.mux4_I[18].x ),
    .TE_B(_0209_),
    .Z(\bus_ow[18] ));
 sky130_fd_sc_hd__ebufn_8 _0990_ (.A(\col[0].genblk1.mux4_I[19].x ),
    .TE_B(_0210_),
    .Z(\bus_ow[19] ));
 sky130_fd_sc_hd__ebufn_8 _0991_ (.A(\col[0].genblk1.mux4_I[20].x ),
    .TE_B(_0211_),
    .Z(\bus_ow[20] ));
 sky130_fd_sc_hd__ebufn_8 _0992_ (.A(\col[0].genblk1.mux4_I[21].x ),
    .TE_B(_0212_),
    .Z(\bus_ow[21] ));
 sky130_fd_sc_hd__ebufn_8 _0993_ (.A(\col[0].genblk1.mux4_I[22].x ),
    .TE_B(_0213_),
    .Z(\bus_ow[22] ));
 sky130_fd_sc_hd__ebufn_8 _0994_ (.A(\col[0].genblk1.mux4_I[23].x ),
    .TE_B(_0214_),
    .Z(\bus_ow[23] ));
 sky130_fd_sc_hd__ebufn_8 _0995_ (.A(\col[2].genblk1.mux4_I[0].x ),
    .TE_B(_0215_),
    .Z(\bus_ow[0] ));
 sky130_fd_sc_hd__ebufn_8 _0996_ (.A(\col[2].genblk1.mux4_I[1].x ),
    .TE_B(_0216_),
    .Z(\bus_ow[1] ));
 sky130_fd_sc_hd__ebufn_8 _0997_ (.A(\col[2].genblk1.mux4_I[2].x ),
    .TE_B(_0217_),
    .Z(\bus_ow[2] ));
 sky130_fd_sc_hd__ebufn_8 _0998_ (.A(\col[2].genblk1.mux4_I[3].x ),
    .TE_B(_0218_),
    .Z(\bus_ow[3] ));
 sky130_fd_sc_hd__ebufn_8 _0999_ (.A(\col[2].genblk1.mux4_I[4].x ),
    .TE_B(_0219_),
    .Z(\bus_ow[4] ));
 sky130_fd_sc_hd__ebufn_8 _1000_ (.A(\col[2].genblk1.mux4_I[5].x ),
    .TE_B(_0220_),
    .Z(\bus_ow[5] ));
 sky130_fd_sc_hd__ebufn_8 _1001_ (.A(\col[2].genblk1.mux4_I[6].x ),
    .TE_B(_0221_),
    .Z(\bus_ow[6] ));
 sky130_fd_sc_hd__ebufn_8 _1002_ (.A(\col[2].genblk1.mux4_I[7].x ),
    .TE_B(_0222_),
    .Z(\bus_ow[7] ));
 sky130_fd_sc_hd__ebufn_8 _1003_ (.A(\col[2].genblk1.mux4_I[8].x ),
    .TE_B(_0223_),
    .Z(\bus_ow[8] ));
 sky130_fd_sc_hd__ebufn_8 _1004_ (.A(\col[2].genblk1.mux4_I[9].x ),
    .TE_B(_0224_),
    .Z(\bus_ow[9] ));
 sky130_fd_sc_hd__ebufn_8 _1005_ (.A(\col[2].genblk1.mux4_I[10].x ),
    .TE_B(_0225_),
    .Z(\bus_ow[10] ));
 sky130_fd_sc_hd__ebufn_8 _1006_ (.A(\col[2].genblk1.mux4_I[11].x ),
    .TE_B(_0226_),
    .Z(\bus_ow[11] ));
 sky130_fd_sc_hd__ebufn_8 _1007_ (.A(\col[2].genblk1.mux4_I[12].x ),
    .TE_B(_0227_),
    .Z(\bus_ow[12] ));
 sky130_fd_sc_hd__ebufn_8 _1008_ (.A(\col[2].genblk1.mux4_I[13].x ),
    .TE_B(_0228_),
    .Z(\bus_ow[13] ));
 sky130_fd_sc_hd__ebufn_8 _1009_ (.A(\col[2].genblk1.mux4_I[14].x ),
    .TE_B(_0229_),
    .Z(\bus_ow[14] ));
 sky130_fd_sc_hd__ebufn_8 _1010_ (.A(\col[2].genblk1.mux4_I[15].x ),
    .TE_B(_0230_),
    .Z(\bus_ow[15] ));
 sky130_fd_sc_hd__ebufn_8 _1011_ (.A(\col[2].genblk1.mux4_I[16].x ),
    .TE_B(_0231_),
    .Z(\bus_ow[16] ));
 sky130_fd_sc_hd__ebufn_8 _1012_ (.A(\col[2].genblk1.mux4_I[17].x ),
    .TE_B(_0232_),
    .Z(\bus_ow[17] ));
 sky130_fd_sc_hd__ebufn_8 _1013_ (.A(\col[2].genblk1.mux4_I[18].x ),
    .TE_B(_0233_),
    .Z(\bus_ow[18] ));
 sky130_fd_sc_hd__ebufn_8 _1014_ (.A(\col[2].genblk1.mux4_I[19].x ),
    .TE_B(_0234_),
    .Z(\bus_ow[19] ));
 sky130_fd_sc_hd__ebufn_8 _1015_ (.A(\col[2].genblk1.mux4_I[20].x ),
    .TE_B(_0235_),
    .Z(\bus_ow[20] ));
 sky130_fd_sc_hd__ebufn_8 _1016_ (.A(\col[2].genblk1.mux4_I[21].x ),
    .TE_B(_0236_),
    .Z(\bus_ow[21] ));
 sky130_fd_sc_hd__ebufn_8 _1017_ (.A(\col[2].genblk1.mux4_I[22].x ),
    .TE_B(_0237_),
    .Z(\bus_ow[22] ));
 sky130_fd_sc_hd__ebufn_8 _1018_ (.A(\col[2].genblk1.mux4_I[23].x ),
    .TE_B(_0238_),
    .Z(\bus_ow[23] ));
 sky130_fd_sc_hd__ebufn_8 _1019_ (.A(\col[4].genblk1.mux4_I[0].x ),
    .TE_B(_0239_),
    .Z(\bus_ow[0] ));
 sky130_fd_sc_hd__ebufn_8 _1020_ (.A(\col[4].genblk1.mux4_I[1].x ),
    .TE_B(_0240_),
    .Z(\bus_ow[1] ));
 sky130_fd_sc_hd__ebufn_8 _1021_ (.A(\col[4].genblk1.mux4_I[2].x ),
    .TE_B(_0241_),
    .Z(\bus_ow[2] ));
 sky130_fd_sc_hd__ebufn_8 _1022_ (.A(\col[4].genblk1.mux4_I[3].x ),
    .TE_B(_0242_),
    .Z(\bus_ow[3] ));
 sky130_fd_sc_hd__ebufn_8 _1023_ (.A(\col[4].genblk1.mux4_I[4].x ),
    .TE_B(_0243_),
    .Z(\bus_ow[4] ));
 sky130_fd_sc_hd__ebufn_8 _1024_ (.A(\col[4].genblk1.mux4_I[5].x ),
    .TE_B(_0244_),
    .Z(\bus_ow[5] ));
 sky130_fd_sc_hd__ebufn_8 _1025_ (.A(\col[4].genblk1.mux4_I[6].x ),
    .TE_B(_0245_),
    .Z(\bus_ow[6] ));
 sky130_fd_sc_hd__ebufn_8 _1026_ (.A(\col[4].genblk1.mux4_I[7].x ),
    .TE_B(_0246_),
    .Z(\bus_ow[7] ));
 sky130_fd_sc_hd__ebufn_8 _1027_ (.A(\col[4].genblk1.mux4_I[8].x ),
    .TE_B(_0247_),
    .Z(\bus_ow[8] ));
 sky130_fd_sc_hd__ebufn_8 _1028_ (.A(\col[4].genblk1.mux4_I[9].x ),
    .TE_B(_0248_),
    .Z(\bus_ow[9] ));
 sky130_fd_sc_hd__ebufn_8 _1029_ (.A(\col[4].genblk1.mux4_I[10].x ),
    .TE_B(_0249_),
    .Z(\bus_ow[10] ));
 sky130_fd_sc_hd__ebufn_8 _1030_ (.A(\col[4].genblk1.mux4_I[11].x ),
    .TE_B(_0250_),
    .Z(\bus_ow[11] ));
 sky130_fd_sc_hd__ebufn_8 _1031_ (.A(\col[4].genblk1.mux4_I[12].x ),
    .TE_B(_0251_),
    .Z(\bus_ow[12] ));
 sky130_fd_sc_hd__ebufn_8 _1032_ (.A(\col[4].genblk1.mux4_I[13].x ),
    .TE_B(_0252_),
    .Z(\bus_ow[13] ));
 sky130_fd_sc_hd__ebufn_8 _1033_ (.A(\col[4].genblk1.mux4_I[14].x ),
    .TE_B(_0253_),
    .Z(\bus_ow[14] ));
 sky130_fd_sc_hd__ebufn_8 _1034_ (.A(\col[4].genblk1.mux4_I[15].x ),
    .TE_B(_0254_),
    .Z(\bus_ow[15] ));
 sky130_fd_sc_hd__ebufn_8 _1035_ (.A(\col[4].genblk1.mux4_I[16].x ),
    .TE_B(_0255_),
    .Z(\bus_ow[16] ));
 sky130_fd_sc_hd__ebufn_8 _1036_ (.A(\col[4].genblk1.mux4_I[17].x ),
    .TE_B(_0256_),
    .Z(\bus_ow[17] ));
 sky130_fd_sc_hd__ebufn_8 _1037_ (.A(\col[4].genblk1.mux4_I[18].x ),
    .TE_B(_0257_),
    .Z(\bus_ow[18] ));
 sky130_fd_sc_hd__ebufn_8 _1038_ (.A(\col[4].genblk1.mux4_I[19].x ),
    .TE_B(_0258_),
    .Z(\bus_ow[19] ));
 sky130_fd_sc_hd__ebufn_8 _1039_ (.A(\col[4].genblk1.mux4_I[20].x ),
    .TE_B(_0259_),
    .Z(\bus_ow[20] ));
 sky130_fd_sc_hd__ebufn_8 _1040_ (.A(\col[4].genblk1.mux4_I[21].x ),
    .TE_B(_0260_),
    .Z(\bus_ow[21] ));
 sky130_fd_sc_hd__ebufn_8 _1041_ (.A(\col[4].genblk1.mux4_I[22].x ),
    .TE_B(_0261_),
    .Z(\bus_ow[22] ));
 sky130_fd_sc_hd__ebufn_8 _1042_ (.A(\col[4].genblk1.mux4_I[23].x ),
    .TE_B(_0262_),
    .Z(\bus_ow[23] ));
 sky130_fd_sc_hd__ebufn_8 _1043_ (.A(\col[6].genblk1.mux4_I[0].x ),
    .TE_B(_0263_),
    .Z(\bus_ow[0] ));
 sky130_fd_sc_hd__ebufn_8 _1044_ (.A(\col[6].genblk1.mux4_I[1].x ),
    .TE_B(_0264_),
    .Z(\bus_ow[1] ));
 sky130_fd_sc_hd__ebufn_8 _1045_ (.A(\col[6].genblk1.mux4_I[2].x ),
    .TE_B(_0265_),
    .Z(\bus_ow[2] ));
 sky130_fd_sc_hd__ebufn_8 _1046_ (.A(\col[6].genblk1.mux4_I[3].x ),
    .TE_B(_0266_),
    .Z(\bus_ow[3] ));
 sky130_fd_sc_hd__ebufn_8 _1047_ (.A(\col[6].genblk1.mux4_I[4].x ),
    .TE_B(_0267_),
    .Z(\bus_ow[4] ));
 sky130_fd_sc_hd__ebufn_8 _1048_ (.A(\col[6].genblk1.mux4_I[5].x ),
    .TE_B(_0268_),
    .Z(\bus_ow[5] ));
 sky130_fd_sc_hd__ebufn_8 _1049_ (.A(\col[6].genblk1.mux4_I[6].x ),
    .TE_B(_0269_),
    .Z(\bus_ow[6] ));
 sky130_fd_sc_hd__ebufn_8 _1050_ (.A(\col[6].genblk1.mux4_I[7].x ),
    .TE_B(_0270_),
    .Z(\bus_ow[7] ));
 sky130_fd_sc_hd__ebufn_8 _1051_ (.A(\col[6].genblk1.mux4_I[8].x ),
    .TE_B(_0271_),
    .Z(\bus_ow[8] ));
 sky130_fd_sc_hd__ebufn_8 _1052_ (.A(\col[6].genblk1.mux4_I[9].x ),
    .TE_B(_0272_),
    .Z(\bus_ow[9] ));
 sky130_fd_sc_hd__ebufn_8 _1053_ (.A(\col[6].genblk1.mux4_I[10].x ),
    .TE_B(_0273_),
    .Z(\bus_ow[10] ));
 sky130_fd_sc_hd__ebufn_8 _1054_ (.A(\col[6].genblk1.mux4_I[11].x ),
    .TE_B(_0274_),
    .Z(\bus_ow[11] ));
 sky130_fd_sc_hd__ebufn_8 _1055_ (.A(\col[6].genblk1.mux4_I[12].x ),
    .TE_B(_0275_),
    .Z(\bus_ow[12] ));
 sky130_fd_sc_hd__ebufn_8 _1056_ (.A(\col[6].genblk1.mux4_I[13].x ),
    .TE_B(_0276_),
    .Z(\bus_ow[13] ));
 sky130_fd_sc_hd__ebufn_8 _1057_ (.A(\col[6].genblk1.mux4_I[14].x ),
    .TE_B(_0277_),
    .Z(\bus_ow[14] ));
 sky130_fd_sc_hd__ebufn_8 _1058_ (.A(\col[6].genblk1.mux4_I[15].x ),
    .TE_B(_0278_),
    .Z(\bus_ow[15] ));
 sky130_fd_sc_hd__ebufn_8 _1059_ (.A(\col[6].genblk1.mux4_I[16].x ),
    .TE_B(_0279_),
    .Z(\bus_ow[16] ));
 sky130_fd_sc_hd__ebufn_8 _1060_ (.A(\col[6].genblk1.mux4_I[17].x ),
    .TE_B(_0280_),
    .Z(\bus_ow[17] ));
 sky130_fd_sc_hd__ebufn_8 _1061_ (.A(\col[6].genblk1.mux4_I[18].x ),
    .TE_B(_0281_),
    .Z(\bus_ow[18] ));
 sky130_fd_sc_hd__ebufn_8 _1062_ (.A(\col[6].genblk1.mux4_I[19].x ),
    .TE_B(_0282_),
    .Z(\bus_ow[19] ));
 sky130_fd_sc_hd__ebufn_8 _1063_ (.A(\col[6].genblk1.mux4_I[20].x ),
    .TE_B(_0283_),
    .Z(\bus_ow[20] ));
 sky130_fd_sc_hd__ebufn_8 _1064_ (.A(\col[6].genblk1.mux4_I[21].x ),
    .TE_B(_0284_),
    .Z(\bus_ow[21] ));
 sky130_fd_sc_hd__ebufn_8 _1065_ (.A(\col[6].genblk1.mux4_I[22].x ),
    .TE_B(_0285_),
    .Z(\bus_ow[22] ));
 sky130_fd_sc_hd__ebufn_8 _1066_ (.A(\col[6].genblk1.mux4_I[23].x ),
    .TE_B(_0286_),
    .Z(\bus_ow[23] ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[0].cell0_I  (.A0(net35),
    .A1(net201),
    .A2(net361),
    .A3(net388),
    .S0(net466),
    .S1(net453),
    .X(\col[0].genblk1.mux4_I[0].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[10].cell0_I  (.A0(net46),
    .A1(net312),
    .A2(net372),
    .A3(net399),
    .S0(net465),
    .S1(net452),
    .X(\col[0].genblk1.mux4_I[10].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[11].cell0_I  (.A0(net57),
    .A1(net323),
    .A2(net373),
    .A3(net400),
    .S0(net465),
    .S1(net452),
    .X(\col[0].genblk1.mux4_I[11].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[12].cell0_I  (.A0(net68),
    .A1(net334),
    .A2(net375),
    .A3(net401),
    .S0(net465),
    .S1(net452),
    .X(\col[0].genblk1.mux4_I[12].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[13].cell0_I  (.A0(net79),
    .A1(net345),
    .A2(net376),
    .A3(net402),
    .S0(net465),
    .S1(net452),
    .X(\col[0].genblk1.mux4_I[13].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[14].cell0_I  (.A0(net90),
    .A1(net350),
    .A2(net377),
    .A3(net403),
    .S0(net464),
    .S1(net451),
    .X(\col[0].genblk1.mux4_I[14].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[15].cell0_I  (.A0(net101),
    .A1(net351),
    .A2(net378),
    .A3(net404),
    .S0(net464),
    .S1(net451),
    .X(\col[0].genblk1.mux4_I[15].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[16].cell0_I  (.A0(net112),
    .A1(net353),
    .A2(net379),
    .A3(net405),
    .S0(net464),
    .S1(net451),
    .X(\col[0].genblk1.mux4_I[16].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[17].cell0_I  (.A0(net123),
    .A1(net354),
    .A2(net380),
    .A3(net406),
    .S0(net464),
    .S1(net451),
    .X(\col[0].genblk1.mux4_I[17].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[18].cell0_I  (.A0(net134),
    .A1(net355),
    .A2(net381),
    .A3(net408),
    .S0(net464),
    .S1(net451),
    .X(\col[0].genblk1.mux4_I[18].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[19].cell0_I  (.A0(net145),
    .A1(net356),
    .A2(net382),
    .A3(net409),
    .S0(net464),
    .S1(net451),
    .X(\col[0].genblk1.mux4_I[19].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[1].cell0_I  (.A0(net146),
    .A1(net212),
    .A2(net362),
    .A3(net389),
    .S0(net466),
    .S1(net453),
    .X(\col[0].genblk1.mux4_I[1].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[20].cell0_I  (.A0(net157),
    .A1(net357),
    .A2(net383),
    .A3(net410),
    .S0(net464),
    .S1(net451),
    .X(\col[0].genblk1.mux4_I[20].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[21].cell0_I  (.A0(net168),
    .A1(net358),
    .A2(net384),
    .A3(net411),
    .S0(net464),
    .S1(net451),
    .X(\col[0].genblk1.mux4_I[21].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[22].cell0_I  (.A0(net179),
    .A1(net359),
    .A2(net386),
    .A3(net412),
    .S0(net464),
    .S1(net451),
    .X(\col[0].genblk1.mux4_I[22].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[23].cell0_I  (.A0(net190),
    .A1(net360),
    .A2(net387),
    .A3(net413),
    .S0(net464),
    .S1(net451),
    .X(\col[0].genblk1.mux4_I[23].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[2].cell0_I  (.A0(net257),
    .A1(net223),
    .A2(net364),
    .A3(net390),
    .S0(net466),
    .S1(net453),
    .X(\col[0].genblk1.mux4_I[2].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[3].cell0_I  (.A0(net352),
    .A1(net234),
    .A2(net365),
    .A3(net391),
    .S0(net466),
    .S1(net453),
    .X(\col[0].genblk1.mux4_I[3].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[4].cell0_I  (.A0(net363),
    .A1(net245),
    .A2(net366),
    .A3(net392),
    .S0(net466),
    .S1(net453),
    .X(\col[0].genblk1.mux4_I[4].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[5].cell0_I  (.A0(net374),
    .A1(net256),
    .A2(net367),
    .A3(net393),
    .S0(net466),
    .S1(net453),
    .X(\col[0].genblk1.mux4_I[5].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[6].cell0_I  (.A0(net385),
    .A1(net268),
    .A2(net368),
    .A3(net394),
    .S0(net466),
    .S1(net452),
    .X(\col[0].genblk1.mux4_I[6].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[7].cell0_I  (.A0(net396),
    .A1(net279),
    .A2(net369),
    .A3(net395),
    .S0(net465),
    .S1(net452),
    .X(\col[0].genblk1.mux4_I[7].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[8].cell0_I  (.A0(net407),
    .A1(net290),
    .A2(net370),
    .A3(net397),
    .S0(net465),
    .S1(net452),
    .X(\col[0].genblk1.mux4_I[8].x ));
 sky130_fd_sc_hd__mux4_2 \col[0].genblk1.mux4_I[9].cell0_I  (.A0(net418),
    .A1(net301),
    .A2(net371),
    .A3(net398),
    .S0(net465),
    .S1(net452),
    .X(\col[0].genblk1.mux4_I[9].x ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_bot_ena_I.genblk1.cell0_I  (.A(net536),
    .B(net448),
    .X(\col[0].zbuf_bot_ena_I.z ));
 sky130_fd_sc_hd__conb_1 \col[0].zbuf_bot_ena_I.genblk1.cell0_I_536  (.HI(net536));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(net511),
    .B(net448),
    .X(\col[0].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(net509),
    .B(net447),
    .X(\col[0].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(net507),
    .B(net447),
    .X(\col[0].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(net505),
    .B(net447),
    .X(\col[0].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(net503),
    .B(net447),
    .X(\col[0].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(net501),
    .B(net447),
    .X(\col[0].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(net499),
    .B(net447),
    .X(\col[0].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(net497),
    .B(net447),
    .X(\col[0].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(net495),
    .B(net448),
    .X(\col[0].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(net493),
    .B(net448),
    .X(\col[0].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(net491),
    .B(net448),
    .X(\col[0].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(net489),
    .B(net448),
    .X(\col[0].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(net487),
    .B(net448),
    .X(\col[0].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(net485),
    .B(net448),
    .X(\col[0].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(net483),
    .B(net448),
    .X(\col[0].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(net481),
    .B(net447),
    .X(\col[0].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(net479),
    .B(net447),
    .X(\col[0].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(net477),
    .B(net447),
    .X(\col[0].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_top_ena_I.genblk1.cell0_I  (.A(net537),
    .B(net436),
    .X(\col[0].zbuf_top_ena_I.z ));
 sky130_fd_sc_hd__conb_1 \col[0].zbuf_top_ena_I.genblk1.cell0_I_537  (.HI(net537));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_top_iw_I[0].genblk1.cell0_I  (.A(net511),
    .B(net436),
    .X(\col[0].zbuf_top_iw_I[0].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_top_iw_I[10].genblk1.cell0_I  (.A(net509),
    .B(net435),
    .X(\col[0].zbuf_top_iw_I[10].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_top_iw_I[11].genblk1.cell0_I  (.A(net507),
    .B(net435),
    .X(\col[0].zbuf_top_iw_I[11].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_top_iw_I[12].genblk1.cell0_I  (.A(net505),
    .B(net435),
    .X(\col[0].zbuf_top_iw_I[12].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_top_iw_I[13].genblk1.cell0_I  (.A(net503),
    .B(net435),
    .X(\col[0].zbuf_top_iw_I[13].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_top_iw_I[14].genblk1.cell0_I  (.A(net501),
    .B(net435),
    .X(\col[0].zbuf_top_iw_I[14].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_top_iw_I[15].genblk1.cell0_I  (.A(net499),
    .B(net435),
    .X(\col[0].zbuf_top_iw_I[15].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_top_iw_I[16].genblk1.cell0_I  (.A(net497),
    .B(net435),
    .X(\col[0].zbuf_top_iw_I[16].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_top_iw_I[17].genblk1.cell0_I  (.A(net495),
    .B(net435),
    .X(\col[0].zbuf_top_iw_I[17].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_top_iw_I[1].genblk1.cell0_I  (.A(net493),
    .B(net436),
    .X(\col[0].zbuf_top_iw_I[1].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_top_iw_I[2].genblk1.cell0_I  (.A(net491),
    .B(net436),
    .X(\col[0].zbuf_top_iw_I[2].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_top_iw_I[3].genblk1.cell0_I  (.A(net489),
    .B(net436),
    .X(\col[0].zbuf_top_iw_I[3].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_top_iw_I[4].genblk1.cell0_I  (.A(net487),
    .B(net436),
    .X(\col[0].zbuf_top_iw_I[4].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_top_iw_I[5].genblk1.cell0_I  (.A(net485),
    .B(net436),
    .X(\col[0].zbuf_top_iw_I[5].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_top_iw_I[6].genblk1.cell0_I  (.A(net483),
    .B(net436),
    .X(\col[0].zbuf_top_iw_I[6].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_top_iw_I[7].genblk1.cell0_I  (.A(net481),
    .B(net436),
    .X(\col[0].zbuf_top_iw_I[7].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_top_iw_I[8].genblk1.cell0_I  (.A(net479),
    .B(net435),
    .X(\col[0].zbuf_top_iw_I[8].z ));
 sky130_fd_sc_hd__and2_1 \col[0].zbuf_top_iw_I[9].genblk1.cell0_I  (.A(net477),
    .B(net435),
    .X(\col[0].zbuf_top_iw_I[9].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_bot_ena_I.genblk1.cell0_I  (.A(net538),
    .B(net434),
    .X(\col[1].zbuf_bot_ena_I.z ));
 sky130_fd_sc_hd__conb_1 \col[1].zbuf_bot_ena_I.genblk1.cell0_I_538  (.HI(net538));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(net511),
    .B(net434),
    .X(\col[1].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(net509),
    .B(net433),
    .X(\col[1].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(net507),
    .B(net433),
    .X(\col[1].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(net505),
    .B(net433),
    .X(\col[1].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(net503),
    .B(net433),
    .X(\col[1].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(net501),
    .B(net433),
    .X(\col[1].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(net499),
    .B(net433),
    .X(\col[1].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(net497),
    .B(net433),
    .X(\col[1].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(net495),
    .B(net433),
    .X(\col[1].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(net493),
    .B(net434),
    .X(\col[1].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(net491),
    .B(net434),
    .X(\col[1].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(net489),
    .B(net434),
    .X(\col[1].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(net487),
    .B(net434),
    .X(\col[1].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(net485),
    .B(net434),
    .X(\col[1].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(net483),
    .B(net434),
    .X(\col[1].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(net481),
    .B(net434),
    .X(\col[1].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(net479),
    .B(net433),
    .X(\col[1].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(net477),
    .B(net433),
    .X(\col[1].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_top_ena_I.genblk1.cell0_I  (.A(net539),
    .B(net432),
    .X(\col[1].zbuf_top_ena_I.z ));
 sky130_fd_sc_hd__conb_1 \col[1].zbuf_top_ena_I.genblk1.cell0_I_539  (.HI(net539));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_top_iw_I[0].genblk1.cell0_I  (.A(net511),
    .B(net432),
    .X(\col[1].zbuf_top_iw_I[0].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_top_iw_I[10].genblk1.cell0_I  (.A(net509),
    .B(net431),
    .X(\col[1].zbuf_top_iw_I[10].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_top_iw_I[11].genblk1.cell0_I  (.A(net507),
    .B(net431),
    .X(\col[1].zbuf_top_iw_I[11].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_top_iw_I[12].genblk1.cell0_I  (.A(net505),
    .B(net431),
    .X(\col[1].zbuf_top_iw_I[12].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_top_iw_I[13].genblk1.cell0_I  (.A(net503),
    .B(net431),
    .X(\col[1].zbuf_top_iw_I[13].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_top_iw_I[14].genblk1.cell0_I  (.A(net501),
    .B(net431),
    .X(\col[1].zbuf_top_iw_I[14].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_top_iw_I[15].genblk1.cell0_I  (.A(net499),
    .B(net431),
    .X(\col[1].zbuf_top_iw_I[15].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_top_iw_I[16].genblk1.cell0_I  (.A(net497),
    .B(net431),
    .X(\col[1].zbuf_top_iw_I[16].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_top_iw_I[17].genblk1.cell0_I  (.A(net495),
    .B(net431),
    .X(\col[1].zbuf_top_iw_I[17].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_top_iw_I[1].genblk1.cell0_I  (.A(net493),
    .B(net432),
    .X(\col[1].zbuf_top_iw_I[1].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_top_iw_I[2].genblk1.cell0_I  (.A(net491),
    .B(net432),
    .X(\col[1].zbuf_top_iw_I[2].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_top_iw_I[3].genblk1.cell0_I  (.A(net489),
    .B(net432),
    .X(\col[1].zbuf_top_iw_I[3].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_top_iw_I[4].genblk1.cell0_I  (.A(net487),
    .B(net432),
    .X(\col[1].zbuf_top_iw_I[4].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_top_iw_I[5].genblk1.cell0_I  (.A(net485),
    .B(net432),
    .X(\col[1].zbuf_top_iw_I[5].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_top_iw_I[6].genblk1.cell0_I  (.A(net483),
    .B(net432),
    .X(\col[1].zbuf_top_iw_I[6].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_top_iw_I[7].genblk1.cell0_I  (.A(net481),
    .B(net432),
    .X(\col[1].zbuf_top_iw_I[7].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_top_iw_I[8].genblk1.cell0_I  (.A(net479),
    .B(net431),
    .X(\col[1].zbuf_top_iw_I[8].z ));
 sky130_fd_sc_hd__and2_1 \col[1].zbuf_top_iw_I[9].genblk1.cell0_I  (.A(net477),
    .B(net431),
    .X(\col[1].zbuf_top_iw_I[9].z ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[0].cell0_I  (.A0(net414),
    .A1(net58),
    .A2(net84),
    .A3(net110),
    .S0(net468),
    .S1(net454),
    .X(\col[2].genblk1.mux4_I[0].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[10].cell0_I  (.A0(net42),
    .A1(net69),
    .A2(net95),
    .A3(net121),
    .S0(net468),
    .S1(net454),
    .X(\col[2].genblk1.mux4_I[10].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[11].cell0_I  (.A0(net43),
    .A1(net70),
    .A2(net96),
    .A3(net122),
    .S0(net468),
    .S1(net454),
    .X(\col[2].genblk1.mux4_I[11].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[12].cell0_I  (.A0(net44),
    .A1(net71),
    .A2(net97),
    .A3(net124),
    .S0(net468),
    .S1(net454),
    .X(\col[2].genblk1.mux4_I[12].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[13].cell0_I  (.A0(net45),
    .A1(net72),
    .A2(net98),
    .A3(net125),
    .S0(net467),
    .S1(net454),
    .X(\col[2].genblk1.mux4_I[13].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[14].cell0_I  (.A0(net47),
    .A1(net73),
    .A2(net99),
    .A3(net126),
    .S0(net467),
    .S1(net456),
    .X(\col[2].genblk1.mux4_I[14].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[15].cell0_I  (.A0(net48),
    .A1(net74),
    .A2(net100),
    .A3(net127),
    .S0(net476),
    .S1(net456),
    .X(\col[2].genblk1.mux4_I[15].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[16].cell0_I  (.A0(net49),
    .A1(net75),
    .A2(net102),
    .A3(net128),
    .S0(net467),
    .S1(net456),
    .X(\col[2].genblk1.mux4_I[16].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[17].cell0_I  (.A0(net50),
    .A1(net76),
    .A2(net103),
    .A3(net129),
    .S0(net467),
    .S1(net456),
    .X(\col[2].genblk1.mux4_I[17].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[18].cell0_I  (.A0(net51),
    .A1(net77),
    .A2(net104),
    .A3(net130),
    .S0(net467),
    .S1(net456),
    .X(\col[2].genblk1.mux4_I[18].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[19].cell0_I  (.A0(net52),
    .A1(net78),
    .A2(net105),
    .A3(net131),
    .S0(net467),
    .S1(net456),
    .X(\col[2].genblk1.mux4_I[19].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[1].cell0_I  (.A0(net415),
    .A1(net59),
    .A2(net85),
    .A3(net111),
    .S0(net468),
    .S1(net454),
    .X(\col[2].genblk1.mux4_I[1].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[20].cell0_I  (.A0(net53),
    .A1(net80),
    .A2(net106),
    .A3(net132),
    .S0(net467),
    .S1(net456),
    .X(\col[2].genblk1.mux4_I[20].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[21].cell0_I  (.A0(net54),
    .A1(net81),
    .A2(net107),
    .A3(net133),
    .S0(net467),
    .S1(net456),
    .X(\col[2].genblk1.mux4_I[21].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[22].cell0_I  (.A0(net55),
    .A1(net82),
    .A2(net108),
    .A3(net135),
    .S0(net467),
    .S1(net456),
    .X(\col[2].genblk1.mux4_I[22].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[23].cell0_I  (.A0(net56),
    .A1(net83),
    .A2(net109),
    .A3(net136),
    .S0(net467),
    .S1(net456),
    .X(\col[2].genblk1.mux4_I[23].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[2].cell0_I  (.A0(net416),
    .A1(net60),
    .A2(net86),
    .A3(net113),
    .S0(net469),
    .S1(net455),
    .X(\col[2].genblk1.mux4_I[2].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[3].cell0_I  (.A0(net417),
    .A1(net61),
    .A2(net87),
    .A3(net114),
    .S0(net469),
    .S1(net455),
    .X(\col[2].genblk1.mux4_I[3].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[4].cell0_I  (.A0(net36),
    .A1(net62),
    .A2(net88),
    .A3(net115),
    .S0(net468),
    .S1(net454),
    .X(\col[2].genblk1.mux4_I[4].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[5].cell0_I  (.A0(net37),
    .A1(net63),
    .A2(net89),
    .A3(net116),
    .S0(net469),
    .S1(net455),
    .X(\col[2].genblk1.mux4_I[5].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[6].cell0_I  (.A0(net38),
    .A1(net64),
    .A2(net91),
    .A3(net117),
    .S0(net469),
    .S1(net455),
    .X(\col[2].genblk1.mux4_I[6].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[7].cell0_I  (.A0(net39),
    .A1(net65),
    .A2(net92),
    .A3(net118),
    .S0(net468),
    .S1(net454),
    .X(\col[2].genblk1.mux4_I[7].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[8].cell0_I  (.A0(net40),
    .A1(net66),
    .A2(net93),
    .A3(net119),
    .S0(net468),
    .S1(net454),
    .X(\col[2].genblk1.mux4_I[8].x ));
 sky130_fd_sc_hd__mux4_1 \col[2].genblk1.mux4_I[9].cell0_I  (.A0(net41),
    .A1(net67),
    .A2(net94),
    .A3(net120),
    .S0(net468),
    .S1(net454),
    .X(\col[2].genblk1.mux4_I[9].x ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_bot_ena_I.genblk1.cell0_I  (.A(net540),
    .B(net446),
    .X(\col[2].zbuf_bot_ena_I.z ));
 sky130_fd_sc_hd__conb_1 \col[2].zbuf_bot_ena_I.genblk1.cell0_I_540  (.HI(net540));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(net511),
    .B(net446),
    .X(\col[2].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(net509),
    .B(net445),
    .X(\col[2].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(net507),
    .B(net445),
    .X(\col[2].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(net505),
    .B(net445),
    .X(\col[2].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(net503),
    .B(net445),
    .X(\col[2].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(net501),
    .B(net445),
    .X(\col[2].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(net499),
    .B(net445),
    .X(\col[2].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(net497),
    .B(net445),
    .X(\col[2].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(net495),
    .B(net445),
    .X(\col[2].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(net493),
    .B(net446),
    .X(\col[2].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(net491),
    .B(net446),
    .X(\col[2].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(net489),
    .B(net446),
    .X(\col[2].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(net487),
    .B(net446),
    .X(\col[2].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(net485),
    .B(net446),
    .X(\col[2].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(net483),
    .B(net446),
    .X(\col[2].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(net481),
    .B(net445),
    .X(\col[2].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(net479),
    .B(net446),
    .X(\col[2].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(net477),
    .B(net445),
    .X(\col[2].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_top_ena_I.genblk1.cell0_I  (.A(net541),
    .B(net430),
    .X(\col[2].zbuf_top_ena_I.z ));
 sky130_fd_sc_hd__conb_1 \col[2].zbuf_top_ena_I.genblk1.cell0_I_541  (.HI(net541));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_top_iw_I[0].genblk1.cell0_I  (.A(net511),
    .B(net430),
    .X(\col[2].zbuf_top_iw_I[0].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_top_iw_I[10].genblk1.cell0_I  (.A(net509),
    .B(net429),
    .X(\col[2].zbuf_top_iw_I[10].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_top_iw_I[11].genblk1.cell0_I  (.A(net507),
    .B(net429),
    .X(\col[2].zbuf_top_iw_I[11].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_top_iw_I[12].genblk1.cell0_I  (.A(net505),
    .B(net429),
    .X(\col[2].zbuf_top_iw_I[12].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_top_iw_I[13].genblk1.cell0_I  (.A(net503),
    .B(net429),
    .X(\col[2].zbuf_top_iw_I[13].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_top_iw_I[14].genblk1.cell0_I  (.A(net501),
    .B(net429),
    .X(\col[2].zbuf_top_iw_I[14].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_top_iw_I[15].genblk1.cell0_I  (.A(net499),
    .B(net429),
    .X(\col[2].zbuf_top_iw_I[15].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_top_iw_I[16].genblk1.cell0_I  (.A(net497),
    .B(net429),
    .X(\col[2].zbuf_top_iw_I[16].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_top_iw_I[17].genblk1.cell0_I  (.A(net495),
    .B(net429),
    .X(\col[2].zbuf_top_iw_I[17].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_top_iw_I[1].genblk1.cell0_I  (.A(net493),
    .B(net430),
    .X(\col[2].zbuf_top_iw_I[1].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_top_iw_I[2].genblk1.cell0_I  (.A(net491),
    .B(net430),
    .X(\col[2].zbuf_top_iw_I[2].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_top_iw_I[3].genblk1.cell0_I  (.A(net489),
    .B(net430),
    .X(\col[2].zbuf_top_iw_I[3].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_top_iw_I[4].genblk1.cell0_I  (.A(net487),
    .B(net430),
    .X(\col[2].zbuf_top_iw_I[4].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_top_iw_I[5].genblk1.cell0_I  (.A(net485),
    .B(net430),
    .X(\col[2].zbuf_top_iw_I[5].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_top_iw_I[6].genblk1.cell0_I  (.A(net483),
    .B(net430),
    .X(\col[2].zbuf_top_iw_I[6].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_top_iw_I[7].genblk1.cell0_I  (.A(net481),
    .B(net430),
    .X(\col[2].zbuf_top_iw_I[7].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_top_iw_I[8].genblk1.cell0_I  (.A(net479),
    .B(net429),
    .X(\col[2].zbuf_top_iw_I[8].z ));
 sky130_fd_sc_hd__and2_1 \col[2].zbuf_top_iw_I[9].genblk1.cell0_I  (.A(net477),
    .B(net429),
    .X(\col[2].zbuf_top_iw_I[9].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_bot_ena_I.genblk1.cell0_I  (.A(net542),
    .B(net428),
    .X(\col[3].zbuf_bot_ena_I.z ));
 sky130_fd_sc_hd__conb_1 \col[3].zbuf_bot_ena_I.genblk1.cell0_I_542  (.HI(net542));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(net511),
    .B(net428),
    .X(\col[3].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(net509),
    .B(net427),
    .X(\col[3].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(net507),
    .B(net427),
    .X(\col[3].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(net505),
    .B(net427),
    .X(\col[3].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(net503),
    .B(net427),
    .X(\col[3].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(net501),
    .B(net427),
    .X(\col[3].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(net499),
    .B(net427),
    .X(\col[3].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(net497),
    .B(net427),
    .X(\col[3].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(net495),
    .B(net427),
    .X(\col[3].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(net493),
    .B(net428),
    .X(\col[3].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(net491),
    .B(net428),
    .X(\col[3].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(net489),
    .B(net428),
    .X(\col[3].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(net487),
    .B(net428),
    .X(\col[3].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(net485),
    .B(net428),
    .X(\col[3].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(net483),
    .B(net428),
    .X(\col[3].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(net481),
    .B(net428),
    .X(\col[3].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(net479),
    .B(net427),
    .X(\col[3].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(net477),
    .B(net427),
    .X(\col[3].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_top_ena_I.genblk1.cell0_I  (.A(net543),
    .B(net425),
    .X(\col[3].zbuf_top_ena_I.z ));
 sky130_fd_sc_hd__conb_1 \col[3].zbuf_top_ena_I.genblk1.cell0_I_543  (.HI(net543));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_top_iw_I[0].genblk1.cell0_I  (.A(net511),
    .B(net426),
    .X(\col[3].zbuf_top_iw_I[0].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_top_iw_I[10].genblk1.cell0_I  (.A(net509),
    .B(net425),
    .X(\col[3].zbuf_top_iw_I[10].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_top_iw_I[11].genblk1.cell0_I  (.A(net507),
    .B(net425),
    .X(\col[3].zbuf_top_iw_I[11].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_top_iw_I[12].genblk1.cell0_I  (.A(net505),
    .B(net425),
    .X(\col[3].zbuf_top_iw_I[12].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_top_iw_I[13].genblk1.cell0_I  (.A(net503),
    .B(net425),
    .X(\col[3].zbuf_top_iw_I[13].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_top_iw_I[14].genblk1.cell0_I  (.A(net501),
    .B(net425),
    .X(\col[3].zbuf_top_iw_I[14].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_top_iw_I[15].genblk1.cell0_I  (.A(net499),
    .B(net425),
    .X(\col[3].zbuf_top_iw_I[15].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_top_iw_I[16].genblk1.cell0_I  (.A(net497),
    .B(net425),
    .X(\col[3].zbuf_top_iw_I[16].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_top_iw_I[17].genblk1.cell0_I  (.A(net495),
    .B(net425),
    .X(\col[3].zbuf_top_iw_I[17].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_top_iw_I[1].genblk1.cell0_I  (.A(net493),
    .B(net426),
    .X(\col[3].zbuf_top_iw_I[1].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_top_iw_I[2].genblk1.cell0_I  (.A(net491),
    .B(net426),
    .X(\col[3].zbuf_top_iw_I[2].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_top_iw_I[3].genblk1.cell0_I  (.A(net489),
    .B(net426),
    .X(\col[3].zbuf_top_iw_I[3].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_top_iw_I[4].genblk1.cell0_I  (.A(net487),
    .B(net426),
    .X(\col[3].zbuf_top_iw_I[4].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_top_iw_I[5].genblk1.cell0_I  (.A(net485),
    .B(net426),
    .X(\col[3].zbuf_top_iw_I[5].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_top_iw_I[6].genblk1.cell0_I  (.A(net483),
    .B(net426),
    .X(\col[3].zbuf_top_iw_I[6].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_top_iw_I[7].genblk1.cell0_I  (.A(net481),
    .B(net426),
    .X(\col[3].zbuf_top_iw_I[7].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_top_iw_I[8].genblk1.cell0_I  (.A(net479),
    .B(net426),
    .X(\col[3].zbuf_top_iw_I[8].z ));
 sky130_fd_sc_hd__and2_1 \col[3].zbuf_top_iw_I[9].genblk1.cell0_I  (.A(net477),
    .B(net425),
    .X(\col[3].zbuf_top_iw_I[9].z ));
 sky130_fd_sc_hd__mux4_2 \col[4].genblk1.mux4_I[0].cell0_I  (.A0(net137),
    .A1(net164),
    .A2(net191),
    .A3(net217),
    .S0(net472),
    .S1(net459),
    .X(\col[4].genblk1.mux4_I[0].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[10].cell0_I  (.A0(net149),
    .A1(net175),
    .A2(net202),
    .A3(net228),
    .S0(net470),
    .S1(net457),
    .X(\col[4].genblk1.mux4_I[10].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[11].cell0_I  (.A0(net150),
    .A1(net176),
    .A2(net203),
    .A3(net229),
    .S0(net471),
    .S1(net457),
    .X(\col[4].genblk1.mux4_I[11].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[12].cell0_I  (.A0(net151),
    .A1(net177),
    .A2(net204),
    .A3(net230),
    .S0(net471),
    .S1(net458),
    .X(\col[4].genblk1.mux4_I[12].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[13].cell0_I  (.A0(net152),
    .A1(net178),
    .A2(net205),
    .A3(net231),
    .S0(net470),
    .S1(net457),
    .X(\col[4].genblk1.mux4_I[13].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[14].cell0_I  (.A0(net153),
    .A1(net180),
    .A2(net206),
    .A3(net232),
    .S0(net470),
    .S1(net457),
    .X(\col[4].genblk1.mux4_I[14].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[15].cell0_I  (.A0(net154),
    .A1(net181),
    .A2(net207),
    .A3(net233),
    .S0(net470),
    .S1(net457),
    .X(\col[4].genblk1.mux4_I[15].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[16].cell0_I  (.A0(net155),
    .A1(net182),
    .A2(net208),
    .A3(net235),
    .S0(net470),
    .S1(net457),
    .X(\col[4].genblk1.mux4_I[16].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[17].cell0_I  (.A0(net156),
    .A1(net183),
    .A2(net209),
    .A3(net236),
    .S0(net470),
    .S1(net457),
    .X(\col[4].genblk1.mux4_I[17].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[18].cell0_I  (.A0(net158),
    .A1(net184),
    .A2(net210),
    .A3(net237),
    .S0(net470),
    .S1(net457),
    .X(\col[4].genblk1.mux4_I[18].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[19].cell0_I  (.A0(net159),
    .A1(net185),
    .A2(net211),
    .A3(net238),
    .S0(net471),
    .S1(net458),
    .X(\col[4].genblk1.mux4_I[19].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[1].cell0_I  (.A0(net138),
    .A1(net165),
    .A2(net192),
    .A3(net218),
    .S0(net472),
    .S1(net459),
    .X(\col[4].genblk1.mux4_I[1].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[20].cell0_I  (.A0(net160),
    .A1(net186),
    .A2(net213),
    .A3(net239),
    .S0(net471),
    .S1(net458),
    .X(\col[4].genblk1.mux4_I[20].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[21].cell0_I  (.A0(net161),
    .A1(net187),
    .A2(net214),
    .A3(net240),
    .S0(net471),
    .S1(net458),
    .X(\col[4].genblk1.mux4_I[21].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[22].cell0_I  (.A0(net162),
    .A1(net188),
    .A2(net215),
    .A3(net241),
    .S0(net471),
    .S1(net458),
    .X(\col[4].genblk1.mux4_I[22].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[23].cell0_I  (.A0(net163),
    .A1(net189),
    .A2(net216),
    .A3(net242),
    .S0(net471),
    .S1(net458),
    .X(\col[4].genblk1.mux4_I[23].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[2].cell0_I  (.A0(net139),
    .A1(net166),
    .A2(net193),
    .A3(net219),
    .S0(net472),
    .S1(net459),
    .X(\col[4].genblk1.mux4_I[2].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[3].cell0_I  (.A0(net140),
    .A1(net167),
    .A2(net194),
    .A3(net220),
    .S0(net472),
    .S1(net459),
    .X(\col[4].genblk1.mux4_I[3].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[4].cell0_I  (.A0(net141),
    .A1(net169),
    .A2(net195),
    .A3(net221),
    .S0(net472),
    .S1(net459),
    .X(\col[4].genblk1.mux4_I[4].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[5].cell0_I  (.A0(net142),
    .A1(net170),
    .A2(net196),
    .A3(net222),
    .S0(net472),
    .S1(net459),
    .X(\col[4].genblk1.mux4_I[5].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[6].cell0_I  (.A0(net143),
    .A1(net171),
    .A2(net197),
    .A3(net224),
    .S0(net470),
    .S1(net457),
    .X(\col[4].genblk1.mux4_I[6].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[7].cell0_I  (.A0(net144),
    .A1(net172),
    .A2(net198),
    .A3(net225),
    .S0(net470),
    .S1(net457),
    .X(\col[4].genblk1.mux4_I[7].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[8].cell0_I  (.A0(net147),
    .A1(net173),
    .A2(net199),
    .A3(net226),
    .S0(net470),
    .S1(net458),
    .X(\col[4].genblk1.mux4_I[8].x ));
 sky130_fd_sc_hd__mux4_1 \col[4].genblk1.mux4_I[9].cell0_I  (.A0(net148),
    .A1(net174),
    .A2(net200),
    .A3(net227),
    .S0(net471),
    .S1(net458),
    .X(\col[4].genblk1.mux4_I[9].x ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_bot_ena_I.genblk1.cell0_I  (.A(net544),
    .B(net444),
    .X(\col[4].zbuf_bot_ena_I.z ));
 sky130_fd_sc_hd__conb_1 \col[4].zbuf_bot_ena_I.genblk1.cell0_I_544  (.HI(net544));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(net511),
    .B(net444),
    .X(\col[4].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(net509),
    .B(net443),
    .X(\col[4].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(net507),
    .B(net443),
    .X(\col[4].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(net505),
    .B(net443),
    .X(\col[4].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(net503),
    .B(net443),
    .X(\col[4].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(net501),
    .B(net443),
    .X(\col[4].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(net499),
    .B(net443),
    .X(\col[4].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(net497),
    .B(net443),
    .X(\col[4].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(net495),
    .B(net443),
    .X(\col[4].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(net493),
    .B(net444),
    .X(\col[4].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(net491),
    .B(net444),
    .X(\col[4].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(net489),
    .B(net444),
    .X(\col[4].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(net487),
    .B(net444),
    .X(\col[4].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(net485),
    .B(net444),
    .X(\col[4].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(net483),
    .B(net444),
    .X(\col[4].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(net481),
    .B(net444),
    .X(\col[4].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(net479),
    .B(net443),
    .X(\col[4].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(net477),
    .B(net443),
    .X(\col[4].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_top_ena_I.genblk1.cell0_I  (.A(net545),
    .B(net424),
    .X(\col[4].zbuf_top_ena_I.z ));
 sky130_fd_sc_hd__conb_1 \col[4].zbuf_top_ena_I.genblk1.cell0_I_545  (.HI(net545));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_top_iw_I[0].genblk1.cell0_I  (.A(net511),
    .B(net424),
    .X(\col[4].zbuf_top_iw_I[0].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_top_iw_I[10].genblk1.cell0_I  (.A(net509),
    .B(net423),
    .X(\col[4].zbuf_top_iw_I[10].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_top_iw_I[11].genblk1.cell0_I  (.A(net507),
    .B(net423),
    .X(\col[4].zbuf_top_iw_I[11].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_top_iw_I[12].genblk1.cell0_I  (.A(net505),
    .B(net423),
    .X(\col[4].zbuf_top_iw_I[12].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_top_iw_I[13].genblk1.cell0_I  (.A(net503),
    .B(net423),
    .X(\col[4].zbuf_top_iw_I[13].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_top_iw_I[14].genblk1.cell0_I  (.A(net501),
    .B(net423),
    .X(\col[4].zbuf_top_iw_I[14].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_top_iw_I[15].genblk1.cell0_I  (.A(net499),
    .B(net423),
    .X(\col[4].zbuf_top_iw_I[15].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_top_iw_I[16].genblk1.cell0_I  (.A(net497),
    .B(net423),
    .X(\col[4].zbuf_top_iw_I[16].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_top_iw_I[17].genblk1.cell0_I  (.A(net495),
    .B(net423),
    .X(\col[4].zbuf_top_iw_I[17].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_top_iw_I[1].genblk1.cell0_I  (.A(net493),
    .B(net424),
    .X(\col[4].zbuf_top_iw_I[1].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_top_iw_I[2].genblk1.cell0_I  (.A(net491),
    .B(net424),
    .X(\col[4].zbuf_top_iw_I[2].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_top_iw_I[3].genblk1.cell0_I  (.A(net489),
    .B(net424),
    .X(\col[4].zbuf_top_iw_I[3].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_top_iw_I[4].genblk1.cell0_I  (.A(net487),
    .B(net424),
    .X(\col[4].zbuf_top_iw_I[4].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_top_iw_I[5].genblk1.cell0_I  (.A(net485),
    .B(net424),
    .X(\col[4].zbuf_top_iw_I[5].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_top_iw_I[6].genblk1.cell0_I  (.A(net483),
    .B(net424),
    .X(\col[4].zbuf_top_iw_I[6].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_top_iw_I[7].genblk1.cell0_I  (.A(net481),
    .B(net424),
    .X(\col[4].zbuf_top_iw_I[7].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_top_iw_I[8].genblk1.cell0_I  (.A(net479),
    .B(net423),
    .X(\col[4].zbuf_top_iw_I[8].z ));
 sky130_fd_sc_hd__and2_1 \col[4].zbuf_top_iw_I[9].genblk1.cell0_I  (.A(net477),
    .B(net423),
    .X(\col[4].zbuf_top_iw_I[9].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_bot_ena_I.genblk1.cell0_I  (.A(net546),
    .B(net422),
    .X(\col[5].zbuf_bot_ena_I.z ));
 sky130_fd_sc_hd__conb_1 \col[5].zbuf_bot_ena_I.genblk1.cell0_I_546  (.HI(net546));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(net512),
    .B(net422),
    .X(\col[5].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(net510),
    .B(net421),
    .X(\col[5].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(net508),
    .B(net421),
    .X(\col[5].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(net506),
    .B(net421),
    .X(\col[5].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(net504),
    .B(net421),
    .X(\col[5].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(net502),
    .B(net421),
    .X(\col[5].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(net500),
    .B(net421),
    .X(\col[5].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(net498),
    .B(net421),
    .X(\col[5].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(net496),
    .B(net421),
    .X(\col[5].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(net494),
    .B(net422),
    .X(\col[5].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(net492),
    .B(net422),
    .X(\col[5].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(net490),
    .B(net422),
    .X(\col[5].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(net488),
    .B(net422),
    .X(\col[5].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(net486),
    .B(net422),
    .X(\col[5].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(net484),
    .B(net422),
    .X(\col[5].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(net482),
    .B(net422),
    .X(\col[5].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(net480),
    .B(net421),
    .X(\col[5].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(net478),
    .B(net421),
    .X(\col[5].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_top_ena_I.genblk1.cell0_I  (.A(net547),
    .B(net420),
    .X(\col[5].zbuf_top_ena_I.z ));
 sky130_fd_sc_hd__conb_1 \col[5].zbuf_top_ena_I.genblk1.cell0_I_547  (.HI(net547));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_top_iw_I[0].genblk1.cell0_I  (.A(net512),
    .B(net420),
    .X(\col[5].zbuf_top_iw_I[0].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_top_iw_I[10].genblk1.cell0_I  (.A(net510),
    .B(net419),
    .X(\col[5].zbuf_top_iw_I[10].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_top_iw_I[11].genblk1.cell0_I  (.A(net508),
    .B(net419),
    .X(\col[5].zbuf_top_iw_I[11].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_top_iw_I[12].genblk1.cell0_I  (.A(net506),
    .B(net419),
    .X(\col[5].zbuf_top_iw_I[12].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_top_iw_I[13].genblk1.cell0_I  (.A(net504),
    .B(net419),
    .X(\col[5].zbuf_top_iw_I[13].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_top_iw_I[14].genblk1.cell0_I  (.A(net502),
    .B(net419),
    .X(\col[5].zbuf_top_iw_I[14].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_top_iw_I[15].genblk1.cell0_I  (.A(net500),
    .B(net419),
    .X(\col[5].zbuf_top_iw_I[15].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_top_iw_I[16].genblk1.cell0_I  (.A(net498),
    .B(net419),
    .X(\col[5].zbuf_top_iw_I[16].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_top_iw_I[17].genblk1.cell0_I  (.A(net496),
    .B(net419),
    .X(\col[5].zbuf_top_iw_I[17].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_top_iw_I[1].genblk1.cell0_I  (.A(net494),
    .B(net420),
    .X(\col[5].zbuf_top_iw_I[1].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_top_iw_I[2].genblk1.cell0_I  (.A(net492),
    .B(net420),
    .X(\col[5].zbuf_top_iw_I[2].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_top_iw_I[3].genblk1.cell0_I  (.A(net490),
    .B(net420),
    .X(\col[5].zbuf_top_iw_I[3].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_top_iw_I[4].genblk1.cell0_I  (.A(net488),
    .B(net420),
    .X(\col[5].zbuf_top_iw_I[4].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_top_iw_I[5].genblk1.cell0_I  (.A(net486),
    .B(net420),
    .X(\col[5].zbuf_top_iw_I[5].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_top_iw_I[6].genblk1.cell0_I  (.A(net484),
    .B(net420),
    .X(\col[5].zbuf_top_iw_I[6].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_top_iw_I[7].genblk1.cell0_I  (.A(net482),
    .B(net420),
    .X(\col[5].zbuf_top_iw_I[7].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_top_iw_I[8].genblk1.cell0_I  (.A(net480),
    .B(net419),
    .X(\col[5].zbuf_top_iw_I[8].z ));
 sky130_fd_sc_hd__and2_1 \col[5].zbuf_top_iw_I[9].genblk1.cell0_I  (.A(net478),
    .B(net419),
    .X(\col[5].zbuf_top_iw_I[9].z ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[0].cell0_I  (.A0(net243),
    .A1(net271),
    .A2(net297),
    .A3(net324),
    .S0(net473),
    .S1(net460),
    .X(\col[6].genblk1.mux4_I[0].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[10].cell0_I  (.A0(net254),
    .A1(net282),
    .A2(net308),
    .A3(net335),
    .S0(net474),
    .S1(net461),
    .X(\col[6].genblk1.mux4_I[10].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[11].cell0_I  (.A0(net255),
    .A1(net283),
    .A2(net309),
    .A3(net336),
    .S0(net473),
    .S1(net460),
    .X(\col[6].genblk1.mux4_I[11].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[12].cell0_I  (.A0(net258),
    .A1(net284),
    .A2(net310),
    .A3(net337),
    .S0(net474),
    .S1(net461),
    .X(\col[6].genblk1.mux4_I[12].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[13].cell0_I  (.A0(net259),
    .A1(net285),
    .A2(net311),
    .A3(net338),
    .S0(net474),
    .S1(net461),
    .X(\col[6].genblk1.mux4_I[13].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[14].cell0_I  (.A0(net260),
    .A1(net286),
    .A2(net313),
    .A3(net339),
    .S0(net474),
    .S1(net461),
    .X(\col[6].genblk1.mux4_I[14].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[15].cell0_I  (.A0(net261),
    .A1(net287),
    .A2(net314),
    .A3(net340),
    .S0(net474),
    .S1(net461),
    .X(\col[6].genblk1.mux4_I[15].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[16].cell0_I  (.A0(net262),
    .A1(net288),
    .A2(net315),
    .A3(net341),
    .S0(net474),
    .S1(net461),
    .X(\col[6].genblk1.mux4_I[16].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[17].cell0_I  (.A0(net263),
    .A1(net289),
    .A2(net316),
    .A3(net342),
    .S0(net475),
    .S1(net462),
    .X(\col[6].genblk1.mux4_I[17].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[18].cell0_I  (.A0(net264),
    .A1(net291),
    .A2(net317),
    .A3(net343),
    .S0(net475),
    .S1(net462),
    .X(\col[6].genblk1.mux4_I[18].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[19].cell0_I  (.A0(net265),
    .A1(net292),
    .A2(net318),
    .A3(net344),
    .S0(net475),
    .S1(net462),
    .X(\col[6].genblk1.mux4_I[19].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[1].cell0_I  (.A0(net244),
    .A1(net272),
    .A2(net298),
    .A3(net325),
    .S0(net473),
    .S1(net460),
    .X(\col[6].genblk1.mux4_I[1].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[20].cell0_I  (.A0(net266),
    .A1(net293),
    .A2(net319),
    .A3(net346),
    .S0(net475),
    .S1(net462),
    .X(\col[6].genblk1.mux4_I[20].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[21].cell0_I  (.A0(net267),
    .A1(net294),
    .A2(net320),
    .A3(net347),
    .S0(net475),
    .S1(net462),
    .X(\col[6].genblk1.mux4_I[21].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[22].cell0_I  (.A0(net269),
    .A1(net295),
    .A2(net321),
    .A3(net348),
    .S0(net475),
    .S1(net462),
    .X(\col[6].genblk1.mux4_I[22].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[23].cell0_I  (.A0(net270),
    .A1(net296),
    .A2(net322),
    .A3(net349),
    .S0(net475),
    .S1(net462),
    .X(\col[6].genblk1.mux4_I[23].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[2].cell0_I  (.A0(net246),
    .A1(net273),
    .A2(net299),
    .A3(net326),
    .S0(net473),
    .S1(net460),
    .X(\col[6].genblk1.mux4_I[2].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[3].cell0_I  (.A0(net247),
    .A1(net274),
    .A2(net300),
    .A3(net327),
    .S0(net473),
    .S1(net460),
    .X(\col[6].genblk1.mux4_I[3].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[4].cell0_I  (.A0(net248),
    .A1(net275),
    .A2(net302),
    .A3(net328),
    .S0(net473),
    .S1(net461),
    .X(\col[6].genblk1.mux4_I[4].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[5].cell0_I  (.A0(net249),
    .A1(net276),
    .A2(net303),
    .A3(net329),
    .S0(net473),
    .S1(net460),
    .X(\col[6].genblk1.mux4_I[5].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[6].cell0_I  (.A0(net250),
    .A1(net277),
    .A2(net304),
    .A3(net330),
    .S0(net473),
    .S1(net460),
    .X(\col[6].genblk1.mux4_I[6].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[7].cell0_I  (.A0(net251),
    .A1(net278),
    .A2(net305),
    .A3(net331),
    .S0(net473),
    .S1(net460),
    .X(\col[6].genblk1.mux4_I[7].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[8].cell0_I  (.A0(net252),
    .A1(net280),
    .A2(net306),
    .A3(net332),
    .S0(net473),
    .S1(net460),
    .X(\col[6].genblk1.mux4_I[8].x ));
 sky130_fd_sc_hd__mux4_1 \col[6].genblk1.mux4_I[9].cell0_I  (.A0(net253),
    .A1(net281),
    .A2(net307),
    .A3(net333),
    .S0(net474),
    .S1(net461),
    .X(\col[6].genblk1.mux4_I[9].x ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_bot_ena_I.genblk1.cell0_I  (.A(net548),
    .B(net450),
    .X(\col[6].zbuf_bot_ena_I.z ));
 sky130_fd_sc_hd__conb_1 \col[6].zbuf_bot_ena_I.genblk1.cell0_I_548  (.HI(net548));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(net512),
    .B(net449),
    .X(\col[6].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(net510),
    .B(net450),
    .X(\col[6].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(net508),
    .B(net450),
    .X(\col[6].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(net506),
    .B(net450),
    .X(\col[6].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(net504),
    .B(net450),
    .X(\col[6].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(net502),
    .B(net450),
    .X(\col[6].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(net500),
    .B(net450),
    .X(\col[6].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(net498),
    .B(net450),
    .X(\col[6].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(net496),
    .B(net450),
    .X(\col[6].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(net494),
    .B(net449),
    .X(\col[6].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(net492),
    .B(net449),
    .X(\col[6].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(net490),
    .B(net449),
    .X(\col[6].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(net488),
    .B(net449),
    .X(\col[6].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(net486),
    .B(net449),
    .X(\col[6].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(net484),
    .B(net449),
    .X(\col[6].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(net482),
    .B(net449),
    .X(\col[6].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(net480),
    .B(net449),
    .X(\col[6].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(net478),
    .B(net449),
    .X(\col[6].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_top_ena_I.genblk1.cell0_I  (.A(net549),
    .B(net441),
    .X(\col[6].zbuf_top_ena_I.z ));
 sky130_fd_sc_hd__conb_1 \col[6].zbuf_top_ena_I.genblk1.cell0_I_549  (.HI(net549));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_top_iw_I[0].genblk1.cell0_I  (.A(net512),
    .B(net442),
    .X(\col[6].zbuf_top_iw_I[0].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_top_iw_I[10].genblk1.cell0_I  (.A(net510),
    .B(net441),
    .X(\col[6].zbuf_top_iw_I[10].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_top_iw_I[11].genblk1.cell0_I  (.A(net508),
    .B(net441),
    .X(\col[6].zbuf_top_iw_I[11].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_top_iw_I[12].genblk1.cell0_I  (.A(net506),
    .B(net441),
    .X(\col[6].zbuf_top_iw_I[12].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_top_iw_I[13].genblk1.cell0_I  (.A(net504),
    .B(net441),
    .X(\col[6].zbuf_top_iw_I[13].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_top_iw_I[14].genblk1.cell0_I  (.A(net502),
    .B(net441),
    .X(\col[6].zbuf_top_iw_I[14].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_top_iw_I[15].genblk1.cell0_I  (.A(net500),
    .B(net441),
    .X(\col[6].zbuf_top_iw_I[15].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_top_iw_I[16].genblk1.cell0_I  (.A(net498),
    .B(net441),
    .X(\col[6].zbuf_top_iw_I[16].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_top_iw_I[17].genblk1.cell0_I  (.A(net496),
    .B(net441),
    .X(\col[6].zbuf_top_iw_I[17].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_top_iw_I[1].genblk1.cell0_I  (.A(net494),
    .B(net442),
    .X(\col[6].zbuf_top_iw_I[1].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_top_iw_I[2].genblk1.cell0_I  (.A(net492),
    .B(net442),
    .X(\col[6].zbuf_top_iw_I[2].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_top_iw_I[3].genblk1.cell0_I  (.A(net490),
    .B(net442),
    .X(\col[6].zbuf_top_iw_I[3].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_top_iw_I[4].genblk1.cell0_I  (.A(net488),
    .B(net442),
    .X(\col[6].zbuf_top_iw_I[4].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_top_iw_I[5].genblk1.cell0_I  (.A(net486),
    .B(net442),
    .X(\col[6].zbuf_top_iw_I[5].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_top_iw_I[6].genblk1.cell0_I  (.A(net484),
    .B(net442),
    .X(\col[6].zbuf_top_iw_I[6].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_top_iw_I[7].genblk1.cell0_I  (.A(net482),
    .B(net442),
    .X(\col[6].zbuf_top_iw_I[7].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_top_iw_I[8].genblk1.cell0_I  (.A(net480),
    .B(net442),
    .X(\col[6].zbuf_top_iw_I[8].z ));
 sky130_fd_sc_hd__and2_1 \col[6].zbuf_top_iw_I[9].genblk1.cell0_I  (.A(net478),
    .B(net441),
    .X(\col[6].zbuf_top_iw_I[9].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_bot_ena_I.genblk1.cell0_I  (.A(net550),
    .B(net440),
    .X(\col[7].zbuf_bot_ena_I.z ));
 sky130_fd_sc_hd__conb_1 \col[7].zbuf_bot_ena_I.genblk1.cell0_I_550  (.HI(net550));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(net512),
    .B(net440),
    .X(\col[7].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(net510),
    .B(net439),
    .X(\col[7].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(net508),
    .B(net439),
    .X(\col[7].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(net506),
    .B(net439),
    .X(\col[7].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(net504),
    .B(net439),
    .X(\col[7].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(net502),
    .B(net439),
    .X(\col[7].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(net500),
    .B(net439),
    .X(\col[7].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(net498),
    .B(net439),
    .X(\col[7].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(net496),
    .B(net439),
    .X(\col[7].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(net494),
    .B(net440),
    .X(\col[7].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(net492),
    .B(net440),
    .X(\col[7].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(net490),
    .B(net440),
    .X(\col[7].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(net488),
    .B(net440),
    .X(\col[7].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(net486),
    .B(net440),
    .X(\col[7].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(net484),
    .B(net440),
    .X(\col[7].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(net482),
    .B(net440),
    .X(\col[7].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(net480),
    .B(net439),
    .X(\col[7].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(net478),
    .B(net439),
    .X(\col[7].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_top_ena_I.genblk1.cell0_I  (.A(net551),
    .B(net438),
    .X(\col[7].zbuf_top_ena_I.z ));
 sky130_fd_sc_hd__conb_1 \col[7].zbuf_top_ena_I.genblk1.cell0_I_551  (.HI(net551));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_top_iw_I[0].genblk1.cell0_I  (.A(net512),
    .B(net438),
    .X(\col[7].zbuf_top_iw_I[0].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_top_iw_I[10].genblk1.cell0_I  (.A(net510),
    .B(net437),
    .X(\col[7].zbuf_top_iw_I[10].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_top_iw_I[11].genblk1.cell0_I  (.A(net508),
    .B(net437),
    .X(\col[7].zbuf_top_iw_I[11].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_top_iw_I[12].genblk1.cell0_I  (.A(net506),
    .B(net437),
    .X(\col[7].zbuf_top_iw_I[12].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_top_iw_I[13].genblk1.cell0_I  (.A(net504),
    .B(net437),
    .X(\col[7].zbuf_top_iw_I[13].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_top_iw_I[14].genblk1.cell0_I  (.A(net502),
    .B(net437),
    .X(\col[7].zbuf_top_iw_I[14].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_top_iw_I[15].genblk1.cell0_I  (.A(net500),
    .B(net437),
    .X(\col[7].zbuf_top_iw_I[15].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_top_iw_I[16].genblk1.cell0_I  (.A(net498),
    .B(net437),
    .X(\col[7].zbuf_top_iw_I[16].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_top_iw_I[17].genblk1.cell0_I  (.A(net496),
    .B(net437),
    .X(\col[7].zbuf_top_iw_I[17].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_top_iw_I[1].genblk1.cell0_I  (.A(net494),
    .B(net438),
    .X(\col[7].zbuf_top_iw_I[1].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_top_iw_I[2].genblk1.cell0_I  (.A(net492),
    .B(net438),
    .X(\col[7].zbuf_top_iw_I[2].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_top_iw_I[3].genblk1.cell0_I  (.A(net490),
    .B(net438),
    .X(\col[7].zbuf_top_iw_I[3].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_top_iw_I[4].genblk1.cell0_I  (.A(net488),
    .B(net438),
    .X(\col[7].zbuf_top_iw_I[4].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_top_iw_I[5].genblk1.cell0_I  (.A(net486),
    .B(net437),
    .X(\col[7].zbuf_top_iw_I[5].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_top_iw_I[6].genblk1.cell0_I  (.A(net484),
    .B(net438),
    .X(\col[7].zbuf_top_iw_I[6].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_top_iw_I[7].genblk1.cell0_I  (.A(net482),
    .B(net438),
    .X(\col[7].zbuf_top_iw_I[7].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_top_iw_I[8].genblk1.cell0_I  (.A(net480),
    .B(net438),
    .X(\col[7].zbuf_top_iw_I[8].z ));
 sky130_fd_sc_hd__and2_1 \col[7].zbuf_top_iw_I[9].genblk1.cell0_I  (.A(net478),
    .B(net437),
    .X(\col[7].zbuf_top_iw_I[9].z ));
 sky130_fd_sc_hd__clkbuf_2 fanout419 (.A(\col[5].zbuf_top_ena_I.e ),
    .X(net419));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout420 (.A(\col[5].zbuf_top_ena_I.e ),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_2 fanout421 (.A(\col[5].zbuf_bot_ena_I.e ),
    .X(net421));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout422 (.A(\col[5].zbuf_bot_ena_I.e ),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_2 fanout423 (.A(\col[4].zbuf_top_ena_I.e ),
    .X(net423));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout424 (.A(\col[4].zbuf_top_ena_I.e ),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_2 fanout425 (.A(\col[3].zbuf_top_ena_I.e ),
    .X(net425));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout426 (.A(\col[3].zbuf_top_ena_I.e ),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_2 fanout427 (.A(\col[3].zbuf_bot_ena_I.e ),
    .X(net427));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout428 (.A(\col[3].zbuf_bot_ena_I.e ),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_2 fanout429 (.A(\col[2].zbuf_top_ena_I.e ),
    .X(net429));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout430 (.A(\col[2].zbuf_top_ena_I.e ),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_2 fanout431 (.A(\col[1].zbuf_top_ena_I.e ),
    .X(net431));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout432 (.A(\col[1].zbuf_top_ena_I.e ),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_2 fanout433 (.A(\col[1].zbuf_bot_ena_I.e ),
    .X(net433));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout434 (.A(\col[1].zbuf_bot_ena_I.e ),
    .X(net434));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout435 (.A(net436),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_2 fanout436 (.A(\col[0].zbuf_top_ena_I.e ),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_2 fanout437 (.A(\col[7].zbuf_top_ena_I.e ),
    .X(net437));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout438 (.A(\col[7].zbuf_top_ena_I.e ),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_2 fanout439 (.A(\col[7].zbuf_bot_ena_I.e ),
    .X(net439));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout440 (.A(\col[7].zbuf_bot_ena_I.e ),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_2 fanout441 (.A(\col[6].zbuf_top_ena_I.e ),
    .X(net441));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout442 (.A(\col[6].zbuf_top_ena_I.e ),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_2 fanout443 (.A(\col[4].zbuf_bot_ena_I.e ),
    .X(net443));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout444 (.A(\col[4].zbuf_bot_ena_I.e ),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_2 fanout445 (.A(\col[2].zbuf_bot_ena_I.e ),
    .X(net445));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout446 (.A(\col[2].zbuf_bot_ena_I.e ),
    .X(net446));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_2 fanout448 (.A(\col[0].zbuf_bot_ena_I.e ),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_2 fanout449 (.A(net450),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_2 fanout450 (.A(\col[6].zbuf_bot_ena_I.e ),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_4 fanout451 (.A(net453),
    .X(net451));
 sky130_fd_sc_hd__buf_2 fanout452 (.A(net453),
    .X(net452));
 sky130_fd_sc_hd__buf_2 fanout453 (.A(net463),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_4 fanout454 (.A(net455),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_2 fanout455 (.A(net463),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_4 fanout456 (.A(net463),
    .X(net456));
 sky130_fd_sc_hd__buf_2 fanout457 (.A(net458),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_4 fanout458 (.A(net459),
    .X(net458));
 sky130_fd_sc_hd__buf_2 fanout459 (.A(net463),
    .X(net459));
 sky130_fd_sc_hd__buf_2 fanout460 (.A(net461),
    .X(net460));
 sky130_fd_sc_hd__buf_2 fanout461 (.A(net462),
    .X(net461));
 sky130_fd_sc_hd__buf_2 fanout462 (.A(net463),
    .X(net462));
 sky130_fd_sc_hd__buf_6 fanout463 (.A(\zbuf_bus_sel_I[1].z ),
    .X(net463));
 sky130_fd_sc_hd__buf_4 fanout464 (.A(net466),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_4 fanout465 (.A(net466),
    .X(net465));
 sky130_fd_sc_hd__buf_4 fanout466 (.A(net476),
    .X(net466));
 sky130_fd_sc_hd__buf_4 fanout467 (.A(net476),
    .X(net467));
 sky130_fd_sc_hd__clkbuf_4 fanout468 (.A(net469),
    .X(net468));
 sky130_fd_sc_hd__clkbuf_2 fanout469 (.A(net476),
    .X(net469));
 sky130_fd_sc_hd__buf_4 fanout470 (.A(net471),
    .X(net470));
 sky130_fd_sc_hd__buf_4 fanout471 (.A(net472),
    .X(net471));
 sky130_fd_sc_hd__clkbuf_4 fanout472 (.A(net476),
    .X(net472));
 sky130_fd_sc_hd__clkbuf_4 fanout473 (.A(net474),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_4 fanout474 (.A(net475),
    .X(net474));
 sky130_fd_sc_hd__clkbuf_4 fanout475 (.A(net476),
    .X(net475));
 sky130_fd_sc_hd__buf_8 fanout476 (.A(\zbuf_bus_sel_I[0].z ),
    .X(net476));
 sky130_fd_sc_hd__buf_6 fanout477 (.A(\col[0].zbuf_bot_iw_I[9].a ),
    .X(net477));
 sky130_fd_sc_hd__clkbuf_4 fanout478 (.A(\col[0].zbuf_bot_iw_I[9].a ),
    .X(net478));
 sky130_fd_sc_hd__buf_6 fanout479 (.A(\col[0].zbuf_bot_iw_I[8].a ),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_4 fanout480 (.A(\col[0].zbuf_bot_iw_I[8].a ),
    .X(net480));
 sky130_fd_sc_hd__buf_6 fanout481 (.A(\col[0].zbuf_bot_iw_I[7].a ),
    .X(net481));
 sky130_fd_sc_hd__clkbuf_4 fanout482 (.A(\col[0].zbuf_bot_iw_I[7].a ),
    .X(net482));
 sky130_fd_sc_hd__buf_6 fanout483 (.A(\col[0].zbuf_bot_iw_I[6].a ),
    .X(net483));
 sky130_fd_sc_hd__clkbuf_4 fanout484 (.A(\col[0].zbuf_bot_iw_I[6].a ),
    .X(net484));
 sky130_fd_sc_hd__buf_6 fanout485 (.A(\col[0].zbuf_bot_iw_I[5].a ),
    .X(net485));
 sky130_fd_sc_hd__clkbuf_4 fanout486 (.A(\col[0].zbuf_bot_iw_I[5].a ),
    .X(net486));
 sky130_fd_sc_hd__buf_6 fanout487 (.A(\col[0].zbuf_bot_iw_I[4].a ),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_4 fanout488 (.A(\col[0].zbuf_bot_iw_I[4].a ),
    .X(net488));
 sky130_fd_sc_hd__buf_6 fanout489 (.A(\col[0].zbuf_bot_iw_I[3].a ),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_4 fanout490 (.A(\col[0].zbuf_bot_iw_I[3].a ),
    .X(net490));
 sky130_fd_sc_hd__buf_6 fanout491 (.A(\col[0].zbuf_bot_iw_I[2].a ),
    .X(net491));
 sky130_fd_sc_hd__clkbuf_4 fanout492 (.A(\col[0].zbuf_bot_iw_I[2].a ),
    .X(net492));
 sky130_fd_sc_hd__buf_6 fanout493 (.A(\col[0].zbuf_bot_iw_I[1].a ),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_4 fanout494 (.A(\col[0].zbuf_bot_iw_I[1].a ),
    .X(net494));
 sky130_fd_sc_hd__buf_6 fanout495 (.A(\col[0].zbuf_bot_iw_I[17].a ),
    .X(net495));
 sky130_fd_sc_hd__clkbuf_4 fanout496 (.A(\col[0].zbuf_bot_iw_I[17].a ),
    .X(net496));
 sky130_fd_sc_hd__buf_6 fanout497 (.A(\col[0].zbuf_bot_iw_I[16].a ),
    .X(net497));
 sky130_fd_sc_hd__clkbuf_4 fanout498 (.A(\col[0].zbuf_bot_iw_I[16].a ),
    .X(net498));
 sky130_fd_sc_hd__buf_6 fanout499 (.A(\col[0].zbuf_bot_iw_I[15].a ),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_4 fanout500 (.A(\col[0].zbuf_bot_iw_I[15].a ),
    .X(net500));
 sky130_fd_sc_hd__buf_6 fanout501 (.A(\col[0].zbuf_bot_iw_I[14].a ),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_4 fanout502 (.A(\col[0].zbuf_bot_iw_I[14].a ),
    .X(net502));
 sky130_fd_sc_hd__buf_6 fanout503 (.A(\col[0].zbuf_bot_iw_I[13].a ),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_4 fanout504 (.A(\col[0].zbuf_bot_iw_I[13].a ),
    .X(net504));
 sky130_fd_sc_hd__buf_6 fanout505 (.A(\col[0].zbuf_bot_iw_I[12].a ),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_4 fanout506 (.A(\col[0].zbuf_bot_iw_I[12].a ),
    .X(net506));
 sky130_fd_sc_hd__buf_6 fanout507 (.A(\col[0].zbuf_bot_iw_I[11].a ),
    .X(net507));
 sky130_fd_sc_hd__clkbuf_4 fanout508 (.A(\col[0].zbuf_bot_iw_I[11].a ),
    .X(net508));
 sky130_fd_sc_hd__buf_8 fanout509 (.A(\col[0].zbuf_bot_iw_I[10].a ),
    .X(net509));
 sky130_fd_sc_hd__clkbuf_4 fanout510 (.A(\col[0].zbuf_bot_iw_I[10].a ),
    .X(net510));
 sky130_fd_sc_hd__buf_6 fanout511 (.A(\col[0].zbuf_bot_iw_I[0].a ),
    .X(net511));
 sky130_fd_sc_hd__clkbuf_4 fanout512 (.A(\col[0].zbuf_bot_iw_I[0].a ),
    .X(net512));
 sky130_fd_sc_hd__clkbuf_2 fanout513 (.A(net514),
    .X(net513));
 sky130_fd_sc_hd__clkbuf_1 fanout514 (.A(net515),
    .X(net514));
 sky130_fd_sc_hd__clkbuf_1 fanout515 (.A(net516),
    .X(net515));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout516 (.A(\zbuf_bus_ena_I.e ),
    .X(net516));
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(addr[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(spine_iw[14]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(um_ow[159]),
    .X(net100));
 sky130_fd_sc_hd__dlymetal6s2s_1 input101 (.A(um_ow[15]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(um_ow[160]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 input103 (.A(um_ow[161]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 input104 (.A(um_ow[162]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(um_ow[163]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(um_ow[164]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 input107 (.A(um_ow[165]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 input108 (.A(um_ow[166]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 input109 (.A(um_ow[167]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(spine_iw[15]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input110 (.A(um_ow[168]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 input111 (.A(um_ow[169]),
    .X(net111));
 sky130_fd_sc_hd__dlymetal6s2s_1 input112 (.A(um_ow[16]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 input113 (.A(um_ow[170]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 input114 (.A(um_ow[171]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 input115 (.A(um_ow[172]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 input116 (.A(um_ow[173]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 input117 (.A(um_ow[174]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 input118 (.A(um_ow[175]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 input119 (.A(um_ow[176]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(spine_iw[16]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input120 (.A(um_ow[177]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 input121 (.A(um_ow[178]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(um_ow[179]),
    .X(net122));
 sky130_fd_sc_hd__dlymetal6s2s_1 input123 (.A(um_ow[17]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(um_ow[180]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 input125 (.A(um_ow[181]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(um_ow[182]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(um_ow[183]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 input128 (.A(um_ow[184]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 input129 (.A(um_ow[185]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(spine_iw[17]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input130 (.A(um_ow[186]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 input131 (.A(um_ow[187]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(um_ow[188]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 input133 (.A(um_ow[189]),
    .X(net133));
 sky130_fd_sc_hd__dlymetal6s2s_1 input134 (.A(um_ow[18]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 input135 (.A(um_ow[190]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 input136 (.A(um_ow[191]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 input137 (.A(um_ow[192]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 input138 (.A(um_ow[193]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 input139 (.A(um_ow[194]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(spine_iw[18]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input140 (.A(um_ow[195]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 input141 (.A(um_ow[196]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 input142 (.A(um_ow[197]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 input143 (.A(um_ow[198]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 input144 (.A(um_ow[199]),
    .X(net144));
 sky130_fd_sc_hd__dlymetal6s2s_1 input145 (.A(um_ow[19]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 input146 (.A(um_ow[1]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 input147 (.A(um_ow[200]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 input148 (.A(um_ow[201]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 input149 (.A(um_ow[202]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(spine_iw[19]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input150 (.A(um_ow[203]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 input151 (.A(um_ow[204]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 input152 (.A(um_ow[205]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 input153 (.A(um_ow[206]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 input154 (.A(um_ow[207]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 input155 (.A(um_ow[208]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_1 input156 (.A(um_ow[209]),
    .X(net156));
 sky130_fd_sc_hd__dlymetal6s2s_1 input157 (.A(um_ow[20]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 input158 (.A(um_ow[210]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 input159 (.A(um_ow[211]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(spine_iw[1]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input160 (.A(um_ow[212]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 input161 (.A(um_ow[213]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 input162 (.A(um_ow[214]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 input163 (.A(um_ow[215]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 input164 (.A(um_ow[216]),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 input165 (.A(um_ow[217]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 input166 (.A(um_ow[218]),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 input167 (.A(um_ow[219]),
    .X(net167));
 sky130_fd_sc_hd__dlymetal6s2s_1 input168 (.A(um_ow[21]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 input169 (.A(um_ow[220]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(spine_iw[20]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input170 (.A(um_ow[221]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 input171 (.A(um_ow[222]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 input172 (.A(um_ow[223]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 input173 (.A(um_ow[224]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 input174 (.A(um_ow[225]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(um_ow[226]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(um_ow[227]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 input177 (.A(um_ow[228]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 input178 (.A(um_ow[229]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_2 input179 (.A(um_ow[22]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(spine_iw[21]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input180 (.A(um_ow[230]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_1 input181 (.A(um_ow[231]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 input182 (.A(um_ow[232]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 input183 (.A(um_ow[233]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 input184 (.A(um_ow[234]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 input185 (.A(um_ow[235]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 input186 (.A(um_ow[236]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 input187 (.A(um_ow[237]),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 input188 (.A(um_ow[238]),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 input189 (.A(um_ow[239]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(spine_iw[22]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input190 (.A(um_ow[23]),
    .X(net190));
 sky130_fd_sc_hd__dlymetal6s2s_1 input191 (.A(um_ow[240]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 input192 (.A(um_ow[241]),
    .X(net192));
 sky130_fd_sc_hd__dlymetal6s2s_1 input193 (.A(um_ow[242]),
    .X(net193));
 sky130_fd_sc_hd__dlymetal6s2s_1 input194 (.A(um_ow[243]),
    .X(net194));
 sky130_fd_sc_hd__dlymetal6s2s_1 input195 (.A(um_ow[244]),
    .X(net195));
 sky130_fd_sc_hd__dlymetal6s2s_1 input196 (.A(um_ow[245]),
    .X(net196));
 sky130_fd_sc_hd__dlymetal6s2s_1 input197 (.A(um_ow[246]),
    .X(net197));
 sky130_fd_sc_hd__dlymetal6s2s_1 input198 (.A(um_ow[247]),
    .X(net198));
 sky130_fd_sc_hd__dlymetal6s2s_1 input199 (.A(um_ow[248]),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(addr[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(spine_iw[23]),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 input200 (.A(um_ow[249]),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_2 input201 (.A(um_ow[24]),
    .X(net201));
 sky130_fd_sc_hd__dlymetal6s2s_1 input202 (.A(um_ow[250]),
    .X(net202));
 sky130_fd_sc_hd__dlymetal6s2s_1 input203 (.A(um_ow[251]),
    .X(net203));
 sky130_fd_sc_hd__dlymetal6s2s_1 input204 (.A(um_ow[252]),
    .X(net204));
 sky130_fd_sc_hd__dlymetal6s2s_1 input205 (.A(um_ow[253]),
    .X(net205));
 sky130_fd_sc_hd__dlymetal6s2s_1 input206 (.A(um_ow[254]),
    .X(net206));
 sky130_fd_sc_hd__dlymetal6s2s_1 input207 (.A(um_ow[255]),
    .X(net207));
 sky130_fd_sc_hd__dlymetal6s2s_1 input208 (.A(um_ow[256]),
    .X(net208));
 sky130_fd_sc_hd__dlymetal6s2s_1 input209 (.A(um_ow[257]),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(spine_iw[24]),
    .X(net21));
 sky130_fd_sc_hd__dlymetal6s2s_1 input210 (.A(um_ow[258]),
    .X(net210));
 sky130_fd_sc_hd__dlymetal6s2s_1 input211 (.A(um_ow[259]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_2 input212 (.A(um_ow[25]),
    .X(net212));
 sky130_fd_sc_hd__dlymetal6s2s_1 input213 (.A(um_ow[260]),
    .X(net213));
 sky130_fd_sc_hd__dlymetal6s2s_1 input214 (.A(um_ow[261]),
    .X(net214));
 sky130_fd_sc_hd__dlymetal6s2s_1 input215 (.A(um_ow[262]),
    .X(net215));
 sky130_fd_sc_hd__dlymetal6s2s_1 input216 (.A(um_ow[263]),
    .X(net216));
 sky130_fd_sc_hd__dlymetal6s2s_1 input217 (.A(um_ow[264]),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_1 input218 (.A(um_ow[265]),
    .X(net218));
 sky130_fd_sc_hd__dlymetal6s2s_1 input219 (.A(um_ow[266]),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(spine_iw[25]),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input220 (.A(um_ow[267]),
    .X(net220));
 sky130_fd_sc_hd__dlymetal6s2s_1 input221 (.A(um_ow[268]),
    .X(net221));
 sky130_fd_sc_hd__dlymetal6s2s_1 input222 (.A(um_ow[269]),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_2 input223 (.A(um_ow[26]),
    .X(net223));
 sky130_fd_sc_hd__dlymetal6s2s_1 input224 (.A(um_ow[270]),
    .X(net224));
 sky130_fd_sc_hd__dlymetal6s2s_1 input225 (.A(um_ow[271]),
    .X(net225));
 sky130_fd_sc_hd__dlymetal6s2s_1 input226 (.A(um_ow[272]),
    .X(net226));
 sky130_fd_sc_hd__dlymetal6s2s_1 input227 (.A(um_ow[273]),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_2 input228 (.A(um_ow[274]),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_2 input229 (.A(um_ow[275]),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(spine_iw[26]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input230 (.A(um_ow[276]),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_2 input231 (.A(um_ow[277]),
    .X(net231));
 sky130_fd_sc_hd__dlymetal6s2s_1 input232 (.A(um_ow[278]),
    .X(net232));
 sky130_fd_sc_hd__dlymetal6s2s_1 input233 (.A(um_ow[279]),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_2 input234 (.A(um_ow[27]),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_2 input235 (.A(um_ow[280]),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_2 input236 (.A(um_ow[281]),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_2 input237 (.A(um_ow[282]),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_2 input238 (.A(um_ow[283]),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_2 input239 (.A(um_ow[284]),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(spine_iw[27]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input240 (.A(um_ow[285]),
    .X(net240));
 sky130_fd_sc_hd__dlymetal6s2s_1 input241 (.A(um_ow[286]),
    .X(net241));
 sky130_fd_sc_hd__dlymetal6s2s_1 input242 (.A(um_ow[287]),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_1 input243 (.A(um_ow[288]),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_1 input244 (.A(um_ow[289]),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_2 input245 (.A(um_ow[28]),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_1 input246 (.A(um_ow[290]),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_1 input247 (.A(um_ow[291]),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_1 input248 (.A(um_ow[292]),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_1 input249 (.A(um_ow[293]),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(spine_iw[28]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input250 (.A(um_ow[294]),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_1 input251 (.A(um_ow[295]),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 input252 (.A(um_ow[296]),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_1 input253 (.A(um_ow[297]),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_1 input254 (.A(um_ow[298]),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_1 input255 (.A(um_ow[299]),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_2 input256 (.A(um_ow[29]),
    .X(net256));
 sky130_fd_sc_hd__dlymetal6s2s_1 input257 (.A(um_ow[2]),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_1 input258 (.A(um_ow[300]),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_1 input259 (.A(um_ow[301]),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(spine_iw[29]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input260 (.A(um_ow[302]),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_1 input261 (.A(um_ow[303]),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_1 input262 (.A(um_ow[304]),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_1 input263 (.A(um_ow[305]),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_1 input264 (.A(um_ow[306]),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_1 input265 (.A(um_ow[307]),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_1 input266 (.A(um_ow[308]),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_1 input267 (.A(um_ow[309]),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_2 input268 (.A(um_ow[30]),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_1 input269 (.A(um_ow[310]),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(spine_iw[2]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input270 (.A(um_ow[311]),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_1 input271 (.A(um_ow[312]),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_1 input272 (.A(um_ow[313]),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_1 input273 (.A(um_ow[314]),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_1 input274 (.A(um_ow[315]),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_1 input275 (.A(um_ow[316]),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_1 input276 (.A(um_ow[317]),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_1 input277 (.A(um_ow[318]),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_1 input278 (.A(um_ow[319]),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_2 input279 (.A(um_ow[31]),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(spine_iw[3]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input280 (.A(um_ow[320]),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_1 input281 (.A(um_ow[321]),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_1 input282 (.A(um_ow[322]),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_1 input283 (.A(um_ow[323]),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_1 input284 (.A(um_ow[324]),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_1 input285 (.A(um_ow[325]),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_1 input286 (.A(um_ow[326]),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_1 input287 (.A(um_ow[327]),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_1 input288 (.A(um_ow[328]),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_1 input289 (.A(um_ow[329]),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(spine_iw[4]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input290 (.A(um_ow[32]),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_1 input291 (.A(um_ow[330]),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_1 input292 (.A(um_ow[331]),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_1 input293 (.A(um_ow[332]),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_1 input294 (.A(um_ow[333]),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_1 input295 (.A(um_ow[334]),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_1 input296 (.A(um_ow[335]),
    .X(net296));
 sky130_fd_sc_hd__dlymetal6s2s_1 input297 (.A(um_ow[336]),
    .X(net297));
 sky130_fd_sc_hd__dlymetal6s2s_1 input298 (.A(um_ow[337]),
    .X(net298));
 sky130_fd_sc_hd__dlymetal6s2s_1 input299 (.A(um_ow[338]),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(addr[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(spine_iw[5]),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 input300 (.A(um_ow[339]),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_2 input301 (.A(um_ow[33]),
    .X(net301));
 sky130_fd_sc_hd__dlymetal6s2s_1 input302 (.A(um_ow[340]),
    .X(net302));
 sky130_fd_sc_hd__dlymetal6s2s_1 input303 (.A(um_ow[341]),
    .X(net303));
 sky130_fd_sc_hd__dlymetal6s2s_1 input304 (.A(um_ow[342]),
    .X(net304));
 sky130_fd_sc_hd__dlymetal6s2s_1 input305 (.A(um_ow[343]),
    .X(net305));
 sky130_fd_sc_hd__dlymetal6s2s_1 input306 (.A(um_ow[344]),
    .X(net306));
 sky130_fd_sc_hd__dlymetal6s2s_1 input307 (.A(um_ow[345]),
    .X(net307));
 sky130_fd_sc_hd__dlymetal6s2s_1 input308 (.A(um_ow[346]),
    .X(net308));
 sky130_fd_sc_hd__dlymetal6s2s_1 input309 (.A(um_ow[347]),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(spine_iw[6]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input310 (.A(um_ow[348]),
    .X(net310));
 sky130_fd_sc_hd__dlymetal6s2s_1 input311 (.A(um_ow[349]),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_2 input312 (.A(um_ow[34]),
    .X(net312));
 sky130_fd_sc_hd__dlymetal6s2s_1 input313 (.A(um_ow[350]),
    .X(net313));
 sky130_fd_sc_hd__dlymetal6s2s_1 input314 (.A(um_ow[351]),
    .X(net314));
 sky130_fd_sc_hd__dlymetal6s2s_1 input315 (.A(um_ow[352]),
    .X(net315));
 sky130_fd_sc_hd__dlymetal6s2s_1 input316 (.A(um_ow[353]),
    .X(net316));
 sky130_fd_sc_hd__dlymetal6s2s_1 input317 (.A(um_ow[354]),
    .X(net317));
 sky130_fd_sc_hd__dlymetal6s2s_1 input318 (.A(um_ow[355]),
    .X(net318));
 sky130_fd_sc_hd__dlymetal6s2s_1 input319 (.A(um_ow[356]),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(spine_iw[7]),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 input320 (.A(um_ow[357]),
    .X(net320));
 sky130_fd_sc_hd__dlymetal6s2s_1 input321 (.A(um_ow[358]),
    .X(net321));
 sky130_fd_sc_hd__dlymetal6s2s_1 input322 (.A(um_ow[359]),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_2 input323 (.A(um_ow[35]),
    .X(net323));
 sky130_fd_sc_hd__dlymetal6s2s_1 input324 (.A(um_ow[360]),
    .X(net324));
 sky130_fd_sc_hd__dlymetal6s2s_1 input325 (.A(um_ow[361]),
    .X(net325));
 sky130_fd_sc_hd__dlymetal6s2s_1 input326 (.A(um_ow[362]),
    .X(net326));
 sky130_fd_sc_hd__dlymetal6s2s_1 input327 (.A(um_ow[363]),
    .X(net327));
 sky130_fd_sc_hd__dlymetal6s2s_1 input328 (.A(um_ow[364]),
    .X(net328));
 sky130_fd_sc_hd__dlymetal6s2s_1 input329 (.A(um_ow[365]),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(spine_iw[8]),
    .X(net33));
 sky130_fd_sc_hd__dlymetal6s2s_1 input330 (.A(um_ow[366]),
    .X(net330));
 sky130_fd_sc_hd__dlymetal6s2s_1 input331 (.A(um_ow[367]),
    .X(net331));
 sky130_fd_sc_hd__dlymetal6s2s_1 input332 (.A(um_ow[368]),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_2 input333 (.A(um_ow[369]),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_2 input334 (.A(um_ow[36]),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_2 input335 (.A(um_ow[370]),
    .X(net335));
 sky130_fd_sc_hd__dlymetal6s2s_1 input336 (.A(um_ow[371]),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_2 input337 (.A(um_ow[372]),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_2 input338 (.A(um_ow[373]),
    .X(net338));
 sky130_fd_sc_hd__dlymetal6s2s_1 input339 (.A(um_ow[374]),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(spine_iw[9]),
    .X(net34));
 sky130_fd_sc_hd__dlymetal6s2s_1 input340 (.A(um_ow[375]),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_2 input341 (.A(um_ow[376]),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_2 input342 (.A(um_ow[377]),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_2 input343 (.A(um_ow[378]),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_2 input344 (.A(um_ow[379]),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_2 input345 (.A(um_ow[37]),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_2 input346 (.A(um_ow[380]),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_2 input347 (.A(um_ow[381]),
    .X(net347));
 sky130_fd_sc_hd__dlymetal6s2s_1 input348 (.A(um_ow[382]),
    .X(net348));
 sky130_fd_sc_hd__dlymetal6s2s_1 input349 (.A(um_ow[383]),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(um_ow[0]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input350 (.A(um_ow[38]),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_2 input351 (.A(um_ow[39]),
    .X(net351));
 sky130_fd_sc_hd__dlymetal6s2s_1 input352 (.A(um_ow[3]),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_2 input353 (.A(um_ow[40]),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_2 input354 (.A(um_ow[41]),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_2 input355 (.A(um_ow[42]),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_2 input356 (.A(um_ow[43]),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_2 input357 (.A(um_ow[44]),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_2 input358 (.A(um_ow[45]),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_2 input359 (.A(um_ow[46]),
    .X(net359));
 sky130_fd_sc_hd__dlymetal6s2s_1 input36 (.A(um_ow[100]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input360 (.A(um_ow[47]),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_1 input361 (.A(um_ow[48]),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_1 input362 (.A(um_ow[49]),
    .X(net362));
 sky130_fd_sc_hd__dlymetal6s2s_1 input363 (.A(um_ow[4]),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_1 input364 (.A(um_ow[50]),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_1 input365 (.A(um_ow[51]),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_1 input366 (.A(um_ow[52]),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_1 input367 (.A(um_ow[53]),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_1 input368 (.A(um_ow[54]),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_1 input369 (.A(um_ow[55]),
    .X(net369));
 sky130_fd_sc_hd__dlymetal6s2s_1 input37 (.A(um_ow[101]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input370 (.A(um_ow[56]),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_1 input371 (.A(um_ow[57]),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_1 input372 (.A(um_ow[58]),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_1 input373 (.A(um_ow[59]),
    .X(net373));
 sky130_fd_sc_hd__dlymetal6s2s_1 input374 (.A(um_ow[5]),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_1 input375 (.A(um_ow[60]),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_1 input376 (.A(um_ow[61]),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_1 input377 (.A(um_ow[62]),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_1 input378 (.A(um_ow[63]),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_1 input379 (.A(um_ow[64]),
    .X(net379));
 sky130_fd_sc_hd__dlymetal6s2s_1 input38 (.A(um_ow[102]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input380 (.A(um_ow[65]),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_1 input381 (.A(um_ow[66]),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_1 input382 (.A(um_ow[67]),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_1 input383 (.A(um_ow[68]),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_1 input384 (.A(um_ow[69]),
    .X(net384));
 sky130_fd_sc_hd__dlymetal6s2s_1 input385 (.A(um_ow[6]),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_1 input386 (.A(um_ow[70]),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_1 input387 (.A(um_ow[71]),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_1 input388 (.A(um_ow[72]),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_1 input389 (.A(um_ow[73]),
    .X(net389));
 sky130_fd_sc_hd__dlymetal6s2s_1 input39 (.A(um_ow[103]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input390 (.A(um_ow[74]),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_1 input391 (.A(um_ow[75]),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_1 input392 (.A(um_ow[76]),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_1 input393 (.A(um_ow[77]),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_1 input394 (.A(um_ow[78]),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_1 input395 (.A(um_ow[79]),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_2 input396 (.A(um_ow[7]),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_1 input397 (.A(um_ow[80]),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_1 input398 (.A(um_ow[81]),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_1 input399 (.A(um_ow[82]),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(addr[3]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input40 (.A(um_ow[104]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input400 (.A(um_ow[83]),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_1 input401 (.A(um_ow[84]),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_1 input402 (.A(um_ow[85]),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_1 input403 (.A(um_ow[86]),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_1 input404 (.A(um_ow[87]),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_1 input405 (.A(um_ow[88]),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_1 input406 (.A(um_ow[89]),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_2 input407 (.A(um_ow[8]),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_1 input408 (.A(um_ow[90]),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_1 input409 (.A(um_ow[91]),
    .X(net409));
 sky130_fd_sc_hd__dlymetal6s2s_1 input41 (.A(um_ow[105]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input410 (.A(um_ow[92]),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_1 input411 (.A(um_ow[93]),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_1 input412 (.A(um_ow[94]),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_1 input413 (.A(um_ow[95]),
    .X(net413));
 sky130_fd_sc_hd__dlymetal6s2s_1 input414 (.A(um_ow[96]),
    .X(net414));
 sky130_fd_sc_hd__dlymetal6s2s_1 input415 (.A(um_ow[97]),
    .X(net415));
 sky130_fd_sc_hd__dlymetal6s2s_1 input416 (.A(um_ow[98]),
    .X(net416));
 sky130_fd_sc_hd__dlymetal6s2s_1 input417 (.A(um_ow[99]),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_2 input418 (.A(um_ow[9]),
    .X(net418));
 sky130_fd_sc_hd__dlymetal6s2s_1 input42 (.A(um_ow[106]),
    .X(net42));
 sky130_fd_sc_hd__dlymetal6s2s_1 input43 (.A(um_ow[107]),
    .X(net43));
 sky130_fd_sc_hd__dlymetal6s2s_1 input44 (.A(um_ow[108]),
    .X(net44));
 sky130_fd_sc_hd__dlymetal6s2s_1 input45 (.A(um_ow[109]),
    .X(net45));
 sky130_fd_sc_hd__dlymetal6s2s_1 input46 (.A(um_ow[10]),
    .X(net46));
 sky130_fd_sc_hd__dlymetal6s2s_1 input47 (.A(um_ow[110]),
    .X(net47));
 sky130_fd_sc_hd__dlymetal6s2s_1 input48 (.A(um_ow[111]),
    .X(net48));
 sky130_fd_sc_hd__dlymetal6s2s_1 input49 (.A(um_ow[112]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(addr[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(um_ow[113]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(um_ow[114]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(um_ow[115]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(um_ow[116]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(um_ow[117]),
    .X(net54));
 sky130_fd_sc_hd__dlymetal6s2s_1 input55 (.A(um_ow[118]),
    .X(net55));
 sky130_fd_sc_hd__dlymetal6s2s_1 input56 (.A(um_ow[119]),
    .X(net56));
 sky130_fd_sc_hd__dlymetal6s2s_1 input57 (.A(um_ow[11]),
    .X(net57));
 sky130_fd_sc_hd__dlymetal6s2s_1 input58 (.A(um_ow[120]),
    .X(net58));
 sky130_fd_sc_hd__dlymetal6s2s_1 input59 (.A(um_ow[121]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(spine_iw[10]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(um_ow[122]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(um_ow[123]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(um_ow[124]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 input63 (.A(um_ow[125]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 input64 (.A(um_ow[126]),
    .X(net64));
 sky130_fd_sc_hd__dlymetal6s2s_1 input65 (.A(um_ow[127]),
    .X(net65));
 sky130_fd_sc_hd__dlymetal6s2s_1 input66 (.A(um_ow[128]),
    .X(net66));
 sky130_fd_sc_hd__dlymetal6s2s_1 input67 (.A(um_ow[129]),
    .X(net67));
 sky130_fd_sc_hd__dlymetal6s2s_1 input68 (.A(um_ow[12]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 input69 (.A(um_ow[130]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(spine_iw[11]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input70 (.A(um_ow[131]),
    .X(net70));
 sky130_fd_sc_hd__dlymetal6s2s_1 input71 (.A(um_ow[132]),
    .X(net71));
 sky130_fd_sc_hd__dlymetal6s2s_1 input72 (.A(um_ow[133]),
    .X(net72));
 sky130_fd_sc_hd__dlymetal6s2s_1 input73 (.A(um_ow[134]),
    .X(net73));
 sky130_fd_sc_hd__dlymetal6s2s_1 input74 (.A(um_ow[135]),
    .X(net74));
 sky130_fd_sc_hd__dlymetal6s2s_1 input75 (.A(um_ow[136]),
    .X(net75));
 sky130_fd_sc_hd__dlymetal6s2s_1 input76 (.A(um_ow[137]),
    .X(net76));
 sky130_fd_sc_hd__dlymetal6s2s_1 input77 (.A(um_ow[138]),
    .X(net77));
 sky130_fd_sc_hd__dlymetal6s2s_1 input78 (.A(um_ow[139]),
    .X(net78));
 sky130_fd_sc_hd__dlymetal6s2s_1 input79 (.A(um_ow[13]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(spine_iw[12]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input80 (.A(um_ow[140]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(um_ow[141]),
    .X(net81));
 sky130_fd_sc_hd__dlymetal6s2s_1 input82 (.A(um_ow[142]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(um_ow[143]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(um_ow[144]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(um_ow[145]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(um_ow[146]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(um_ow[147]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(um_ow[148]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(um_ow[149]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(spine_iw[13]),
    .X(net9));
 sky130_fd_sc_hd__dlymetal6s2s_1 input90 (.A(um_ow[14]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(um_ow[150]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(um_ow[151]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(um_ow[152]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(um_ow[153]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(um_ow[154]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(um_ow[155]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(um_ow[156]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 input98 (.A(um_ow[157]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 input99 (.A(um_ow[158]),
    .X(net99));
 sky130_fd_sc_hd__conb_1 tt_mux_517 (.LO(net517));
 sky130_fd_sc_hd__conb_1 tt_mux_518 (.LO(net518));
 sky130_fd_sc_hd__conb_1 tt_mux_519 (.LO(net519));
 sky130_fd_sc_hd__conb_1 tt_mux_520 (.LO(net520));
 sky130_fd_sc_hd__conb_1 tt_mux_521 (.LO(net521));
 sky130_fd_sc_hd__conb_1 tt_mux_522 (.LO(net522));
 sky130_fd_sc_hd__conb_1 tt_mux_523 (.LO(net523));
 sky130_fd_sc_hd__conb_1 tt_mux_524 (.LO(net524));
 sky130_fd_sc_hd__conb_1 tt_mux_525 (.LO(net525));
 sky130_fd_sc_hd__conb_1 tt_mux_526 (.LO(net526));
 sky130_fd_sc_hd__conb_1 tt_mux_527 (.LO(net527));
 sky130_fd_sc_hd__conb_1 tt_mux_528 (.LO(net528));
 sky130_fd_sc_hd__conb_1 tt_mux_529 (.LO(net529));
 sky130_fd_sc_hd__conb_1 tt_mux_530 (.LO(net530));
 sky130_fd_sc_hd__conb_1 tt_mux_531 (.LO(net531));
 sky130_fd_sc_hd__conb_1 tt_mux_532 (.LO(net532));
 sky130_fd_sc_hd__conb_1 tt_mux_533 (.LO(net533));
 sky130_fd_sc_hd__conb_1 tt_mux_534 (.LO(net534));
 sky130_fd_sc_hd__conb_1 tt_mux_535 (.LO(net535));
 sky130_fd_sc_hd__conb_1 tt_mux_552 (.HI(net552));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_ena_I.genblk1.cell0_I  (.A(net16),
    .B(net516),
    .X(\zbuf_bus_ena_I.genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_ena_I.genblk1.cell1_I  (.A(\zbuf_bus_ena_I.genblk1.l ),
    .X(\zbuf_bus_ena_I.z ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[0].genblk1.cell0_I  (.A(net8),
    .B(net513),
    .X(\zbuf_bus_iw_I[0].genblk1.l ));
 sky130_fd_sc_hd__buf_6 \zbuf_bus_iw_I[0].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[0].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[0].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[10].genblk1.cell0_I  (.A(net19),
    .B(net515),
    .X(\zbuf_bus_iw_I[10].genblk1.l ));
 sky130_fd_sc_hd__buf_6 \zbuf_bus_iw_I[10].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[10].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[10].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[11].genblk1.cell0_I  (.A(net20),
    .B(net515),
    .X(\zbuf_bus_iw_I[11].genblk1.l ));
 sky130_fd_sc_hd__buf_6 \zbuf_bus_iw_I[11].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[11].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[11].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[12].genblk1.cell0_I  (.A(net21),
    .B(net515),
    .X(\zbuf_bus_iw_I[12].genblk1.l ));
 sky130_fd_sc_hd__buf_6 \zbuf_bus_iw_I[12].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[12].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[12].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[13].genblk1.cell0_I  (.A(net22),
    .B(net515),
    .X(\zbuf_bus_iw_I[13].genblk1.l ));
 sky130_fd_sc_hd__buf_6 \zbuf_bus_iw_I[13].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[13].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[13].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[14].genblk1.cell0_I  (.A(net23),
    .B(net513),
    .X(\zbuf_bus_iw_I[14].genblk1.l ));
 sky130_fd_sc_hd__buf_6 \zbuf_bus_iw_I[14].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[14].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[14].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[15].genblk1.cell0_I  (.A(net24),
    .B(net513),
    .X(\zbuf_bus_iw_I[15].genblk1.l ));
 sky130_fd_sc_hd__buf_6 \zbuf_bus_iw_I[15].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[15].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[15].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[16].genblk1.cell0_I  (.A(net25),
    .B(net513),
    .X(\zbuf_bus_iw_I[16].genblk1.l ));
 sky130_fd_sc_hd__buf_6 \zbuf_bus_iw_I[16].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[16].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[16].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[17].genblk1.cell0_I  (.A(net26),
    .B(net513),
    .X(\zbuf_bus_iw_I[17].genblk1.l ));
 sky130_fd_sc_hd__buf_6 \zbuf_bus_iw_I[17].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[17].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[17].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[1].genblk1.cell0_I  (.A(net9),
    .B(net513),
    .X(\zbuf_bus_iw_I[1].genblk1.l ));
 sky130_fd_sc_hd__buf_6 \zbuf_bus_iw_I[1].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[1].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[1].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[2].genblk1.cell0_I  (.A(net10),
    .B(net513),
    .X(\zbuf_bus_iw_I[2].genblk1.l ));
 sky130_fd_sc_hd__buf_6 \zbuf_bus_iw_I[2].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[2].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[2].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[3].genblk1.cell0_I  (.A(net11),
    .B(net513),
    .X(\zbuf_bus_iw_I[3].genblk1.l ));
 sky130_fd_sc_hd__buf_6 \zbuf_bus_iw_I[3].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[3].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[3].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[4].genblk1.cell0_I  (.A(net12),
    .B(net514),
    .X(\zbuf_bus_iw_I[4].genblk1.l ));
 sky130_fd_sc_hd__buf_6 \zbuf_bus_iw_I[4].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[4].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[4].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[5].genblk1.cell0_I  (.A(net13),
    .B(net514),
    .X(\zbuf_bus_iw_I[5].genblk1.l ));
 sky130_fd_sc_hd__buf_6 \zbuf_bus_iw_I[5].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[5].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[5].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[6].genblk1.cell0_I  (.A(net14),
    .B(net514),
    .X(\zbuf_bus_iw_I[6].genblk1.l ));
 sky130_fd_sc_hd__buf_6 \zbuf_bus_iw_I[6].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[6].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[6].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[7].genblk1.cell0_I  (.A(net15),
    .B(net513),
    .X(\zbuf_bus_iw_I[7].genblk1.l ));
 sky130_fd_sc_hd__buf_6 \zbuf_bus_iw_I[7].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[7].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[7].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[8].genblk1.cell0_I  (.A(net17),
    .B(net513),
    .X(\zbuf_bus_iw_I[8].genblk1.l ));
 sky130_fd_sc_hd__buf_6 \zbuf_bus_iw_I[8].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[8].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[8].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_iw_I[9].genblk1.cell0_I  (.A(net18),
    .B(net514),
    .X(\zbuf_bus_iw_I[9].genblk1.l ));
 sky130_fd_sc_hd__buf_6 \zbuf_bus_iw_I[9].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[9].genblk1.l ),
    .X(\col[0].zbuf_bot_iw_I[9].a ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_sel_I[0].genblk1.cell0_I  (.A(net32),
    .B(net516),
    .X(\zbuf_bus_sel_I[0].genblk1.l ));
 sky130_fd_sc_hd__buf_6 \zbuf_bus_sel_I[0].genblk1.cell1_I  (.A(\zbuf_bus_sel_I[0].genblk1.l ),
    .X(\zbuf_bus_sel_I[0].z ));
 sky130_fd_sc_hd__and2_1 \zbuf_bus_sel_I[1].genblk1.cell0_I  (.A(net27),
    .B(net516),
    .X(\zbuf_bus_sel_I[1].genblk1.l ));
 sky130_fd_sc_hd__clkbuf_1 \zbuf_bus_sel_I[1].genblk1.cell1_I  (.A(\zbuf_bus_sel_I[1].genblk1.l ),
    .X(\zbuf_bus_sel_I[1].z ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_sel_I[2].genblk1.cell0_I  (.A(net28),
    .B(net516),
    .X(\zbuf_bus_sel_I[2].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_sel_I[2].genblk1.cell1_I  (.A(\zbuf_bus_sel_I[2].genblk1.l ),
    .X(\zbuf_bus_sel_I[2].z ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_sel_I[3].genblk1.cell0_I  (.A(net29),
    .B(net516),
    .X(\zbuf_bus_sel_I[3].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_sel_I[3].genblk1.cell1_I  (.A(\zbuf_bus_sel_I[3].genblk1.l ),
    .X(\zbuf_bus_sel_I[3].z ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_sel_I[4].genblk1.cell0_I  (.A(net30),
    .B(net516),
    .X(\zbuf_bus_sel_I[4].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_sel_I[4].genblk1.cell1_I  (.A(\zbuf_bus_sel_I[4].genblk1.l ),
    .X(\zbuf_bus_sel_I[4].z ));
 assign k_one = net552;
 assign k_zero = net517;
 assign spine_ow[0] = net518;
 assign spine_ow[25] = net519;
 assign um_k_zero[0] = net520;
 assign um_k_zero[10] = net530;
 assign um_k_zero[11] = net531;
 assign um_k_zero[12] = net532;
 assign um_k_zero[13] = net533;
 assign um_k_zero[14] = net534;
 assign um_k_zero[15] = net535;
 assign um_k_zero[1] = net521;
 assign um_k_zero[2] = net522;
 assign um_k_zero[3] = net523;
 assign um_k_zero[4] = net524;
 assign um_k_zero[5] = net525;
 assign um_k_zero[6] = net526;
 assign um_k_zero[7] = net527;
 assign um_k_zero[8] = net528;
 assign um_k_zero[9] = net529;
endmodule

