// This is the unpowered netlist.
module user_project_wrapper (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire \tt_top1.io_oeb[0] ;
 wire \tt_top1.io_oeb[16] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.clk ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ena ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.k_zero ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[0].um_bot_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.clk ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ena ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.k_zero ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[0].um_top_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.clk ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ena ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.k_zero ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[1].um_bot_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.clk ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ena ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.k_zero ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[1].um_top_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.clk ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ena ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.k_zero ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[2].um_bot_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.clk ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ena ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.k_zero ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[2].um_top_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.clk ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.ena ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.clk ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ena ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.k_zero ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[3].um_top_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.clk ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ena ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.k_zero ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[4].um_bot_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.clk ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ena ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.k_zero ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[4].um_top_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.clk ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.ena ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.clk ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ena ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.k_zero ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[5].um_top_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.clk ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.ena ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.clk ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ena ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.k_zero ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[6].um_top_I.ow[9] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.clk ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.ena ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.clk ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ena ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[10] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[11] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[12] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[13] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[14] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[15] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[16] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[17] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[1] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[2] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[3] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[4] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[5] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[6] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[7] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[8] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.iw[9] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.k_zero ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[0] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[10] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[11] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[12] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[13] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[14] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[15] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[16] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[17] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[18] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[19] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[1] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[20] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[21] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[22] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[23] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[2] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[3] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[4] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[5] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[6] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[7] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[8] ;
 wire \tt_top1.branch[0].col_um[7].um_top_I.ow[9] ;
 wire \tt_top1.branch[0].l_addr[0] ;
 wire \tt_top1.branch[0].l_k_one ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.clk ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ena ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.k_zero ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[0].um_bot_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.clk ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ena ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.k_zero ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[0].um_top_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.clk ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ena ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.k_zero ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[1].um_bot_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.clk ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ena ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.k_zero ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[1].um_top_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.clk ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ena ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.k_zero ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[2].um_bot_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.clk ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ena ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.k_zero ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[2].um_top_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.clk ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ena ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.k_zero ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[3].um_bot_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.clk ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ena ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.k_zero ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[3].um_top_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.clk ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ena ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.k_zero ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[4].um_bot_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.clk ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ena ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.k_zero ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[4].um_top_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.clk ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ena ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.k_zero ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[5].um_bot_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.clk ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ena ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.k_zero ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[5].um_top_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.clk ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ena ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.k_zero ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[6].um_bot_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.clk ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ena ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.k_zero ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[6].um_top_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.clk ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ena ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.k_zero ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[7].um_bot_I.ow[9] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.clk ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ena ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[10] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[11] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[12] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[13] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[14] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[15] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[16] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[17] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[1] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[2] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[3] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[4] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[5] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[6] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[7] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[8] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.iw[9] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.k_zero ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[0] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[10] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[11] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[12] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[13] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[14] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[15] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[16] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[17] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[18] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[19] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[1] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[20] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[21] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[22] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[23] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[2] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[3] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[4] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[5] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[6] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[7] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[8] ;
 wire \tt_top1.branch[1].col_um[7].um_top_I.ow[9] ;
 wire \tt_top1.branch[1].l_addr[0] ;
 wire \tt_top1.branch[1].l_addr[1] ;
 wire \tt_top1.spine_iw[0] ;
 wire \tt_top1.spine_iw[10] ;
 wire \tt_top1.spine_iw[11] ;
 wire \tt_top1.spine_iw[12] ;
 wire \tt_top1.spine_iw[13] ;
 wire \tt_top1.spine_iw[14] ;
 wire \tt_top1.spine_iw[15] ;
 wire \tt_top1.spine_iw[16] ;
 wire \tt_top1.spine_iw[17] ;
 wire \tt_top1.spine_iw[18] ;
 wire \tt_top1.spine_iw[19] ;
 wire \tt_top1.spine_iw[1] ;
 wire \tt_top1.spine_iw[20] ;
 wire \tt_top1.spine_iw[21] ;
 wire \tt_top1.spine_iw[22] ;
 wire \tt_top1.spine_iw[23] ;
 wire \tt_top1.spine_iw[24] ;
 wire \tt_top1.spine_iw[25] ;
 wire \tt_top1.spine_iw[26] ;
 wire \tt_top1.spine_iw[27] ;
 wire \tt_top1.spine_iw[28] ;
 wire \tt_top1.spine_iw[29] ;
 wire \tt_top1.spine_iw[2] ;
 wire \tt_top1.spine_iw[30] ;
 wire \tt_top1.spine_iw[3] ;
 wire \tt_top1.spine_iw[4] ;
 wire \tt_top1.spine_iw[5] ;
 wire \tt_top1.spine_iw[6] ;
 wire \tt_top1.spine_iw[7] ;
 wire \tt_top1.spine_iw[8] ;
 wire \tt_top1.spine_iw[9] ;
 wire \tt_top1.spine_ow[0] ;
 wire \tt_top1.spine_ow[10] ;
 wire \tt_top1.spine_ow[11] ;
 wire \tt_top1.spine_ow[12] ;
 wire \tt_top1.spine_ow[13] ;
 wire \tt_top1.spine_ow[14] ;
 wire \tt_top1.spine_ow[15] ;
 wire \tt_top1.spine_ow[16] ;
 wire \tt_top1.spine_ow[17] ;
 wire \tt_top1.spine_ow[18] ;
 wire \tt_top1.spine_ow[19] ;
 wire \tt_top1.spine_ow[1] ;
 wire \tt_top1.spine_ow[20] ;
 wire \tt_top1.spine_ow[21] ;
 wire \tt_top1.spine_ow[22] ;
 wire \tt_top1.spine_ow[23] ;
 wire \tt_top1.spine_ow[24] ;
 wire \tt_top1.spine_ow[25] ;
 wire \tt_top1.spine_ow[2] ;
 wire \tt_top1.spine_ow[3] ;
 wire \tt_top1.spine_ow[4] ;
 wire \tt_top1.spine_ow[5] ;
 wire \tt_top1.spine_ow[6] ;
 wire \tt_top1.spine_ow[7] ;
 wire \tt_top1.spine_ow[8] ;
 wire \tt_top1.spine_ow[9] ;

 tt_um_as1802 \tt_top1.branch[0].col_um[0].um_bot_I.block_0_0.tt_um_I  (.clk(\tt_top1.branch[0].col_um[0].um_bot_I.clk ),
    .ena(\tt_top1.branch[0].col_um[0].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[0].um_bot_I.iw[1] ),
    .ui_in({\tt_top1.branch[0].col_um[0].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[0].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[0].um_bot_I.ow[23] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[22] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[21] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[20] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[19] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[18] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[17] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[0].um_bot_I.ow[15] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[14] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[13] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[12] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[11] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[10] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[9] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[0].um_bot_I.ow[7] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[6] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[5] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[4] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[3] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[2] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[1] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[0] }));
 tt_um_loopback \tt_top1.branch[0].col_um[0].um_top_I.block_1_0.tt_um_I  (.clk(\tt_top1.branch[0].col_um[0].um_top_I.clk ),
    .ena(\tt_top1.branch[0].col_um[0].um_top_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[0].um_top_I.iw[1] ),
    .ui_in({\tt_top1.branch[0].col_um[0].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[0].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[0].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[0].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[0].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[0] }));
 tt_um_urish_simon \tt_top1.branch[0].col_um[1].um_bot_I.block_0_1.tt_um_I  (.clk(\tt_top1.branch[0].col_um[1].um_bot_I.clk ),
    .ena(\tt_top1.branch[0].col_um[1].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[1].um_bot_I.iw[1] ),
    .ui_in({\tt_top1.branch[0].col_um[1].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[1].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[1].um_bot_I.ow[23] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[22] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[21] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[20] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[19] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[18] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[17] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[1].um_bot_I.ow[15] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[14] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[13] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[12] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[11] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[10] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[9] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[1].um_bot_I.ow[7] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[6] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[5] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[4] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[3] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[2] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[1] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[0] }));
 tt_um_power_test \tt_top1.branch[0].col_um[1].um_top_I.block_1_1.tt_um_I  (.clk(\tt_top1.branch[0].col_um[1].um_top_I.clk ),
    .ena(\tt_top1.branch[0].col_um[1].um_top_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[1].um_top_I.iw[1] ),
    .ui_in({\tt_top1.branch[0].col_um[1].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[1].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[1].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[1].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[1].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[0] }));
 tt_um_tomkeddie_a \tt_top1.branch[0].col_um[2].um_bot_I.block_0_2.tt_um_I  (.clk(\tt_top1.branch[0].col_um[2].um_bot_I.clk ),
    .ena(\tt_top1.branch[0].col_um[2].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[2].um_bot_I.iw[1] ),
    .ui_in({\tt_top1.branch[0].col_um[2].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[2].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[2].um_bot_I.ow[23] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[22] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[21] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[20] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[19] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[18] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[17] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[2].um_bot_I.ow[15] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[14] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[13] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[12] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[11] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[10] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[9] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[2].um_bot_I.ow[7] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[6] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[5] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[4] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[3] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[2] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[1] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[0] }));
 tt_um_test \tt_top1.branch[0].col_um[2].um_top_I.block_1_2.tt_um_I  (.clk(\tt_top1.branch[0].col_um[2].um_top_I.clk ),
    .ena(\tt_top1.branch[0].col_um[2].um_top_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[2].um_top_I.iw[1] ),
    .ui_in({\tt_top1.branch[0].col_um[2].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[2].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[2].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[2].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[2].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[0] }));
 tt_um_test \tt_top1.branch[0].col_um[3].um_top_I.block_1_3.tt_um_I  (.clk(\tt_top1.branch[0].col_um[3].um_top_I.clk ),
    .ena(\tt_top1.branch[0].col_um[3].um_top_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[3].um_top_I.iw[1] ),
    .ui_in({\tt_top1.branch[0].col_um[3].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[3].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[3].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[3].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[3].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[0] }));
 tt_um_urish_dffram \tt_top1.branch[0].col_um[4].um_bot_I.block_0_4.tt_um_I  (.clk(\tt_top1.branch[0].col_um[4].um_bot_I.clk ),
    .ena(\tt_top1.branch[0].col_um[4].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[4].um_bot_I.iw[1] ),
    .ui_in({\tt_top1.branch[0].col_um[4].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[4].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[4].um_bot_I.ow[23] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[22] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[21] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[20] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[19] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[18] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[17] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[4].um_bot_I.ow[15] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[14] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[13] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[12] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[11] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[10] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[9] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[4].um_bot_I.ow[7] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[6] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[5] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[4] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[3] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[2] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[1] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[0] }));
 tt_um_test \tt_top1.branch[0].col_um[4].um_top_I.block_1_4.tt_um_I  (.clk(\tt_top1.branch[0].col_um[4].um_top_I.clk ),
    .ena(\tt_top1.branch[0].col_um[4].um_top_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[4].um_top_I.iw[1] ),
    .ui_in({\tt_top1.branch[0].col_um[4].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[4].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[4].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[4].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[4].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[0] }));
 tt_um_test \tt_top1.branch[0].col_um[5].um_top_I.block_1_5.tt_um_I  (.clk(\tt_top1.branch[0].col_um[5].um_top_I.clk ),
    .ena(\tt_top1.branch[0].col_um[5].um_top_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[5].um_top_I.iw[1] ),
    .ui_in({\tt_top1.branch[0].col_um[5].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[5].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[5].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[5].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[5].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[0] }));
 tt_um_test \tt_top1.branch[0].col_um[6].um_top_I.block_1_6.tt_um_I  (.clk(\tt_top1.branch[0].col_um[6].um_top_I.clk ),
    .ena(\tt_top1.branch[0].col_um[6].um_top_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[6].um_top_I.iw[1] ),
    .ui_in({\tt_top1.branch[0].col_um[6].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[6].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[6].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[6].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[6].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[0] }));
 tt_um_test \tt_top1.branch[0].col_um[7].um_top_I.block_1_7.tt_um_I  (.clk(\tt_top1.branch[0].col_um[7].um_top_I.clk ),
    .ena(\tt_top1.branch[0].col_um[7].um_top_I.ena ),
    .rst_n(\tt_top1.branch[0].col_um[7].um_top_I.iw[1] ),
    .ui_in({\tt_top1.branch[0].col_um[7].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[0].col_um[7].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[0].col_um[7].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[0].col_um[7].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[0].col_um[7].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[0] }));
 tt_mux \tt_top1.branch[0].mux_I  (.k_one(\tt_top1.branch[0].l_k_one ),
    .k_zero(\tt_top1.branch[0].l_addr[0] ),
    .addr({\tt_top1.branch[0].l_addr[0] ,
    \tt_top1.branch[0].l_addr[0] ,
    \tt_top1.branch[0].l_addr[0] ,
    \tt_top1.branch[0].l_addr[0] ,
    \tt_top1.branch[0].l_addr[0] }),
    .spine_iw({\tt_top1.spine_iw[30] ,
    \tt_top1.spine_iw[29] ,
    \tt_top1.spine_iw[28] ,
    \tt_top1.spine_iw[27] ,
    \tt_top1.spine_iw[26] ,
    \tt_top1.spine_iw[25] ,
    \tt_top1.spine_iw[24] ,
    \tt_top1.spine_iw[23] ,
    \tt_top1.spine_iw[22] ,
    \tt_top1.spine_iw[21] ,
    \tt_top1.spine_iw[20] ,
    \tt_top1.spine_iw[19] ,
    \tt_top1.spine_iw[18] ,
    \tt_top1.spine_iw[17] ,
    \tt_top1.spine_iw[16] ,
    \tt_top1.spine_iw[15] ,
    \tt_top1.spine_iw[14] ,
    \tt_top1.spine_iw[13] ,
    \tt_top1.spine_iw[12] ,
    \tt_top1.spine_iw[11] ,
    \tt_top1.spine_iw[10] ,
    \tt_top1.spine_iw[9] ,
    \tt_top1.spine_iw[8] ,
    \tt_top1.spine_iw[7] ,
    \tt_top1.spine_iw[6] ,
    \tt_top1.spine_iw[5] ,
    \tt_top1.spine_iw[4] ,
    \tt_top1.spine_iw[3] ,
    \tt_top1.spine_iw[2] ,
    \tt_top1.spine_iw[1] ,
    \tt_top1.spine_iw[0] }),
    .spine_ow({\tt_top1.spine_ow[25] ,
    \tt_top1.spine_ow[24] ,
    \tt_top1.spine_ow[23] ,
    \tt_top1.spine_ow[22] ,
    \tt_top1.spine_ow[21] ,
    \tt_top1.spine_ow[20] ,
    \tt_top1.spine_ow[19] ,
    \tt_top1.spine_ow[18] ,
    \tt_top1.spine_ow[17] ,
    \tt_top1.spine_ow[16] ,
    \tt_top1.spine_ow[15] ,
    \tt_top1.spine_ow[14] ,
    \tt_top1.spine_ow[13] ,
    \tt_top1.spine_ow[12] ,
    \tt_top1.spine_ow[11] ,
    \tt_top1.spine_ow[10] ,
    \tt_top1.spine_ow[9] ,
    \tt_top1.spine_ow[8] ,
    \tt_top1.spine_ow[7] ,
    \tt_top1.spine_ow[6] ,
    \tt_top1.spine_ow[5] ,
    \tt_top1.spine_ow[4] ,
    \tt_top1.spine_ow[3] ,
    \tt_top1.spine_ow[2] ,
    \tt_top1.spine_ow[1] ,
    \tt_top1.spine_ow[0] }),
    .um_ena({\tt_top1.branch[0].col_um[7].um_top_I.ena ,
    \tt_top1.branch[0].col_um[7].um_bot_I.ena ,
    \tt_top1.branch[0].col_um[6].um_top_I.ena ,
    \tt_top1.branch[0].col_um[6].um_bot_I.ena ,
    \tt_top1.branch[0].col_um[5].um_top_I.ena ,
    \tt_top1.branch[0].col_um[5].um_bot_I.ena ,
    \tt_top1.branch[0].col_um[4].um_top_I.ena ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ena ,
    \tt_top1.branch[0].col_um[3].um_top_I.ena ,
    \tt_top1.branch[0].col_um[3].um_bot_I.ena ,
    \tt_top1.branch[0].col_um[2].um_top_I.ena ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ena ,
    \tt_top1.branch[0].col_um[1].um_top_I.ena ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ena ,
    \tt_top1.branch[0].col_um[0].um_top_I.ena ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ena }),
    .um_iw({\tt_top1.branch[0].col_um[7].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[10] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[2] ,
    \tt_top1.branch[0].col_um[7].um_top_I.iw[1] ,
    \tt_top1.branch[0].col_um[7].um_top_I.clk ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[10] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[2] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.iw[1] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.clk ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[10] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[2] ,
    \tt_top1.branch[0].col_um[6].um_top_I.iw[1] ,
    \tt_top1.branch[0].col_um[6].um_top_I.clk ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[10] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[2] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.iw[1] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.clk ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[10] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[2] ,
    \tt_top1.branch[0].col_um[5].um_top_I.iw[1] ,
    \tt_top1.branch[0].col_um[5].um_top_I.clk ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[10] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[2] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.iw[1] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.clk ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[10] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[2] ,
    \tt_top1.branch[0].col_um[4].um_top_I.iw[1] ,
    \tt_top1.branch[0].col_um[4].um_top_I.clk ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[10] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[2] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.iw[1] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.clk ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[10] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[2] ,
    \tt_top1.branch[0].col_um[3].um_top_I.iw[1] ,
    \tt_top1.branch[0].col_um[3].um_top_I.clk ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[10] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[2] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.iw[1] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.clk ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[10] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[2] ,
    \tt_top1.branch[0].col_um[2].um_top_I.iw[1] ,
    \tt_top1.branch[0].col_um[2].um_top_I.clk ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[10] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[2] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.iw[1] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.clk ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[10] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[2] ,
    \tt_top1.branch[0].col_um[1].um_top_I.iw[1] ,
    \tt_top1.branch[0].col_um[1].um_top_I.clk ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[10] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[2] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.iw[1] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.clk ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[17] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[16] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[15] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[14] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[13] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[12] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[11] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[10] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[9] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[8] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[7] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[6] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[5] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[4] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[3] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[2] ,
    \tt_top1.branch[0].col_um[0].um_top_I.iw[1] ,
    \tt_top1.branch[0].col_um[0].um_top_I.clk ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[17] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[16] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[15] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[14] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[13] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[12] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[11] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[10] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[9] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[8] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[7] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[6] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[5] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[4] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[3] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[2] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.iw[1] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.clk }),
    .um_k_zero({\tt_top1.branch[0].col_um[7].um_top_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_top_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_top_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[4].um_top_I.k_zero ,
    \tt_top1.branch[0].col_um[4].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_top_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[2].um_top_I.k_zero ,
    \tt_top1.branch[0].col_um[2].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[1].um_top_I.k_zero ,
    \tt_top1.branch[0].col_um[1].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[0].um_top_I.k_zero ,
    \tt_top1.branch[0].col_um[0].um_bot_I.k_zero }),
    .um_ow({\tt_top1.branch[0].col_um[7].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[16] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[8] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[7].um_top_I.ow[0] ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[16] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[8] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[6].um_top_I.ow[0] ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[16] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[8] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[5].um_top_I.ow[0] ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[16] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[8] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[4].um_top_I.ow[0] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[23] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[22] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[21] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[20] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[19] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[18] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[17] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[16] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[15] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[14] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[13] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[12] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[11] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[10] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[9] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[8] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[7] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[6] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[5] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[4] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[3] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[2] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[1] ,
    \tt_top1.branch[0].col_um[4].um_bot_I.ow[0] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[16] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[8] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[3].um_top_I.ow[0] ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[16] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[8] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[2].um_top_I.ow[0] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[23] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[22] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[21] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[20] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[19] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[18] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[17] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[16] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[15] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[14] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[13] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[12] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[11] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[10] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[9] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[8] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[7] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[6] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[5] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[4] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[3] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[2] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[1] ,
    \tt_top1.branch[0].col_um[2].um_bot_I.ow[0] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[16] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[8] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[1].um_top_I.ow[0] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[23] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[22] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[21] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[20] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[19] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[18] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[17] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[16] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[15] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[14] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[13] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[12] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[11] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[10] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[9] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[8] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[7] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[6] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[5] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[4] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[3] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[2] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[1] ,
    \tt_top1.branch[0].col_um[1].um_bot_I.ow[0] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[23] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[22] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[21] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[20] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[19] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[18] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[17] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[16] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[15] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[14] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[13] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[12] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[11] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[10] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[9] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[8] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[7] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[6] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[5] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[4] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[3] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[2] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[1] ,
    \tt_top1.branch[0].col_um[0].um_top_I.ow[0] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[23] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[22] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[21] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[20] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[19] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[18] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[17] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[16] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[15] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[14] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[13] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[12] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[11] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[10] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[9] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[8] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[7] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[6] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[5] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[4] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[3] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[2] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[1] ,
    \tt_top1.branch[0].col_um[0].um_bot_I.ow[0] }));
 tt_um_TrainLED2_top \tt_top1.branch[1].col_um[0].um_bot_I.block_0_16.tt_um_I  (.clk(\tt_top1.branch[1].col_um[0].um_bot_I.clk ),
    .ena(\tt_top1.branch[1].col_um[0].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[0].um_bot_I.iw[1] ),
    .ui_in({\tt_top1.branch[1].col_um[0].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[0].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[0].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[0].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[0].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[0] }));
 tt_um_loopback \tt_top1.branch[1].col_um[0].um_top_I.block_1_16.tt_um_I  (.clk(\tt_top1.branch[1].col_um[0].um_top_I.clk ),
    .ena(\tt_top1.branch[1].col_um[0].um_top_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[0].um_top_I.iw[1] ),
    .ui_in({\tt_top1.branch[1].col_um[0].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[0].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[0].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[0].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[0].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[0] }));
 tt_um_moyes0_top_module \tt_top1.branch[1].col_um[1].um_bot_I.block_0_17.tt_um_I  (.clk(\tt_top1.branch[1].col_um[1].um_bot_I.clk ),
    .ena(\tt_top1.branch[1].col_um[1].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[1].um_bot_I.iw[1] ),
    .ui_in({\tt_top1.branch[1].col_um[1].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[1].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[1].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[1].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[1].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[0] }));
 tt_um_test \tt_top1.branch[1].col_um[1].um_top_I.block_1_17.tt_um_I  (.clk(\tt_top1.branch[1].col_um[1].um_top_I.clk ),
    .ena(\tt_top1.branch[1].col_um[1].um_top_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[1].um_top_I.iw[1] ),
    .ui_in({\tt_top1.branch[1].col_um[1].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[1].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[1].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[1].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[1].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[0] }));
 tt_um_vga_clock \tt_top1.branch[1].col_um[2].um_bot_I.block_0_18.tt_um_I  (.clk(\tt_top1.branch[1].col_um[2].um_bot_I.clk ),
    .ena(\tt_top1.branch[1].col_um[2].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[2].um_bot_I.iw[1] ),
    .ui_in({\tt_top1.branch[1].col_um[2].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[2].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[2].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[2].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[2].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[0] }));
 tt_um_test \tt_top1.branch[1].col_um[2].um_top_I.block_1_18.tt_um_I  (.clk(\tt_top1.branch[1].col_um[2].um_top_I.clk ),
    .ena(\tt_top1.branch[1].col_um[2].um_top_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[2].um_top_I.iw[1] ),
    .ui_in({\tt_top1.branch[1].col_um[2].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[2].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[2].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[2].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[2].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[0] }));
 tt_um_kiwih_tt_top \tt_top1.branch[1].col_um[3].um_bot_I.block_0_19.tt_um_I  (.clk(\tt_top1.branch[1].col_um[3].um_bot_I.clk ),
    .ena(\tt_top1.branch[1].col_um[3].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[3].um_bot_I.iw[1] ),
    .ui_in({\tt_top1.branch[1].col_um[3].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[3].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[3].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[3].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[3].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[0] }));
 tt_um_test \tt_top1.branch[1].col_um[3].um_top_I.block_1_19.tt_um_I  (.clk(\tt_top1.branch[1].col_um[3].um_top_I.clk ),
    .ena(\tt_top1.branch[1].col_um[3].um_top_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[3].um_top_I.iw[1] ),
    .ui_in({\tt_top1.branch[1].col_um[3].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[3].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[3].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[3].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[3].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[0] }));
 tt_um_ternaryPC_radixconvert \tt_top1.branch[1].col_um[4].um_bot_I.block_0_20.tt_um_I  (.clk(\tt_top1.branch[1].col_um[4].um_bot_I.clk ),
    .ena(\tt_top1.branch[1].col_um[4].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[4].um_bot_I.iw[1] ),
    .ui_in({\tt_top1.branch[1].col_um[4].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[4].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[4].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[4].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[4].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[0] }));
 tt_um_test \tt_top1.branch[1].col_um[4].um_top_I.block_1_20.tt_um_I  (.clk(\tt_top1.branch[1].col_um[4].um_top_I.clk ),
    .ena(\tt_top1.branch[1].col_um[4].um_top_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[4].um_top_I.iw[1] ),
    .ui_in({\tt_top1.branch[1].col_um[4].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[4].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[4].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[4].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[4].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[0] }));
 tt_um_wokwi_366318576852367361 \tt_top1.branch[1].col_um[5].um_bot_I.block_0_21.tt_um_I  (.clk(\tt_top1.branch[1].col_um[5].um_bot_I.clk ),
    .ena(\tt_top1.branch[1].col_um[5].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[5].um_bot_I.iw[1] ),
    .ui_in({\tt_top1.branch[1].col_um[5].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[5].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[5].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[5].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[5].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[0] }));
 tt_um_test \tt_top1.branch[1].col_um[5].um_top_I.block_1_21.tt_um_I  (.clk(\tt_top1.branch[1].col_um[5].um_top_I.clk ),
    .ena(\tt_top1.branch[1].col_um[5].um_top_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[5].um_top_I.iw[1] ),
    .ui_in({\tt_top1.branch[1].col_um[5].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[5].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[5].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[5].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[5].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[0] }));
 tt_um_MichaelBell_hovalaag \tt_top1.branch[1].col_um[6].um_bot_I.block_0_22.tt_um_I  (.clk(\tt_top1.branch[1].col_um[6].um_bot_I.clk ),
    .ena(\tt_top1.branch[1].col_um[6].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[6].um_bot_I.iw[1] ),
    .ui_in({\tt_top1.branch[1].col_um[6].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[6].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[6].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[6].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[6].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[0] }));
 tt_um_test \tt_top1.branch[1].col_um[6].um_top_I.block_1_22.tt_um_I  (.clk(\tt_top1.branch[1].col_um[6].um_top_I.clk ),
    .ena(\tt_top1.branch[1].col_um[6].um_top_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[6].um_top_I.iw[1] ),
    .ui_in({\tt_top1.branch[1].col_um[6].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[6].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[6].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[6].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[6].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[0] }));
 tt_um_cam \tt_top1.branch[1].col_um[7].um_bot_I.block_0_23.tt_um_I  (.clk(\tt_top1.branch[1].col_um[7].um_bot_I.clk ),
    .ena(\tt_top1.branch[1].col_um[7].um_bot_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[7].um_bot_I.iw[1] ),
    .ui_in({\tt_top1.branch[1].col_um[7].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[7].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[7].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[7].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[7].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[0] }));
 tt_um_test \tt_top1.branch[1].col_um[7].um_top_I.block_1_23.tt_um_I  (.clk(\tt_top1.branch[1].col_um[7].um_top_I.clk ),
    .ena(\tt_top1.branch[1].col_um[7].um_top_I.ena ),
    .rst_n(\tt_top1.branch[1].col_um[7].um_top_I.iw[1] ),
    .ui_in({\tt_top1.branch[1].col_um[7].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[2] }),
    .uio_in({\tt_top1.branch[1].col_um[7].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[10] }),
    .uio_oe({\tt_top1.branch[1].col_um[7].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[16] }),
    .uio_out({\tt_top1.branch[1].col_um[7].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[8] }),
    .uo_out({\tt_top1.branch[1].col_um[7].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[0] }));
 tt_mux \tt_top1.branch[1].mux_I  (.k_one(\tt_top1.branch[1].l_addr[0] ),
    .k_zero(\tt_top1.branch[1].l_addr[1] ),
    .addr({\tt_top1.branch[1].l_addr[1] ,
    \tt_top1.branch[1].l_addr[1] ,
    \tt_top1.branch[1].l_addr[1] ,
    \tt_top1.branch[1].l_addr[1] ,
    \tt_top1.branch[1].l_addr[0] }),
    .spine_iw({\tt_top1.spine_iw[30] ,
    \tt_top1.spine_iw[29] ,
    \tt_top1.spine_iw[28] ,
    \tt_top1.spine_iw[27] ,
    \tt_top1.spine_iw[26] ,
    \tt_top1.spine_iw[25] ,
    \tt_top1.spine_iw[24] ,
    \tt_top1.spine_iw[23] ,
    \tt_top1.spine_iw[22] ,
    \tt_top1.spine_iw[21] ,
    \tt_top1.spine_iw[20] ,
    \tt_top1.spine_iw[19] ,
    \tt_top1.spine_iw[18] ,
    \tt_top1.spine_iw[17] ,
    \tt_top1.spine_iw[16] ,
    \tt_top1.spine_iw[15] ,
    \tt_top1.spine_iw[14] ,
    \tt_top1.spine_iw[13] ,
    \tt_top1.spine_iw[12] ,
    \tt_top1.spine_iw[11] ,
    \tt_top1.spine_iw[10] ,
    \tt_top1.spine_iw[9] ,
    \tt_top1.spine_iw[8] ,
    \tt_top1.spine_iw[7] ,
    \tt_top1.spine_iw[6] ,
    \tt_top1.spine_iw[5] ,
    \tt_top1.spine_iw[4] ,
    \tt_top1.spine_iw[3] ,
    \tt_top1.spine_iw[2] ,
    \tt_top1.spine_iw[1] ,
    \tt_top1.spine_iw[0] }),
    .spine_ow({\tt_top1.spine_ow[25] ,
    \tt_top1.spine_ow[24] ,
    \tt_top1.spine_ow[23] ,
    \tt_top1.spine_ow[22] ,
    \tt_top1.spine_ow[21] ,
    \tt_top1.spine_ow[20] ,
    \tt_top1.spine_ow[19] ,
    \tt_top1.spine_ow[18] ,
    \tt_top1.spine_ow[17] ,
    \tt_top1.spine_ow[16] ,
    \tt_top1.spine_ow[15] ,
    \tt_top1.spine_ow[14] ,
    \tt_top1.spine_ow[13] ,
    \tt_top1.spine_ow[12] ,
    \tt_top1.spine_ow[11] ,
    \tt_top1.spine_ow[10] ,
    \tt_top1.spine_ow[9] ,
    \tt_top1.spine_ow[8] ,
    \tt_top1.spine_ow[7] ,
    \tt_top1.spine_ow[6] ,
    \tt_top1.spine_ow[5] ,
    \tt_top1.spine_ow[4] ,
    \tt_top1.spine_ow[3] ,
    \tt_top1.spine_ow[2] ,
    \tt_top1.spine_ow[1] ,
    \tt_top1.spine_ow[0] }),
    .um_ena({\tt_top1.branch[1].col_um[7].um_top_I.ena ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ena ,
    \tt_top1.branch[1].col_um[6].um_top_I.ena ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ena ,
    \tt_top1.branch[1].col_um[5].um_top_I.ena ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ena ,
    \tt_top1.branch[1].col_um[4].um_top_I.ena ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ena ,
    \tt_top1.branch[1].col_um[3].um_top_I.ena ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ena ,
    \tt_top1.branch[1].col_um[2].um_top_I.ena ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ena ,
    \tt_top1.branch[1].col_um[1].um_top_I.ena ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ena ,
    \tt_top1.branch[1].col_um[0].um_top_I.ena ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ena }),
    .um_iw({\tt_top1.branch[1].col_um[7].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[10] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[2] ,
    \tt_top1.branch[1].col_um[7].um_top_I.iw[1] ,
    \tt_top1.branch[1].col_um[7].um_top_I.clk ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[10] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[2] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.iw[1] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.clk ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[10] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[2] ,
    \tt_top1.branch[1].col_um[6].um_top_I.iw[1] ,
    \tt_top1.branch[1].col_um[6].um_top_I.clk ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[10] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[2] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.iw[1] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.clk ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[10] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[2] ,
    \tt_top1.branch[1].col_um[5].um_top_I.iw[1] ,
    \tt_top1.branch[1].col_um[5].um_top_I.clk ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[10] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[2] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.iw[1] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.clk ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[10] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[2] ,
    \tt_top1.branch[1].col_um[4].um_top_I.iw[1] ,
    \tt_top1.branch[1].col_um[4].um_top_I.clk ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[10] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[2] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.iw[1] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.clk ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[10] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[2] ,
    \tt_top1.branch[1].col_um[3].um_top_I.iw[1] ,
    \tt_top1.branch[1].col_um[3].um_top_I.clk ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[10] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[2] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.iw[1] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.clk ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[10] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[2] ,
    \tt_top1.branch[1].col_um[2].um_top_I.iw[1] ,
    \tt_top1.branch[1].col_um[2].um_top_I.clk ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[10] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[2] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.iw[1] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.clk ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[10] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[2] ,
    \tt_top1.branch[1].col_um[1].um_top_I.iw[1] ,
    \tt_top1.branch[1].col_um[1].um_top_I.clk ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[10] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[2] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.iw[1] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.clk ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[17] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[16] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[15] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[14] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[13] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[12] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[11] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[10] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[9] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[8] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[7] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[6] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[5] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[4] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[3] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[2] ,
    \tt_top1.branch[1].col_um[0].um_top_I.iw[1] ,
    \tt_top1.branch[1].col_um[0].um_top_I.clk ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[17] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[16] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[15] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[14] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[13] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[12] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[11] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[10] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[9] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[8] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[7] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[6] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[5] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[4] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[3] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[2] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.iw[1] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.clk }),
    .um_k_zero({\tt_top1.branch[1].col_um[7].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[7].um_bot_I.k_zero ,
    \tt_top1.branch[1].col_um[6].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[6].um_bot_I.k_zero ,
    \tt_top1.branch[1].col_um[5].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[5].um_bot_I.k_zero ,
    \tt_top1.branch[1].col_um[4].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[4].um_bot_I.k_zero ,
    \tt_top1.branch[1].col_um[3].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[3].um_bot_I.k_zero ,
    \tt_top1.branch[1].col_um[2].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[2].um_bot_I.k_zero ,
    \tt_top1.branch[1].col_um[1].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[1].um_bot_I.k_zero ,
    \tt_top1.branch[1].col_um[0].um_top_I.k_zero ,
    \tt_top1.branch[1].col_um[0].um_bot_I.k_zero }),
    .um_ow({\tt_top1.branch[1].col_um[7].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[16] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[8] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[7].um_top_I.ow[0] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[16] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[8] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[7].um_bot_I.ow[0] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[16] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[8] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[6].um_top_I.ow[0] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[16] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[8] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[6].um_bot_I.ow[0] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[16] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[8] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[5].um_top_I.ow[0] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[16] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[8] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[5].um_bot_I.ow[0] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[16] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[8] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[4].um_top_I.ow[0] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[16] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[8] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[4].um_bot_I.ow[0] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[16] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[8] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[3].um_top_I.ow[0] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[16] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[8] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[3].um_bot_I.ow[0] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[16] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[8] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[2].um_top_I.ow[0] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[16] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[8] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[2].um_bot_I.ow[0] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[16] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[8] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[1].um_top_I.ow[0] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[16] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[8] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[1].um_bot_I.ow[0] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[23] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[22] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[21] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[20] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[19] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[18] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[17] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[16] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[15] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[14] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[13] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[12] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[11] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[10] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[9] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[8] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[7] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[6] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[5] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[4] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[3] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[2] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[1] ,
    \tt_top1.branch[1].col_um[0].um_top_I.ow[0] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[23] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[22] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[21] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[20] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[19] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[18] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[17] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[16] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[15] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[14] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[13] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[12] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[11] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[10] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[9] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[8] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[7] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[6] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[5] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[4] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[3] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[2] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[1] ,
    \tt_top1.branch[1].col_um[0].um_bot_I.ow[0] }));
 tt_ctrl \tt_top1.ctrl_I  (.ctrl_ena(io_in[32]),
    .ctrl_sel_inc(io_in[34]),
    .ctrl_sel_rst_n(io_in[36]),
    .k_one(\tt_top1.io_oeb[0] ),
    .k_zero(\tt_top1.io_oeb[16] ),
    .pad_ui_in({io_in[15],
    io_in[14],
    io_in[13],
    io_in[12],
    io_in[11],
    io_in[10],
    io_in[9],
    io_in[8],
    io_in[7],
    io_in[6]}),
    .pad_uio_in({io_in[31],
    io_in[30],
    io_in[29],
    io_in[28],
    io_in[27],
    io_in[26],
    io_in[25],
    io_in[24]}),
    .pad_uio_oe_n({io_oeb[31],
    io_oeb[30],
    io_oeb[29],
    io_oeb[28],
    io_oeb[27],
    io_oeb[26],
    io_oeb[25],
    io_oeb[24]}),
    .pad_uio_out({io_out[31],
    io_out[30],
    io_out[29],
    io_out[28],
    io_out[27],
    io_out[26],
    io_out[25],
    io_out[24]}),
    .pad_uo_out({io_out[23],
    io_out[22],
    io_out[21],
    io_out[20],
    io_out[19],
    io_out[18],
    io_out[17],
    io_out[16]}),
    .spine_iw({\tt_top1.spine_iw[30] ,
    \tt_top1.spine_iw[29] ,
    \tt_top1.spine_iw[28] ,
    \tt_top1.spine_iw[27] ,
    \tt_top1.spine_iw[26] ,
    \tt_top1.spine_iw[25] ,
    \tt_top1.spine_iw[24] ,
    \tt_top1.spine_iw[23] ,
    \tt_top1.spine_iw[22] ,
    \tt_top1.spine_iw[21] ,
    \tt_top1.spine_iw[20] ,
    \tt_top1.spine_iw[19] ,
    \tt_top1.spine_iw[18] ,
    \tt_top1.spine_iw[17] ,
    \tt_top1.spine_iw[16] ,
    \tt_top1.spine_iw[15] ,
    \tt_top1.spine_iw[14] ,
    \tt_top1.spine_iw[13] ,
    \tt_top1.spine_iw[12] ,
    \tt_top1.spine_iw[11] ,
    \tt_top1.spine_iw[10] ,
    \tt_top1.spine_iw[9] ,
    \tt_top1.spine_iw[8] ,
    \tt_top1.spine_iw[7] ,
    \tt_top1.spine_iw[6] ,
    \tt_top1.spine_iw[5] ,
    \tt_top1.spine_iw[4] ,
    \tt_top1.spine_iw[3] ,
    \tt_top1.spine_iw[2] ,
    \tt_top1.spine_iw[1] ,
    \tt_top1.spine_iw[0] }),
    .spine_ow({\tt_top1.spine_ow[25] ,
    \tt_top1.spine_ow[24] ,
    \tt_top1.spine_ow[23] ,
    \tt_top1.spine_ow[22] ,
    \tt_top1.spine_ow[21] ,
    \tt_top1.spine_ow[20] ,
    \tt_top1.spine_ow[19] ,
    \tt_top1.spine_ow[18] ,
    \tt_top1.spine_ow[17] ,
    \tt_top1.spine_ow[16] ,
    \tt_top1.spine_ow[15] ,
    \tt_top1.spine_ow[14] ,
    \tt_top1.spine_ow[13] ,
    \tt_top1.spine_ow[12] ,
    \tt_top1.spine_ow[11] ,
    \tt_top1.spine_ow[10] ,
    \tt_top1.spine_ow[9] ,
    \tt_top1.spine_ow[8] ,
    \tt_top1.spine_ow[7] ,
    \tt_top1.spine_ow[6] ,
    \tt_top1.spine_ow[5] ,
    \tt_top1.spine_ow[4] ,
    \tt_top1.spine_ow[3] ,
    \tt_top1.spine_ow[2] ,
    \tt_top1.spine_ow[1] ,
    \tt_top1.spine_ow[0] }));
 assign io_oeb[0] = \tt_top1.io_oeb[0] ;
 assign io_oeb[10] = \tt_top1.io_oeb[0] ;
 assign io_oeb[11] = \tt_top1.io_oeb[0] ;
 assign io_oeb[12] = \tt_top1.io_oeb[0] ;
 assign io_oeb[13] = \tt_top1.io_oeb[0] ;
 assign io_oeb[14] = \tt_top1.io_oeb[0] ;
 assign io_oeb[15] = \tt_top1.io_oeb[0] ;
 assign io_oeb[16] = \tt_top1.io_oeb[16] ;
 assign io_oeb[17] = \tt_top1.io_oeb[16] ;
 assign io_oeb[18] = \tt_top1.io_oeb[16] ;
 assign io_oeb[19] = \tt_top1.io_oeb[16] ;
 assign io_oeb[1] = \tt_top1.io_oeb[0] ;
 assign io_oeb[20] = \tt_top1.io_oeb[16] ;
 assign io_oeb[21] = \tt_top1.io_oeb[16] ;
 assign io_oeb[22] = \tt_top1.io_oeb[16] ;
 assign io_oeb[23] = \tt_top1.io_oeb[16] ;
 assign io_oeb[2] = \tt_top1.io_oeb[0] ;
 assign io_oeb[32] = \tt_top1.io_oeb[0] ;
 assign io_oeb[33] = \tt_top1.io_oeb[16] ;
 assign io_oeb[34] = \tt_top1.io_oeb[0] ;
 assign io_oeb[35] = \tt_top1.io_oeb[16] ;
 assign io_oeb[36] = \tt_top1.io_oeb[0] ;
 assign io_oeb[37] = \tt_top1.io_oeb[16] ;
 assign io_oeb[3] = \tt_top1.io_oeb[0] ;
 assign io_oeb[4] = \tt_top1.io_oeb[16] ;
 assign io_oeb[5] = \tt_top1.io_oeb[16] ;
 assign io_oeb[6] = \tt_top1.io_oeb[0] ;
 assign io_oeb[7] = \tt_top1.io_oeb[0] ;
 assign io_oeb[8] = \tt_top1.io_oeb[0] ;
 assign io_oeb[9] = \tt_top1.io_oeb[0] ;
 assign io_out[0] = \tt_top1.io_oeb[0] ;
 assign io_out[10] = \tt_top1.io_oeb[0] ;
 assign io_out[11] = \tt_top1.io_oeb[0] ;
 assign io_out[12] = \tt_top1.io_oeb[0] ;
 assign io_out[13] = \tt_top1.io_oeb[0] ;
 assign io_out[14] = \tt_top1.io_oeb[0] ;
 assign io_out[15] = \tt_top1.io_oeb[0] ;
 assign io_out[1] = \tt_top1.io_oeb[0] ;
 assign io_out[2] = \tt_top1.io_oeb[0] ;
 assign io_out[32] = \tt_top1.io_oeb[16] ;
 assign io_out[33] = \tt_top1.io_oeb[16] ;
 assign io_out[34] = \tt_top1.io_oeb[16] ;
 assign io_out[35] = \tt_top1.io_oeb[16] ;
 assign io_out[36] = \tt_top1.io_oeb[16] ;
 assign io_out[37] = \tt_top1.io_oeb[16] ;
 assign io_out[3] = \tt_top1.io_oeb[0] ;
 assign io_out[4] = \tt_top1.io_oeb[16] ;
 assign io_out[5] = user_clock2;
 assign io_out[6] = \tt_top1.io_oeb[0] ;
 assign io_out[7] = \tt_top1.io_oeb[0] ;
 assign io_out[8] = \tt_top1.io_oeb[0] ;
 assign io_out[9] = \tt_top1.io_oeb[0] ;
endmodule

